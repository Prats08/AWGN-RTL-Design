/* Top Level for AWGN */

module AWGN(input clk, input reset, output reg Valid, output reg [15:0] X0_Out, output reg [15:0] X1_Out);

wire [31:0] Taus1, Taus2;
reg [47:0] LogIn;
wire [30:0] LogOut;
reg [30:0] LogOut2;
wire [16:0] SqrtOut;
wire [15:0] Sin11, Cos11;

reg [15:0] Angle, X0, X1, X01, X11;
reg [15:0] Sin, Sin1, Sin2, Sin3, Sin4, Sin5, Sin6, Sin7, Sin8;
reg [15:0] Cos, Cos1, Cos2, Cos3, Cos4, Cos5, Cos6, Cos7, Cos8;
reg [31:0] RegX0, RegX1;


reg Valid0, Valid1, Valid2, Valid3, Valid4, Valid5, Valid6, Valid7, Valid8, Valid9, Valid10, Valid11, Valid12, Valid13, Valid14, Valid15;

always @(posedge clk)
begin

		Valid0 <= !reset;
		Valid1 <= Valid0;
		Valid2 <= Valid1;
		Valid3 <= Valid2;
		Valid4 <= Valid3;
		Valid5 <= Valid4;
		Valid6 <= Valid5;
		Valid7 <= Valid6;
		Valid8 <= Valid7;
		Valid9 <= Valid8;
		Valid10 <= Valid9;
		Valid11 <= Valid10;
		Valid12 <= Valid11;
		Valid13 <= Valid12;
		Valid14 <= Valid13;
		Valid15 <= Valid14;
		Valid <= Valid15;

	if(!reset)
	begin

		// Cycle 1 Taus

		// Cycle 2
		LogIn <= {Taus1[31:0], Taus2[31:16]};
		Angle <= Taus2[15:0];
		
		// Pipelining
		Sin2 <= Sin11;	Cos2 <= Cos11;	// 3 Cycles	
		Sin3 <= Sin2;	Cos3 <= Cos2;	// 4 Cycles	
		Sin4 <= Sin3;	Cos4 <= Cos3;	// 5 Cycles
		Sin5 <= Sin4;	Cos5 <= Cos4;	// 6 Cycles
		Sin6 <= Sin5;	Cos6 <= Cos5;	// 7 Cycles
		Sin7 <= Sin6;	Cos7 <= Cos6;	// 8 Cycles
		Sin8 <= Sin7;	Cos8 <= Cos7;	// 9 Cycles
		Sin <= Sin8;	Cos <= Cos8;	// 10 Cycles
//		Sin <= Sin1;	Cos <= Cos1;	// 11 Cycles

		LogOut2 <= LogOut;		// Register between Log and Cosine Block

		// Cycle 12
		X0[15] <= Sin[15];
		X1[15] <= Cos[15];


		RegX0 <= Sin[14:0] * SqrtOut[16:0];
		RegX1 <= Cos[14:0] * SqrtOut[16:0];

		// Cycle 13		 
		X0[14:11] <= RegX0[31:28];
		X0[10:0] <= RegX0[27:17];

		X1[14:11] <= RegX1[31:28];
		X1[10:0] <= RegX1[27:17];

		// Cycle 14

		X01 <= X0;
		X11 <= X1;

		// Cycle 15

		X0_Out <= X01;
		X1_Out <= X11;

	end // reset

	else begin
		Valid <= 1'b0;
		Valid0 <= 1'b0;
		Valid1 <= 1'b0;
		Valid2 <= 1'b0;
		Valid3 <= 1'b0;
		Valid4 <= 1'b0;
		Valid5 <= 1'b0;
		Valid6 <= 1'b0;
		Valid7 <= 1'b0;
		Valid8 <= 1'b0;
		Valid9 <= 1'b0;
		Valid10 <= 1'b0;
		Valid11 <= 1'b0;
		Valid12 <= 1'b0;
		Valid13 <= 1'b0;
		Valid14 <= 1'b0;
		Valid15 <= 1'b0;

		X0_Out <= 15'b0;
		X1_Out <= 15'b0;
	end

end

Taus T1(clk, reset, Taus1[31:0]);	// 1 Cycle
Taus T2(clk, reset, Taus2[31:0]);	// 1 Cycle

LOG_POLY L1(clk, reset, LogIn, LogOut);		// 6 Cycles + 1 Cycle
SQRT_POLY S1(clk,reset, LogOut2, SqrtOut);	// 3 Cycles

SinBlock SinInst1(clk,reset, 1'b0, Angle, Sin11);	// 2 Cycle
SinBlock CosInst1(clk,reset, 1'b1, Angle, Cos11);	// 2 Cycle

endmodule

/* 32-bit Tausworthe Uniform Random Number Generator */

module Taus(input clk, input reset, output reg [31:0] Tout);

	reg [31:0] s0, s1, s2, b0, b1, b2;

always @(posedge clk) begin

	if(!reset)


	begin

		b0 <= ((( s0 << 13) ^ s0) >> 19);

		s0 <= ((( s0 & 32'hFFFFFFFE) << 12 ) ^ b0);

		b1 <= ((( s1 << 2) ^ s1) >> 25);

		s1 <= ((( s1 & 32'hFFFF_FFF8) << 4 ) ^ b1);

		b2 <= ((( s2 << 3) ^ s2) >> 11);
	
		s2 <= ((( s2 & 32'hFFFF_FFF0) << 17 ) ^ b2);


		Tout <= s0 ^ s1 ^ s2;

	end

	else begin

		b0 <= 32'b00000000_00000000_00000000_00000000;
		b1 <= 32'b00000000_00000000_00000000_00000000;
		b2 <= 32'b00000000_00000000_00000000_00000000;
		s0 <= 32'b00000000_00000000_00000000_00000010;
		s1 <= 32'b00000000_00000000_00000000_00000111;
		s2 <= 32'b00000000_00000000_00000000_00000101;
	end
end


endmodule


/* Verilog code for The Logarithm block of AWGN Project

	Log takes input of 48 bits in Q48 format.
	Output is 32 bits wide in Q23 format.

	Method: Polyfit coffecients are found using MATLAB. A memory is created to store those coefficients.

	Latency = 6
*/


module LOG_POLY(input clk, input reset, input [47:0] LogIn, output reg [30:0] LogOut);

reg [29:0] Log_C2[256];
reg [21:0] Log_C1[256];
reg [12:0] Log_C0[256];

reg [95:0] LogInSquare;
reg [125:0] Term1;
reg [69:0] Term2;
reg [26:0] Term3;

reg [23:0] FractionBit;
reg [6:0] IntegerBits;
reg [29:0] Log;

reg [47:0] LogIn2;
reg [125:0] Term11;
reg [69:0] Term21;
reg [26:0] Term31;
reg [22:0] LogPipe;

always @(posedge clk)
begin
	if(!reset)
	begin

		//CYCLE 1
		LogInSquare <= LogIn * LogIn;
		LogIn2 <= LogIn;

		//CYCLE 2		
		Term1 <= LogInSquare * Log_C2[LogIn2[47:40]];
		Term2 <= LogIn2 * Log_C1[LogIn2[47:40]];
		Term3 <= { Log_C0[LogIn2[47:40]], 14'b00000000_000000 };

		//CYCLE 3
		Term11 <= Term1;
		Term21 <= Term2;
		Term31 <= Term3;

		FractionBit <= Term1[111:89] - Term2[60:38] + Term3 [23:1];

		//CYCLE 4
		IntegerBits <=  Term11[118:112] - Term21[67:61] + Term31 [26:24] + FractionBit[23];
		LogPipe[22:0] <= FractionBit[22:0];

		//CYCLE 5
		Log[22:0] <= LogPipe[22:0];
		Log[29:23] <= IntegerBits[6:0];

		//CYCLE 6
		LogOut <= Log * 2;

	end

	else begin

		//LogOut <= 31'b0;

	// C2 Coefficient Table

		Log_C2[0] <= 30'b111111111111111111111111111111;
		Log_C2[1] <= 30'b111011110010100011100010001111;
		Log_C2[2] <= 30'b010100110101110010110001110101;
		Log_C2[3] <= 30'b001010100010101011001001011011;
		Log_C2[4] <= 30'b000110010110101101001111011101;
		Log_C2[5] <= 30'b000100001111110001101111110100;
		Log_C2[6] <= 30'b000011000010011000111000010010;
		Log_C2[7] <= 30'b000010010001111010100010101111;
		Log_C2[8] <= 30'b000001110001100011011001111100;
		Log_C2[9] <= 30'b000001011010111000001110000011;
		Log_C2[10] <= 30'b000001001010011000000101111001;
		Log_C2[11] <= 30'b000000111101111111100110010010;
		Log_C2[12] <= 30'b000000110100011101110000010101;
		Log_C2[13] <= 30'b000000101100111110011100110111;
		Log_C2[14] <= 30'b000000100110111110111010101110;
		Log_C2[15] <= 30'b000000100010000111001111001110;
		Log_C2[16] <= 30'b000000011110000110100001010100;
		Log_C2[17] <= 30'b000000011010110000100011111111;
		Log_C2[18] <= 30'b000000010111111100010111100010;
		Log_C2[19] <= 30'b000000010101100011001100000011;
		Log_C2[20] <= 30'b000000010011011111111000011011;
		Log_C2[21] <= 30'b000000010001101110011110010000;
		Log_C2[22] <= 30'b000000010000001011110110011101;
		Log_C2[23] <= 30'b000000001110110101100011010101;
		Log_C2[24] <= 30'b000000001101101001100110110010;
		Log_C2[25] <= 30'b000000001100100110011010111001;
		Log_C2[26] <= 30'b000000001011101010101100101001;
		Log_C2[27] <= 30'b000000001010110101010111110100;
		Log_C2[28] <= 30'b000000001010000101100011111100;
		Log_C2[29] <= 30'b000000001001011010100010000000;
		Log_C2[30] <= 30'b000000001000110011101010100001;
		Log_C2[31] <= 30'b000000001000010000011100001011;
		Log_C2[32] <= 30'b000000000111110000011010110000;
		Log_C2[33] <= 30'b000000000111010011001110000111;
		Log_C2[34] <= 30'b000000000110111000100001101000;
		Log_C2[35] <= 30'b000000000110100000000011011111;
		Log_C2[36] <= 30'b000000000110001001100100010101;
		Log_C2[37] <= 30'b000000000101110100110110110000;
		Log_C2[38] <= 30'b000000000101100001101111001001;
		Log_C2[39] <= 30'b000000000101010000000011010010;
		Log_C2[40] <= 30'b000000000100111111101010010000;
		Log_C2[41] <= 30'b000000000100110000011100001000;
		Log_C2[42] <= 30'b000000000100100010010001111101;
		Log_C2[43] <= 30'b000000000100010101000101100100;
		Log_C2[44] <= 30'b000000000100001000110001011110;
		Log_C2[45] <= 30'b000000000011111101010000110000;
		Log_C2[46] <= 30'b000000000011110010011111000100;
		Log_C2[47] <= 30'b000000000011101000011000011111;
		Log_C2[48] <= 30'b000000000011011110111001011110;
		Log_C2[49] <= 30'b000000000011010101111110111001;
		Log_C2[50] <= 30'b000000000011001101100101110111;
		Log_C2[51] <= 30'b000000000011000101101011110101;
		Log_C2[52] <= 30'b000000000010111110001110011011;
		Log_C2[53] <= 30'b000000000010110111001011100010;
		Log_C2[54] <= 30'b000000000010110000100001010000;
		Log_C2[55] <= 30'b000000000010101010001101110011;
		Log_C2[56] <= 30'b000000000010100100001111100101;
		Log_C2[57] <= 30'b000000000010011110100101001000;
		Log_C2[58] <= 30'b000000000010011001001101000110;
		Log_C2[59] <= 30'b000000000010010100000110010001;
		Log_C2[60] <= 30'b000000000010001111001111100001;
		Log_C2[61] <= 30'b000000000010001010100111110100;
		Log_C2[62] <= 30'b000000000010000110001110001011;
		Log_C2[63] <= 30'b000000000010000010000001101111;
		Log_C2[64] <= 30'b000000000001111110000001101100;
		Log_C2[65] <= 30'b000000000001111010001101010010;
		Log_C2[66] <= 30'b000000000001110110100011110101;
		Log_C2[67] <= 30'b000000000001110011000100101010;
		Log_C2[68] <= 30'b000000000001101111101111001101;
		Log_C2[69] <= 30'b000000000001101100100010111000;
		Log_C2[70] <= 30'b000000000001101001011111001101;
		Log_C2[71] <= 30'b000000000001100110100011101011;
		Log_C2[72] <= 30'b000000000001100011101111110110;
		Log_C2[73] <= 30'b000000000001100001000011010100;
		Log_C2[74] <= 30'b000000000001011110011101101100;
		Log_C2[75] <= 30'b000000000001011011111110100110;
		Log_C2[76] <= 30'b000000000001011001100101101101;
		Log_C2[77] <= 30'b000000000001010111010010101100;
		Log_C2[78] <= 30'b000000000001010101000101010000;
		Log_C2[79] <= 30'b000000000001010010111101001000;
		Log_C2[80] <= 30'b000000000001010000111010000011;
		Log_C2[81] <= 30'b000000000001001110111011110000;
		Log_C2[82] <= 30'b000000000001001101000010000001;
		Log_C2[83] <= 30'b000000000001001011001100101001;
		Log_C2[84] <= 30'b000000000001001001011011011010;
		Log_C2[85] <= 30'b000000000001000111101110001000;
		Log_C2[86] <= 30'b000000000001000110000100100111;
		Log_C2[87] <= 30'b000000000001000100011110101100;
		Log_C2[88] <= 30'b000000000001000010111100001101;
		Log_C2[89] <= 30'b000000000001000001011101000000;
		Log_C2[90] <= 30'b000000000001000000000000111011;
		Log_C2[91] <= 30'b000000000000111110100111110111;
		Log_C2[92] <= 30'b000000000000111101010001101011;
		Log_C2[93] <= 30'b000000000000111011111110001111;
		Log_C2[94] <= 30'b000000000000111010101101011100;
		Log_C2[95] <= 30'b000000000000111001011111001010;
		Log_C2[96] <= 30'b000000000000111000010011010011;
		Log_C2[97] <= 30'b000000000000110111001001110001;
		Log_C2[98] <= 30'b000000000000110110000010011101;
		Log_C2[99] <= 30'b000000000000110100111101010010;
		Log_C2[100] <= 30'b000000000000110011111010001011;
		Log_C2[101] <= 30'b000000000000110010111001000010;
		Log_C2[102] <= 30'b000000000000110001111001110011;
		Log_C2[103] <= 30'b000000000000110000111100011000;
		Log_C2[104] <= 30'b000000000000110000000000101101;
		Log_C2[105] <= 30'b000000000000101111000110101111;
		Log_C2[106] <= 30'b000000000000101110001110011001;
		Log_C2[107] <= 30'b000000000000101101010111100110;
		Log_C2[108] <= 30'b000000000000101100100010010101;
		Log_C2[109] <= 30'b000000000000101011101110100000;
		Log_C2[110] <= 30'b000000000000101010111100000101;
		Log_C2[111] <= 30'b000000000000101010001011000000;
		Log_C2[112] <= 30'b000000000000101001011011001111;
		Log_C2[113] <= 30'b000000000000101000101100101110;
		Log_C2[114] <= 30'b000000000000100111111111011011;
		Log_C2[115] <= 30'b000000000000100111010011010011;
		Log_C2[116] <= 30'b000000000000100110101000010011;
		Log_C2[117] <= 30'b000000000000100101111110011010;
		Log_C2[118] <= 30'b000000000000100101010101100011;
		Log_C2[119] <= 30'b000000000000100100101101101111;
		Log_C2[120] <= 30'b000000000000100100000110111001;
		Log_C2[121] <= 30'b000000000000100011100001000000;
		Log_C2[122] <= 30'b000000000000100010111100000011;
		Log_C2[123] <= 30'b000000000000100010010111111111;
		Log_C2[124] <= 30'b000000000000100001110100110010;
		Log_C2[125] <= 30'b000000000000100001010010011011;
		Log_C2[126] <= 30'b000000000000100000110000111000;
		Log_C2[127] <= 30'b000000000000100000010000000111;
		Log_C2[128] <= 30'b000000000000011111110000000111;
		Log_C2[129] <= 30'b000000000000011111010000110110;
		Log_C2[130] <= 30'b000000000000011110110010010011;
		Log_C2[131] <= 30'b000000000000011110010100011100;
		Log_C2[132] <= 30'b000000000000011101110111010001;
		Log_C2[133] <= 30'b000000000000011101011010101111;
		Log_C2[134] <= 30'b000000000000011100111110110110;
		Log_C2[135] <= 30'b000000000000011100100011100100;
		Log_C2[136] <= 30'b000000000000011100001000111001;
		Log_C2[137] <= 30'b000000000000011011101110110011;
		Log_C2[138] <= 30'b000000000000011011010101010000;
		Log_C2[139] <= 30'b000000000000011010111100010001;
		Log_C2[140] <= 30'b000000000000011010100011110100;
		Log_C2[141] <= 30'b000000000000011010001011110111;
		Log_C2[142] <= 30'b000000000000011001110100011011;
		Log_C2[143] <= 30'b000000000000011001011101011111;
		Log_C2[144] <= 30'b000000000000011001000111000000;
		Log_C2[145] <= 30'b000000000000011000110000111111;
		Log_C2[146] <= 30'b000000000000011000011011011011;
		Log_C2[147] <= 30'b000000000000011000000110010011;
		Log_C2[148] <= 30'b000000000000010111110001100110;
		Log_C2[149] <= 30'b000000000000010111011101010100;
		Log_C2[150] <= 30'b000000000000010111001001011011;
		Log_C2[151] <= 30'b000000000000010110110101111100;
		Log_C2[152] <= 30'b000000000000010110100010110100;
		Log_C2[153] <= 30'b000000000000010110010000000101;
		Log_C2[154] <= 30'b000000000000010101111101101101;
		Log_C2[155] <= 30'b000000000000010101101011101100;
		Log_C2[156] <= 30'b000000000000010101011010000001;
		Log_C2[157] <= 30'b000000000000010101001000101011;
		Log_C2[158] <= 30'b000000000000010100110111101010;
		Log_C2[159] <= 30'b000000000000010100100110111101;
		Log_C2[160] <= 30'b000000000000010100010110100101;
		Log_C2[161] <= 30'b000000000000010100000110011111;
		Log_C2[162] <= 30'b000000000000010011110110101101;
		Log_C2[163] <= 30'b000000000000010011100111001101;
		Log_C2[164] <= 30'b000000000000010011011000000000;
		Log_C2[165] <= 30'b000000000000010011001001000100;
		Log_C2[166] <= 30'b000000000000010010111010011001;
		Log_C2[167] <= 30'b000000000000010010101011111110;
		Log_C2[168] <= 30'b000000000000010010011101110101;
		Log_C2[169] <= 30'b000000000000010010001111111011;
		Log_C2[170] <= 30'b000000000000010010000010010000;
		Log_C2[171] <= 30'b000000000000010001110100110110;
		Log_C2[172] <= 30'b000000000000010001100111101001;
		Log_C2[173] <= 30'b000000000000010001011010101100;
		Log_C2[174] <= 30'b000000000000010001001101111101;
		Log_C2[175] <= 30'b000000000000010001000001011011;
		Log_C2[176] <= 30'b000000000000010000110101000111;
		Log_C2[177] <= 30'b000000000000010000101001000001;
		Log_C2[178] <= 30'b000000000000010000011101000111;
		Log_C2[179] <= 30'b000000000000010000010001011010;
		Log_C2[180] <= 30'b000000000000010000000101111010;
		Log_C2[181] <= 30'b000000000000001111111010100110;
		Log_C2[182] <= 30'b000000000000001111101111011101;
		Log_C2[183] <= 30'b000000000000001111100100100000;
		Log_C2[184] <= 30'b000000000000001111011001101111;
		Log_C2[185] <= 30'b000000000000001111001111001000;
		Log_C2[186] <= 30'b000000000000001111000100101101;
		Log_C2[187] <= 30'b000000000000001110111010011100;
		Log_C2[188] <= 30'b000000000000001110110000010110;
		Log_C2[189] <= 30'b000000000000001110100110011010;
		Log_C2[190] <= 30'b000000000000001110011100100111;
		Log_C2[191] <= 30'b000000000000001110010010111111;
		Log_C2[192] <= 30'b000000000000001110001001100000;
		Log_C2[193] <= 30'b000000000000001110000000001011;
		Log_C2[194] <= 30'b000000000000001101110110111110;
		Log_C2[195] <= 30'b000000000000001101101101111011;
		Log_C2[196] <= 30'b000000000000001101100101000001;
		Log_C2[197] <= 30'b000000000000001101011100001111;
		Log_C2[198] <= 30'b000000000000001101010011100110;
		Log_C2[199] <= 30'b000000000000001101001011000101;
		Log_C2[200] <= 30'b000000000000001101000010101100;
		Log_C2[201] <= 30'b000000000000001100111010011011;
		Log_C2[202] <= 30'b000000000000001100110010010010;
		Log_C2[203] <= 30'b000000000000001100101010010000;
		Log_C2[204] <= 30'b000000000000001100100010010110;
		Log_C2[205] <= 30'b000000000000001100011010100100;
		Log_C2[206] <= 30'b000000000000001100010010111001;
		Log_C2[207] <= 30'b000000000000001100001011010100;
		Log_C2[208] <= 30'b000000000000001100000011110111;
		Log_C2[209] <= 30'b000000000000001011111100100001;
		Log_C2[210] <= 30'b000000000000001011110101010001;
		Log_C2[211] <= 30'b000000000000001011101110001000;
		Log_C2[212] <= 30'b000000000000001011100111000101;
		Log_C2[213] <= 30'b000000000000001011100000001000;
		Log_C2[214] <= 30'b000000000000001011011001010010;
		Log_C2[215] <= 30'b000000000000001011010010100010;
		Log_C2[216] <= 30'b000000000000001011001011111000;
		Log_C2[217] <= 30'b000000000000001011000101010011;
		Log_C2[218] <= 30'b000000000000001010111110110101;
		Log_C2[219] <= 30'b000000000000001010111000011100;
		Log_C2[220] <= 30'b000000000000001010110010001001;
		Log_C2[221] <= 30'b000000000000001010101011111011;
		Log_C2[222] <= 30'b000000000000001010100101110010;
		Log_C2[223] <= 30'b000000000000001010011111101111;
		Log_C2[224] <= 30'b000000000000001010011001110001;
		Log_C2[225] <= 30'b000000000000001010010011111000;
		Log_C2[226] <= 30'b000000000000001010001110000100;
		Log_C2[227] <= 30'b000000000000001010001000010100;
		Log_C2[228] <= 30'b000000000000001010000010101010;
		Log_C2[229] <= 30'b000000000000001001111101000100;
		Log_C2[230] <= 30'b000000000000001001110111100011;
		Log_C2[231] <= 30'b000000000000001001110010000111;
		Log_C2[232] <= 30'b000000000000001001101100101111;
		Log_C2[233] <= 30'b000000000000001001100111011011;
		Log_C2[234] <= 30'b000000000000001001100010001100;
		Log_C2[235] <= 30'b000000000000001001011101000001;
		Log_C2[236] <= 30'b000000000000001001010111111010;
		Log_C2[237] <= 30'b000000000000001001010010111000;
		Log_C2[238] <= 30'b000000000000001001001101111001;
		Log_C2[239] <= 30'b000000000000001001001000111111;
		Log_C2[240] <= 30'b000000000000001001000100001000;
		Log_C2[241] <= 30'b000000000000001000111111010101;
		Log_C2[242] <= 30'b000000000000001000111010100110;
		Log_C2[243] <= 30'b000000000000001000110101111011;
		Log_C2[244] <= 30'b000000000000001000110001010011;
		Log_C2[245] <= 30'b000000000000001000101100101111;
		Log_C2[246] <= 30'b000000000000001000101000001110;
		Log_C2[247] <= 30'b000000000000001000100011110001;
		Log_C2[248] <= 30'b000000000000001000011111011000;
		Log_C2[249] <= 30'b000000000000001000011011000010;
		Log_C2[250] <= 30'b000000000000001000010110101111;
		Log_C2[251] <= 30'b000000000000001000010010011111;
		Log_C2[252] <= 30'b000000000000001000001110010011;
		Log_C2[253] <= 30'b000000000000001000001010001010;
		Log_C2[254] <= 30'b000000000000001000000110000011;
		Log_C2[255] <= 30'b000000000000001000000010000000;


	// C1 Coefficient Table

		Log_C1[0] <= 22'b1111111111111111111111;
		Log_C1[1] <= 22'b1011000100000100110111;
		Log_C1[2] <= 22'b0110011110111000010000;
		Log_C1[3] <= 22'b0100100110011110011011;
		Log_C1[4] <= 22'b0011100100011100101001;
		Log_C1[5] <= 22'b0010111010101010110110;
		Log_C1[6] <= 22'b0010011101110101010110;
		Log_C1[7] <= 22'b0010001000101110011011;
		Log_C1[8] <= 22'b0001111000100110100011;
		Log_C1[9] <= 22'b0001101011111000100100;
		Log_C1[10] <= 22'b0001100001100110000000;
		Log_C1[11] <= 22'b0001011001000110001100;
		Log_C1[12] <= 22'b0001010001111101100010;
		Log_C1[13] <= 22'b0001001011111000101000;
		Log_C1[14] <= 22'b0001000110101001011011;
		Log_C1[15] <= 22'b0001000010000101100001;
		Log_C1[16] <= 22'b0000111110000101000010;
		Log_C1[17] <= 22'b0000111010100001111000;
		Log_C1[18] <= 22'b0000110111010111010011;
		Log_C1[19] <= 22'b0000110100100001100001;
		Log_C1[20] <= 22'b0000110001111101011111;
		Log_C1[21] <= 22'b0000101111101000101101;
		Log_C1[22] <= 22'b0000101101100001001011;
		Log_C1[23] <= 22'b0000101011100101001011;
		Log_C1[24] <= 22'b0000101001110011010011;
		Log_C1[25] <= 22'b0000101000001010010110;
		Log_C1[26] <= 22'b0000100110101001010101;
		Log_C1[27] <= 22'b0000100101001111011000;
		Log_C1[28] <= 22'b0000100011111011101111;
		Log_C1[29] <= 22'b0000100010101101110001;
		Log_C1[30] <= 22'b0000100001100100111010;
		Log_C1[31] <= 22'b0000100000100000101011;
		Log_C1[32] <= 22'b0000011111100000101001;
		Log_C1[33] <= 22'b0000011110100100011100;
		Log_C1[34] <= 22'b0000011101101011101110;
		Log_C1[35] <= 22'b0000011100110110001101;
		Log_C1[36] <= 22'b0000011100000011100111;
		Log_C1[37] <= 22'b0000011011010011101110;
		Log_C1[38] <= 22'b0000011010100110010101;
		Log_C1[39] <= 22'b0000011001111011001110;
		Log_C1[40] <= 22'b0000011001010010010000;
		Log_C1[41] <= 22'b0000011000101011010000;
		Log_C1[42] <= 22'b0000011000000110000110;
		Log_C1[43] <= 22'b0000010111100010101001;
		Log_C1[44] <= 22'b0000010111000000110010;
		Log_C1[45] <= 22'b0000010110100000011010;
		Log_C1[46] <= 22'b0000010110000001011011;
		Log_C1[47] <= 22'b0000010101100011110000;
		Log_C1[48] <= 22'b0000010101000111010011;
		Log_C1[49] <= 22'b0000010100101100000000;
		Log_C1[50] <= 22'b0000010100010001110010;
		Log_C1[51] <= 22'b0000010011111000100101;
		Log_C1[52] <= 22'b0000010011100000010110;
		Log_C1[53] <= 22'b0000010011001001000000;
		Log_C1[54] <= 22'b0000010010110010100010;
		Log_C1[55] <= 22'b0000010010011100110111;
		Log_C1[56] <= 22'b0000010010000111111101;
		Log_C1[57] <= 22'b0000010001110011110010;
		Log_C1[58] <= 22'b0000010001100000010011;
		Log_C1[59] <= 22'b0000010001001101011110;
		Log_C1[60] <= 22'b0000010000111011010001;
		Log_C1[61] <= 22'b0000010000101001101001;
		Log_C1[62] <= 22'b0000010000011000100110;
		Log_C1[63] <= 22'b0000010000001000000101;
		Log_C1[64] <= 22'b0000001111111000000101;
		Log_C1[65] <= 22'b0000001111101000100100;
		Log_C1[66] <= 22'b0000001111011001100001;
		Log_C1[67] <= 22'b0000001111001010111011;
		Log_C1[68] <= 22'b0000001110111100110000;
		Log_C1[69] <= 22'b0000001110101110111111;
		Log_C1[70] <= 22'b0000001110100001100111;
		Log_C1[71] <= 22'b0000001110010100100110;
		Log_C1[72] <= 22'b0000001110000111111101;
		Log_C1[73] <= 22'b0000001101111011101010;
		Log_C1[74] <= 22'b0000001101101111101100;
		Log_C1[75] <= 22'b0000001101100100000010;
		Log_C1[76] <= 22'b0000001101011000101100;
		Log_C1[77] <= 22'b0000001101001101101001;
		Log_C1[78] <= 22'b0000001101000010110111;
		Log_C1[79] <= 22'b0000001100111000010111;
		Log_C1[80] <= 22'b0000001100101110001000;
		Log_C1[81] <= 22'b0000001100100100001000;
		Log_C1[82] <= 22'b0000001100011010011001;
		Log_C1[83] <= 22'b0000001100010000111000;
		Log_C1[84] <= 22'b0000001100000111100101;
		Log_C1[85] <= 22'b0000001011111110100001;
		Log_C1[86] <= 22'b0000001011110101101010;
		Log_C1[87] <= 22'b0000001011101100111111;
		Log_C1[88] <= 22'b0000001011100100100010;
		Log_C1[89] <= 22'b0000001011011100010000;
		Log_C1[90] <= 22'b0000001011010100001010;
		Log_C1[91] <= 22'b0000001011001100010000;
		Log_C1[92] <= 22'b0000001011000100100000;
		Log_C1[93] <= 22'b0000001010111100111011;
		Log_C1[94] <= 22'b0000001010110101100001;
		Log_C1[95] <= 22'b0000001010101110010000;
		Log_C1[96] <= 22'b0000001010100111001001;
		Log_C1[97] <= 22'b0000001010100000001011;
		Log_C1[98] <= 22'b0000001010011001010110;
		Log_C1[99] <= 22'b0000001010010010101010;
		Log_C1[100] <= 22'b0000001010001100000111;
		Log_C1[101] <= 22'b0000001010000101101100;
		Log_C1[102] <= 22'b0000001001111111011000;
		Log_C1[103] <= 22'b0000001001111001001101;
		Log_C1[104] <= 22'b0000001001110011001001;
		Log_C1[105] <= 22'b0000001001101101001101;
		Log_C1[106] <= 22'b0000001001100111010111;
		Log_C1[107] <= 22'b0000001001100001101001;
		Log_C1[108] <= 22'b0000001001011100000001;
		Log_C1[109] <= 22'b0000001001010110100000;
		Log_C1[110] <= 22'b0000001001010001000110;
		Log_C1[111] <= 22'b0000001001001011110001;
		Log_C1[112] <= 22'b0000001001000110100011;
		Log_C1[113] <= 22'b0000001001000001011010;
		Log_C1[114] <= 22'b0000001000111100011000;
		Log_C1[115] <= 22'b0000001000110111011011;
		Log_C1[116] <= 22'b0000001000110010100011;
		Log_C1[117] <= 22'b0000001000101101110000;
		Log_C1[118] <= 22'b0000001000101001000011;
		Log_C1[119] <= 22'b0000001000100100011011;
		Log_C1[120] <= 22'b0000001000011111111000;
		Log_C1[121] <= 22'b0000001000011011011001;
		Log_C1[122] <= 22'b0000001000010110111111;
		Log_C1[123] <= 22'b0000001000010010101010;
		Log_C1[124] <= 22'b0000001000001110011001;
		Log_C1[125] <= 22'b0000001000001010001101;
		Log_C1[126] <= 22'b0000001000000110000101;
		Log_C1[127] <= 22'b0000001000000010000001;
		Log_C1[128] <= 22'b0000000111111110000001;
		Log_C1[129] <= 22'b0000000111111010000101;
		Log_C1[130] <= 22'b0000000111110110001100;
		Log_C1[131] <= 22'b0000000111110010011000;
		Log_C1[132] <= 22'b0000000111101110100111;
		Log_C1[133] <= 22'b0000000111101010111010;
		Log_C1[134] <= 22'b0000000111100111010001;
		Log_C1[135] <= 22'b0000000111100011101010;
		Log_C1[136] <= 22'b0000000111100000001000;
		Log_C1[137] <= 22'b0000000111011100101000;
		Log_C1[138] <= 22'b0000000111011001001100;
		Log_C1[139] <= 22'b0000000111010101110011;
		Log_C1[140] <= 22'b0000000111010010011101;
		Log_C1[141] <= 22'b0000000111001111001010;
		Log_C1[142] <= 22'b0000000111001011111010;
		Log_C1[143] <= 22'b0000000111001000101101;
		Log_C1[144] <= 22'b0000000111000101100010;
		Log_C1[145] <= 22'b0000000111000010011011;
		Log_C1[146] <= 22'b0000000110111111010110;
		Log_C1[147] <= 22'b0000000110111100010100;
		Log_C1[148] <= 22'b0000000110111001010101;
		Log_C1[149] <= 22'b0000000110110110011000;
		Log_C1[150] <= 22'b0000000110110011011101;
		Log_C1[151] <= 22'b0000000110110000100101;
		Log_C1[152] <= 22'b0000000110101101110000;
		Log_C1[153] <= 22'b0000000110101010111101;
		Log_C1[154] <= 22'b0000000110101000001100;
		Log_C1[155] <= 22'b0000000110100101011101;
		Log_C1[156] <= 22'b0000000110100010110001;
		Log_C1[157] <= 22'b0000000110100000000111;
		Log_C1[158] <= 22'b0000000110011101011111;
		Log_C1[159] <= 22'b0000000110011010111001;
		Log_C1[160] <= 22'b0000000110011000010101;
		Log_C1[161] <= 22'b0000000110010101110011;
		Log_C1[162] <= 22'b0000000110010011010011;
		Log_C1[163] <= 22'b0000000110010000110101;
		Log_C1[164] <= 22'b0000000110001110011001;
		Log_C1[165] <= 22'b0000000110001011111111;
		Log_C1[166] <= 22'b0000000110001001100111;
		Log_C1[167] <= 22'b0000000110000111010001;
		Log_C1[168] <= 22'b0000000110000100111100;
		Log_C1[169] <= 22'b0000000110000010101001;
		Log_C1[170] <= 22'b0000000110000000011000;
		Log_C1[171] <= 22'b0000000101111110001001;
		Log_C1[172] <= 22'b0000000101111011111011;
		Log_C1[173] <= 22'b0000000101111001101111;
		Log_C1[174] <= 22'b0000000101110111100100;
		Log_C1[175] <= 22'b0000000101110101011011;
		Log_C1[176] <= 22'b0000000101110011010100;
		Log_C1[177] <= 22'b0000000101110001001110;
		Log_C1[178] <= 22'b0000000101101111001010;
		Log_C1[179] <= 22'b0000000101101101000111;
		Log_C1[180] <= 22'b0000000101101011000101;
		Log_C1[181] <= 22'b0000000101101001000101;
		Log_C1[182] <= 22'b0000000101100111000111;
		Log_C1[183] <= 22'b0000000101100101001001;
		Log_C1[184] <= 22'b0000000101100011001101;
		Log_C1[185] <= 22'b0000000101100001010011;
		Log_C1[186] <= 22'b0000000101011111011010;
		Log_C1[187] <= 22'b0000000101011101100010;
		Log_C1[188] <= 22'b0000000101011011101011;
		Log_C1[189] <= 22'b0000000101011001110110;
		Log_C1[190] <= 22'b0000000101011000000001;
		Log_C1[191] <= 22'b0000000101010110001110;
		Log_C1[192] <= 22'b0000000101010100011101;
		Log_C1[193] <= 22'b0000000101010010101100;
		Log_C1[194] <= 22'b0000000101010000111101;
		Log_C1[195] <= 22'b0000000101001111001110;
		Log_C1[196] <= 22'b0000000101001101100001;
		Log_C1[197] <= 22'b0000000101001011110101;
		Log_C1[198] <= 22'b0000000101001010001010;
		Log_C1[199] <= 22'b0000000101001000100000;
		Log_C1[200] <= 22'b0000000101000110110111;
		Log_C1[201] <= 22'b0000000101000101001111;
		Log_C1[202] <= 22'b0000000101000011101001;
		Log_C1[203] <= 22'b0000000101000010000011;
		Log_C1[204] <= 22'b0000000101000000011110;
		Log_C1[205] <= 22'b0000000100111110111010;
		Log_C1[206] <= 22'b0000000100111101010111;
		Log_C1[207] <= 22'b0000000100111011110110;
		Log_C1[208] <= 22'b0000000100111010010101;
		Log_C1[209] <= 22'b0000000100111000110101;
		Log_C1[210] <= 22'b0000000100110111010101;
		Log_C1[211] <= 22'b0000000100110101110111;
		Log_C1[212] <= 22'b0000000100110100011010;
		Log_C1[213] <= 22'b0000000100110010111101;
		Log_C1[214] <= 22'b0000000100110001100010;
		Log_C1[215] <= 22'b0000000100110000000111;
		Log_C1[216] <= 22'b0000000100101110101101;
		Log_C1[217] <= 22'b0000000100101101010100;
		Log_C1[218] <= 22'b0000000100101011111100;
		Log_C1[219] <= 22'b0000000100101010100100;
		Log_C1[220] <= 22'b0000000100101001001110;
		Log_C1[221] <= 22'b0000000100100111111000;
		Log_C1[222] <= 22'b0000000100100110100011;
		Log_C1[223] <= 22'b0000000100100101001110;
		Log_C1[224] <= 22'b0000000100100011111011;
		Log_C1[225] <= 22'b0000000100100010101000;
		Log_C1[226] <= 22'b0000000100100001010110;
		Log_C1[227] <= 22'b0000000100100000000101;
		Log_C1[228] <= 22'b0000000100011110110100;
		Log_C1[229] <= 22'b0000000100011101100100;
		Log_C1[230] <= 22'b0000000100011100010101;
		Log_C1[231] <= 22'b0000000100011011000110;
		Log_C1[232] <= 22'b0000000100011001111000;
		Log_C1[233] <= 22'b0000000100011000101011;
		Log_C1[234] <= 22'b0000000100010111011110;
		Log_C1[235] <= 22'b0000000100010110010010;
		Log_C1[236] <= 22'b0000000100010101000111;
		Log_C1[237] <= 22'b0000000100010011111100;
		Log_C1[238] <= 22'b0000000100010010110010;
		Log_C1[239] <= 22'b0000000100010001101001;
		Log_C1[240] <= 22'b0000000100010000100000;
		Log_C1[241] <= 22'b0000000100001111011000;
		Log_C1[242] <= 22'b0000000100001110010000;
		Log_C1[243] <= 22'b0000000100001101001001;
		Log_C1[244] <= 22'b0000000100001100000011;
		Log_C1[245] <= 22'b0000000100001010111101;
		Log_C1[246] <= 22'b0000000100001001110111;
		Log_C1[247] <= 22'b0000000100001000110011;
		Log_C1[248] <= 22'b0000000100000111101111;
		Log_C1[249] <= 22'b0000000100000110101011;
		Log_C1[250] <= 22'b0000000100000101101000;
		Log_C1[251] <= 22'b0000000100000100100101;
		Log_C1[252] <= 22'b0000000100000011100011;
		Log_C1[253] <= 22'b0000000100000010100010;
		Log_C1[254] <= 22'b0000000100000001100001;
		Log_C1[255] <= 22'b0000000100000000100000;

	// C0 Coefficient Table
		Log_C0[0] <= 13'b1111111111111;
		Log_C0[1] <= 13'b1101011000001;
		Log_C0[2] <= 13'b1100010010101;
		Log_C0[3] <= 13'b1011100110100;
		Log_C0[4] <= 13'b1011000101111;
		Log_C0[5] <= 13'b1010101100000;
		Log_C0[6] <= 13'b1010010110100;
		Log_C0[7] <= 13'b1010000100001;
		Log_C0[8] <= 13'b1001110100000;
		Log_C0[9] <= 13'b1001100101110;
		Log_C0[10] <= 13'b1001011000111;
		Log_C0[11] <= 13'b1001001101010;
		Log_C0[12] <= 13'b1001000010101;
		Log_C0[13] <= 13'b1000111000110;
		Log_C0[14] <= 13'b1000101111100;
		Log_C0[15] <= 13'b1000100111000;
		Log_C0[16] <= 13'b1000011111000;
		Log_C0[17] <= 13'b1000010111100;
		Log_C0[18] <= 13'b1000010000011;
		Log_C0[19] <= 13'b1000001001101;
		Log_C0[20] <= 13'b1000000011010;
		Log_C0[21] <= 13'b0111111101001;
		Log_C0[22] <= 13'b0111110111010;
		Log_C0[23] <= 13'b0111110001110;
		Log_C0[24] <= 13'b0111101100011;
		Log_C0[25] <= 13'b0111100111010;
		Log_C0[26] <= 13'b0111100010011;
		Log_C0[27] <= 13'b0111011101101;
		Log_C0[28] <= 13'b0111011001000;
		Log_C0[29] <= 13'b0111010100101;
		Log_C0[30] <= 13'b0111010000011;
		Log_C0[31] <= 13'b0111001100010;
		Log_C0[32] <= 13'b0111001000010;
		Log_C0[33] <= 13'b0111000100011;
		Log_C0[34] <= 13'b0111000000100;
		Log_C0[35] <= 13'b0110111100111;
		Log_C0[36] <= 13'b0110111001011;
		Log_C0[37] <= 13'b0110110101111;
		Log_C0[38] <= 13'b0110110010100;
		Log_C0[39] <= 13'b0110101111010;
		Log_C0[40] <= 13'b0110101100000;
		Log_C0[41] <= 13'b0110101000111;
		Log_C0[42] <= 13'b0110100101111;
		Log_C0[43] <= 13'b0110100010111;
		Log_C0[44] <= 13'b0110100000000;
		Log_C0[45] <= 13'b0110011101001;
		Log_C0[46] <= 13'b0110011010011;
		Log_C0[47] <= 13'b0110010111101;
		Log_C0[48] <= 13'b0110010101000;
		Log_C0[49] <= 13'b0110010010011;
		Log_C0[50] <= 13'b0110001111110;
		Log_C0[51] <= 13'b0110001101010;
		Log_C0[52] <= 13'b0110001010110;
		Log_C0[53] <= 13'b0110001000011;
		Log_C0[54] <= 13'b0110000110000;
		Log_C0[55] <= 13'b0110000011110;
		Log_C0[56] <= 13'b0110000001011;
		Log_C0[57] <= 13'b0101111111001;
		Log_C0[58] <= 13'b0101111101000;
		Log_C0[59] <= 13'b0101111010110;
		Log_C0[60] <= 13'b0101111000101;
		Log_C0[61] <= 13'b0101110110100;
		Log_C0[62] <= 13'b0101110100100;
		Log_C0[63] <= 13'b0101110010100;
		Log_C0[64] <= 13'b0101110000100;
		Log_C0[65] <= 13'b0101101110100;
		Log_C0[66] <= 13'b0101101100100;
		Log_C0[67] <= 13'b0101101010101;
		Log_C0[68] <= 13'b0101101000110;
		Log_C0[69] <= 13'b0101100110111;
		Log_C0[70] <= 13'b0101100101001;
		Log_C0[71] <= 13'b0101100011010;
		Log_C0[72] <= 13'b0101100001100;
		Log_C0[73] <= 13'b0101011111110;
		Log_C0[74] <= 13'b0101011110000;
		Log_C0[75] <= 13'b0101011100010;
		Log_C0[76] <= 13'b0101011010101;
		Log_C0[77] <= 13'b0101011001000;
		Log_C0[78] <= 13'b0101010111010;
		Log_C0[79] <= 13'b0101010101110;
		Log_C0[80] <= 13'b0101010100001;
		Log_C0[81] <= 13'b0101010010100;
		Log_C0[82] <= 13'b0101010001000;
		Log_C0[83] <= 13'b0101001111011;
		Log_C0[84] <= 13'b0101001101111;
		Log_C0[85] <= 13'b0101001100011;
		Log_C0[86] <= 13'b0101001010111;
		Log_C0[87] <= 13'b0101001001011;
		Log_C0[88] <= 13'b0101001000000;
		Log_C0[89] <= 13'b0101000110100;
		Log_C0[90] <= 13'b0101000101001;
		Log_C0[91] <= 13'b0101000011110;
		Log_C0[92] <= 13'b0101000010010;
		Log_C0[93] <= 13'b0101000000111;
		Log_C0[94] <= 13'b0100111111101;
		Log_C0[95] <= 13'b0100111110010;
		Log_C0[96] <= 13'b0100111100111;
		Log_C0[97] <= 13'b0100111011101;
		Log_C0[98] <= 13'b0100111010010;
		Log_C0[99] <= 13'b0100111001000;
		Log_C0[100] <= 13'b0100110111101;
		Log_C0[101] <= 13'b0100110110011;
		Log_C0[102] <= 13'b0100110101001;
		Log_C0[103] <= 13'b0100110011111;
		Log_C0[104] <= 13'b0100110010110;
		Log_C0[105] <= 13'b0100110001100;
		Log_C0[106] <= 13'b0100110000010;
		Log_C0[107] <= 13'b0100101111001;
		Log_C0[108] <= 13'b0100101101111;
		Log_C0[109] <= 13'b0100101100110;
		Log_C0[110] <= 13'b0100101011100;
		Log_C0[111] <= 13'b0100101010011;
		Log_C0[112] <= 13'b0100101001010;
		Log_C0[113] <= 13'b0100101000001;
		Log_C0[114] <= 13'b0100100111000;
		Log_C0[115] <= 13'b0100100101111;
		Log_C0[116] <= 13'b0100100100110;
		Log_C0[117] <= 13'b0100100011101;
		Log_C0[118] <= 13'b0100100010101;
		Log_C0[119] <= 13'b0100100001100;
		Log_C0[120] <= 13'b0100100000100;
		Log_C0[121] <= 13'b0100011111011;
		Log_C0[122] <= 13'b0100011110011;
		Log_C0[123] <= 13'b0100011101010;
		Log_C0[124] <= 13'b0100011100010;
		Log_C0[125] <= 13'b0100011011010;
		Log_C0[126] <= 13'b0100011010010;
		Log_C0[127] <= 13'b0100011001010;
		Log_C0[128] <= 13'b0100011000010;
		Log_C0[129] <= 13'b0100010111010;
		Log_C0[130] <= 13'b0100010110010;
		Log_C0[131] <= 13'b0100010101010;
		Log_C0[132] <= 13'b0100010100010;
		Log_C0[133] <= 13'b0100010011011;
		Log_C0[134] <= 13'b0100010010011;
		Log_C0[135] <= 13'b0100010001011;
		Log_C0[136] <= 13'b0100010000100;
		Log_C0[137] <= 13'b0100001111100;
		Log_C0[138] <= 13'b0100001110101;
		Log_C0[139] <= 13'b0100001101110;
		Log_C0[140] <= 13'b0100001100110;
		Log_C0[141] <= 13'b0100001011111;
		Log_C0[142] <= 13'b0100001011000;
		Log_C0[143] <= 13'b0100001010001;
		Log_C0[144] <= 13'b0100001001010;
		Log_C0[145] <= 13'b0100001000011;
		Log_C0[146] <= 13'b0100000111100;
		Log_C0[147] <= 13'b0100000110101;
		Log_C0[148] <= 13'b0100000101110;
		Log_C0[149] <= 13'b0100000100111;
		Log_C0[150] <= 13'b0100000100000;
		Log_C0[151] <= 13'b0100000011001;
		Log_C0[152] <= 13'b0100000010010;
		Log_C0[153] <= 13'b0100000001100;
		Log_C0[154] <= 13'b0100000000101;
		Log_C0[155] <= 13'b0011111111111;
		Log_C0[156] <= 13'b0011111111000;
		Log_C0[157] <= 13'b0011111110001;
		Log_C0[158] <= 13'b0011111101011;
		Log_C0[159] <= 13'b0011111100100;
		Log_C0[160] <= 13'b0011111011110;
		Log_C0[161] <= 13'b0011111011000;
		Log_C0[162] <= 13'b0011111010001;
		Log_C0[163] <= 13'b0011111001011;
		Log_C0[164] <= 13'b0011111000101;
		Log_C0[165] <= 13'b0011110111111;
		Log_C0[166] <= 13'b0011110111001;
		Log_C0[167] <= 13'b0011110110010;
		Log_C0[168] <= 13'b0011110101100;
		Log_C0[169] <= 13'b0011110100110;
		Log_C0[170] <= 13'b0011110100000;
		Log_C0[171] <= 13'b0011110011010;
		Log_C0[172] <= 13'b0011110010100;
		Log_C0[173] <= 13'b0011110001110;
		Log_C0[174] <= 13'b0011110001000;
		Log_C0[175] <= 13'b0011110000011;
		Log_C0[176] <= 13'b0011101111101;
		Log_C0[177] <= 13'b0011101110111;
		Log_C0[178] <= 13'b0011101110001;
		Log_C0[179] <= 13'b0011101101100;
		Log_C0[180] <= 13'b0011101100110;
		Log_C0[181] <= 13'b0011101100000;
		Log_C0[182] <= 13'b0011101011011;
		Log_C0[183] <= 13'b0011101010101;
		Log_C0[184] <= 13'b0011101001111;
		Log_C0[185] <= 13'b0011101001010;
		Log_C0[186] <= 13'b0011101000100;
		Log_C0[187] <= 13'b0011100111111;
		Log_C0[188] <= 13'b0011100111001;
		Log_C0[189] <= 13'b0011100110100;
		Log_C0[190] <= 13'b0011100101111;
		Log_C0[191] <= 13'b0011100101001;
		Log_C0[192] <= 13'b0011100100100;
		Log_C0[193] <= 13'b0011100011111;
		Log_C0[194] <= 13'b0011100011001;
		Log_C0[195] <= 13'b0011100010100;
		Log_C0[196] <= 13'b0011100001111;
		Log_C0[197] <= 13'b0011100001010;
		Log_C0[198] <= 13'b0011100000100;
		Log_C0[199] <= 13'b0011011111111;
		Log_C0[200] <= 13'b0011011111010;
		Log_C0[201] <= 13'b0011011110101;
		Log_C0[202] <= 13'b0011011110000;
		Log_C0[203] <= 13'b0011011101011;
		Log_C0[204] <= 13'b0011011100110;
		Log_C0[205] <= 13'b0011011100001;
		Log_C0[206] <= 13'b0011011011100;
		Log_C0[207] <= 13'b0011011010111;
		Log_C0[208] <= 13'b0011011010010;
		Log_C0[209] <= 13'b0011011001101;
		Log_C0[210] <= 13'b0011011001000;
		Log_C0[211] <= 13'b0011011000100;
		Log_C0[212] <= 13'b0011010111111;
		Log_C0[213] <= 13'b0011010111010;
		Log_C0[214] <= 13'b0011010110101;
		Log_C0[215] <= 13'b0011010110000;
		Log_C0[216] <= 13'b0011010101100;
		Log_C0[217] <= 13'b0011010100111;
		Log_C0[218] <= 13'b0011010100010;
		Log_C0[219] <= 13'b0011010011110;
		Log_C0[220] <= 13'b0011010011001;
		Log_C0[221] <= 13'b0011010010100;
		Log_C0[222] <= 13'b0011010010000;
		Log_C0[223] <= 13'b0011010001011;
		Log_C0[224] <= 13'b0011010000110;
		Log_C0[225] <= 13'b0011010000010;
		Log_C0[226] <= 13'b0011001111101;
		Log_C0[227] <= 13'b0011001111001;
		Log_C0[228] <= 13'b0011001110100;
		Log_C0[229] <= 13'b0011001110000;
		Log_C0[230] <= 13'b0011001101011;
		Log_C0[231] <= 13'b0011001100111;
		Log_C0[232] <= 13'b0011001100011;
		Log_C0[233] <= 13'b0011001011110;
		Log_C0[234] <= 13'b0011001011010;
		Log_C0[235] <= 13'b0011001010101;
		Log_C0[236] <= 13'b0011001010001;
		Log_C0[237] <= 13'b0011001001101;
		Log_C0[238] <= 13'b0011001001001;
		Log_C0[239] <= 13'b0011001000100;
		Log_C0[240] <= 13'b0011001000000;
		Log_C0[241] <= 13'b0011000111100;
		Log_C0[242] <= 13'b0011000110111;
		Log_C0[243] <= 13'b0011000110011;
		Log_C0[244] <= 13'b0011000101111;
		Log_C0[245] <= 13'b0011000101011;
		Log_C0[246] <= 13'b0011000100111;
		Log_C0[247] <= 13'b0011000100011;
		Log_C0[248] <= 13'b0011000011110;
		Log_C0[249] <= 13'b0011000011010;
		Log_C0[250] <= 13'b0011000010110;
		Log_C0[251] <= 13'b0011000010010;
		Log_C0[252] <= 13'b0011000001110;
		Log_C0[253] <= 13'b0011000001010;
		Log_C0[254] <= 13'b0011000000110;
		Log_C0[255] <= 13'b0011000000010;

	end
end
endmodule

/* Verilog code for The Logarithm block of AWGN Project

	Log takes input of 31 bits in Q23 format.
	Output is 17 bits wide in Q13 format.

	Method: Polyfit coffecients are found using MATLAB. A memory is created to store those coefficients.

	Latency = 3;

*/


module SQRT_POLY(input clk, input reset, input [30:0] RootIn, output reg [16:0] RootOut);

bit [11:0] Sqrt_C1[64];
bit [19:0] Sqrt_C0[64];

reg [42:0] Term1;
reg [19:0] Term2;

reg [42:0] Term11;
reg [19:0] Term21;
reg [12:0] Root;

reg [13:0] FractionBit;
reg [3:0] IntegerBits;

always @(posedge clk)
begin
	if(!reset)
	begin

		// Cycle 1
		Term1 <= RootIn * Sqrt_C1[RootIn[30:25]];
		Term2 <= Sqrt_C0[RootIn[30:25]];


		// Cycle 2
		FractionBit <= Term1[35:23] + Term2[16:4];
		//Pipelining
		Term11 <= Term1;
		Term21 <= Term2;

		// Cycle 3
		IntegerBits <=  Term11[39:36] + Term21[19:17] + FractionBit[13];
		Root[12:0] <=  FractionBit[12:0];	// Pipelining

		RootOut[12:0] <= Root[12:0];		
		RootOut[16:13] <= IntegerBits[3:0];

	end

	else begin

	// C1 Coefficient Table

		Sqrt_C1[0] <= 12'b100100010001;
		Sqrt_C1[1] <= 12'b010010101001;
		Sqrt_C1[2] <= 12'b001110010111;
		Sqrt_C1[3] <= 12'b001100000111;
		Sqrt_C1[4] <= 12'b001010101011;
		Sqrt_C1[5] <= 12'b001001101010;
		Sqrt_C1[6] <= 12'b001000111000;
		Sqrt_C1[7] <= 12'b001000010001;
		Sqrt_C1[8] <= 12'b000111110001;
		Sqrt_C1[9] <= 12'b000111010110;
		Sqrt_C1[10] <= 12'b000110111111;
		Sqrt_C1[11] <= 12'b000110101011;
		Sqrt_C1[12] <= 12'b000110011010;
		Sqrt_C1[13] <= 12'b000110001010;
		Sqrt_C1[14] <= 12'b000101111100;
		Sqrt_C1[15] <= 12'b000101110000;
		Sqrt_C1[16] <= 12'b000101100101;
		Sqrt_C1[17] <= 12'b000101011010;
		Sqrt_C1[18] <= 12'b000101010001;
		Sqrt_C1[19] <= 12'b000101001000;
		Sqrt_C1[20] <= 12'b000101000000;
		Sqrt_C1[21] <= 12'b000100111000;
		Sqrt_C1[22] <= 12'b000100110001;
		Sqrt_C1[23] <= 12'b000100101011;
		Sqrt_C1[24] <= 12'b000100100101;
		Sqrt_C1[25] <= 12'b000100011111;
		Sqrt_C1[26] <= 12'b000100011001;
		Sqrt_C1[27] <= 12'b000100010100;
		Sqrt_C1[28] <= 12'b000100001111;
		Sqrt_C1[29] <= 12'b000100001011;
		Sqrt_C1[30] <= 12'b000100000110;
		Sqrt_C1[31] <= 12'b000100000010;
		Sqrt_C1[32] <= 12'b000011111110;
		Sqrt_C1[33] <= 12'b000011111010;
		Sqrt_C1[34] <= 12'b000011110111;
		Sqrt_C1[35] <= 12'b000011110011;
		Sqrt_C1[36] <= 12'b000011110000;
		Sqrt_C1[37] <= 12'b000011101100;
		Sqrt_C1[38] <= 12'b000011101001;
		Sqrt_C1[39] <= 12'b000011100110;
		Sqrt_C1[40] <= 12'b000011100100;
		Sqrt_C1[41] <= 12'b000011100001;
		Sqrt_C1[42] <= 12'b000011011110;
		Sqrt_C1[43] <= 12'b000011011100;
		Sqrt_C1[44] <= 12'b000011011001;
		Sqrt_C1[45] <= 12'b000011010111;
		Sqrt_C1[46] <= 12'b000011010100;
		Sqrt_C1[47] <= 12'b000011010010;
		Sqrt_C1[48] <= 12'b000011010000;
		Sqrt_C1[49] <= 12'b000011001110;
		Sqrt_C1[50] <= 12'b000011001100;
		Sqrt_C1[51] <= 12'b000011001010;
		Sqrt_C1[52] <= 12'b000011001000;
		Sqrt_C1[53] <= 12'b000011000110;
		Sqrt_C1[54] <= 12'b000011000100;
		Sqrt_C1[55] <= 12'b000011000010;
		Sqrt_C1[56] <= 12'b000011000001;
		Sqrt_C1[57] <= 12'b000010111111;
		Sqrt_C1[58] <= 12'b000010111101;
		Sqrt_C1[59] <= 12'b000010111100;
		Sqrt_C1[60] <= 12'b000010111010;
		Sqrt_C1[61] <= 12'b000010111001;
		Sqrt_C1[62] <= 12'b000010110111;
		Sqrt_C1[63] <= 12'b000010110110;

	// C0 Coefficient Table

		Sqrt_C0[0] <= 20'b00001100000001100001;
		Sqrt_C0[1] <= 20'b00011011001101011001;
		Sqrt_C0[2] <= 20'b00100011100011000010;
		Sqrt_C0[3] <= 20'b00101010001100011011;
		Sqrt_C0[4] <= 20'b00101111111001111101;
		Sqrt_C0[5] <= 20'b00110100111111110000;
		Sqrt_C0[6] <= 20'b00111001101000100111;
		Sqrt_C0[7] <= 20'b00111101111011001000;
		Sqrt_C0[8] <= 20'b01000001111011101111;
		Sqrt_C0[9] <= 20'b01000101101101100011;
		Sqrt_C0[10] <= 20'b01001001010010110111;
		Sqrt_C0[11] <= 20'b01001100101101011101;
		Sqrt_C0[12] <= 20'b01001111111110101101;
		Sqrt_C0[13] <= 20'b01010011000111101101;
		Sqrt_C0[14] <= 20'b01010110001001010111;
		Sqrt_C0[15] <= 20'b01011001000100011101;
		Sqrt_C0[16] <= 20'b01011011111001100101;
		Sqrt_C0[17] <= 20'b01011110101001010010;
		Sqrt_C0[18] <= 20'b01100001010100000010;
		Sqrt_C0[19] <= 20'b01100011111010001101;
		Sqrt_C0[20] <= 20'b01100110011100001011;
		Sqrt_C0[21] <= 20'b01101000111010001111;
		Sqrt_C0[22] <= 20'b01101011010100101010;
		Sqrt_C0[23] <= 20'b01101101101011101100;
		Sqrt_C0[24] <= 20'b01101111111111100010;
		Sqrt_C0[25] <= 20'b01110010010000011000;
		Sqrt_C0[26] <= 20'b01110100011110011010;
		Sqrt_C0[27] <= 20'b01110110101001110010;
		Sqrt_C0[28] <= 20'b01111000110010101010;
		Sqrt_C0[29] <= 20'b01111010111001001001;
		Sqrt_C0[30] <= 20'b01111100111101010111;
		Sqrt_C0[31] <= 20'b01111110111111011011;
		Sqrt_C0[32] <= 20'b10000000111111011100;
		Sqrt_C0[33] <= 20'b10000010111101100000;
		Sqrt_C0[34] <= 20'b10000100111001101101;
		Sqrt_C0[35] <= 20'b10000110110100000111;
		Sqrt_C0[36] <= 20'b10001000101100110011;
		Sqrt_C0[37] <= 20'b10001010100011110110;
		Sqrt_C0[38] <= 20'b10001100011001010101;
		Sqrt_C0[39] <= 20'b10001110001101010010;
		Sqrt_C0[40] <= 20'b10001111111111110010;
		Sqrt_C0[41] <= 20'b10010001110000111000;
		Sqrt_C0[42] <= 20'b10010011100000100111;
		Sqrt_C0[43] <= 20'b10010101001111000010;
		Sqrt_C0[44] <= 20'b10010110111100001101;
		Sqrt_C0[45] <= 20'b10011000101000001010;
		Sqrt_C0[46] <= 20'b10011010010010111011;
		Sqrt_C0[47] <= 20'b10011011111100100011;
		Sqrt_C0[48] <= 20'b10011101100101000100;
		Sqrt_C0[49] <= 20'b10011111001100100000;
		Sqrt_C0[50] <= 20'b10100000110010111010;
		Sqrt_C0[51] <= 20'b10100010011000010100;
		Sqrt_C0[52] <= 20'b10100011111100101110;
		Sqrt_C0[53] <= 20'b10100101100000001100;
		Sqrt_C0[54] <= 20'b10100111000010101111;
		Sqrt_C0[55] <= 20'b10101000100100011000;
		Sqrt_C0[56] <= 20'b10101010000101001001;
		Sqrt_C0[57] <= 20'b10101011100101000011;
		Sqrt_C0[58] <= 20'b10101101000100001000;
		Sqrt_C0[59] <= 20'b10101110100010011001;
		Sqrt_C0[60] <= 20'b10101111111111111000;
		Sqrt_C0[61] <= 20'b10110001011100100110;
		Sqrt_C0[62] <= 20'b10110010111000100011;
		Sqrt_C0[63] <= 20'b10110100010011110010;

	end
end
endmodule

/* Module to calculate sin of the input signal (16,16) bits 

Func - 	0 for sine
	1 for Cosine

Latency = 2 clock cycle

*/

module SinBlock(input clk, input reset, input func, input [15:0] x, output reg [15:0] sinValue);

reg [11:0] Sin_C1[128];
reg [18:0] Sin_C0[128];

reg [25:0] Term1;
reg [32:0] Term2;
reg sValue, s1;
reg [6:0] Address;

always @(posedge clk)
begin
	if(!reset)
	begin

		// Cycle 1 get address
	
		
		// Cycle 2
		Term1 <= Sin_C1[Address] * x[13:0];
		Term2 <= Sin_C0[Address];
		s1 <= sValue;

		// Cycle 3
		sinValue [14:0] <= Term1[25:11] + Term2[32:18];
		sinValue [15] <= s1;

		case( {func, x[15:14]} )
		// Sine Calculation
	
		3'b000 : begin
				sValue <= 1'b0;
				Address <= (7'b1111_111 - x[14:8]);
			end

		3'b001 : begin
				sValue <= 1'b0;
				Address <= x[14:8];
			end
	
		3'b010 : begin
				sValue <= 1'b1;
				Address <= (7'b1111_111 - x[14:8]);
			end
	
		3'b011 : begin
				sValue <= 1'b1;
				Address <= x[14:8];
			end

		// Cosine Calculation

		3'b100 : begin
				sValue <= 1'b0;
				Address <= x[14:8];
			end

		3'b101 : begin
				sValue <= 1'b1;
				Address <= (7'b1111_111 - x[14:8]);
			end

		3'b110 : begin
				sValue <= 1'b1;
				Address <= x[14:8];
			end
	
		3'b111 : begin
				sValue <= 1'b0;
				Address <= (7'b1111_111 - x[14:8]);
			end	

		endcase


	end // reset

	else
	begin

		Sin_C0[0] <= 19'b1000000000000000011;
		Sin_C0[1] <= 19'b1000000000000101011;
		Sin_C0[2] <= 19'b1000000000001111010;
		Sin_C0[3] <= 19'b1000000000011110000;
		Sin_C0[4] <= 19'b1000000000110001110;
		Sin_C0[5] <= 19'b1000000001001010011;
		Sin_C0[6] <= 19'b1000000001100111111;
		Sin_C0[7] <= 19'b1000000010001010010;
		Sin_C0[8] <= 19'b1000000010110001101;
		Sin_C0[9] <= 19'b1000000011011101110;
		Sin_C0[10] <= 19'b1000000100001110110;
		Sin_C0[11] <= 19'b1000000101000100100;
		Sin_C0[12] <= 19'b1000000101111111000;
		Sin_C0[13] <= 19'b1000000110111110011;
		Sin_C0[14] <= 19'b1000001000000010100;
		Sin_C0[15] <= 19'b1000001001001011010;
		Sin_C0[16] <= 19'b1000001010011000101;
		Sin_C0[17] <= 19'b1000001011101010110;
		Sin_C0[18] <= 19'b1000001101000001011;
		Sin_C0[19] <= 19'b1000001110011100101;
		Sin_C0[20] <= 19'b1000001111111100011;
		Sin_C0[21] <= 19'b1000010001100000101;
		Sin_C0[22] <= 19'b1000010011001001010;
		Sin_C0[23] <= 19'b1000010100110110010;
		Sin_C0[24] <= 19'b1000010110100111100;
		Sin_C0[25] <= 19'b1000011000011101001;
		Sin_C0[26] <= 19'b1000011010010111000;
		Sin_C0[27] <= 19'b1000011100010101000;
		Sin_C0[28] <= 19'b1000011110010111000;
		Sin_C0[29] <= 19'b1000100000011101010;
		Sin_C0[30] <= 19'b1000100010100111011;
		Sin_C0[31] <= 19'b1000100100110101011;
		Sin_C0[32] <= 19'b1000100111000111010;
		Sin_C0[33] <= 19'b1000101001011100111;
		Sin_C0[34] <= 19'b1000101011110110010;
		Sin_C0[35] <= 19'b1000101110010011011;
		Sin_C0[36] <= 19'b1000110000110011111;
		Sin_C0[37] <= 19'b1000110011011000000;
		Sin_C0[38] <= 19'b1000110101111111100;
		Sin_C0[39] <= 19'b1000111000101010011;
		Sin_C0[40] <= 19'b1000111011011000011;
		Sin_C0[41] <= 19'b1000111110001001101;
		Sin_C0[42] <= 19'b1001000000111110000;
		Sin_C0[43] <= 19'b1001000011110101011;
		Sin_C0[44] <= 19'b1001000110101111100;
		Sin_C0[45] <= 19'b1001001001101100101;
		Sin_C0[46] <= 19'b1001001100101100011;
		Sin_C0[47] <= 19'b1001001111101110110;
		Sin_C0[48] <= 19'b1001010010110011110;
		Sin_C0[49] <= 19'b1001010101111011001;
		Sin_C0[50] <= 19'b1001011001000100111;
		Sin_C0[51] <= 19'b1001011100010000111;
		Sin_C0[52] <= 19'b1001011111011110111;
		Sin_C0[53] <= 19'b1001100010101111001;
		Sin_C0[54] <= 19'b1001100110000001001;
		Sin_C0[55] <= 19'b1001101001010101000;
		Sin_C0[56] <= 19'b1001101100101010101;
		Sin_C0[57] <= 19'b1001110000000001111;
		Sin_C0[58] <= 19'b1001110011011010101;
		Sin_C0[59] <= 19'b1001110110110100110;
		Sin_C0[60] <= 19'b1001111010010000001;
		Sin_C0[61] <= 19'b1001111101101100101;
		Sin_C0[62] <= 19'b1010000001001010010;
		Sin_C0[63] <= 19'b1010000100101000110;
		Sin_C0[64] <= 19'b1010001000001000000;
		Sin_C0[65] <= 19'b1010001011101000001;
		Sin_C0[66] <= 19'b1010001111001000101;
		Sin_C0[67] <= 19'b1010010010101001101;
		Sin_C0[68] <= 19'b1010010110001011000;
		Sin_C0[69] <= 19'b1010011001101100100;
		Sin_C0[70] <= 19'b1010011101001110001;
		Sin_C0[71] <= 19'b1010100000101111110;
		Sin_C0[72] <= 19'b1010100100010001001;
		Sin_C0[73] <= 19'b1010100111110010010;
		Sin_C0[74] <= 19'b1010101011010010111;
		Sin_C0[75] <= 19'b1010101110110011000;
		Sin_C0[76] <= 19'b1010110010010010011;
		Sin_C0[77] <= 19'b1010110101110001000;
		Sin_C0[78] <= 19'b1010111001001110101;
		Sin_C0[79] <= 19'b1010111100101011001;
		Sin_C0[80] <= 19'b1011000000000110100;
		Sin_C0[81] <= 19'b1011000011100000100;
		Sin_C0[82] <= 19'b1011000110111001000;
		Sin_C0[83] <= 19'b1011001010001111111;
		Sin_C0[84] <= 19'b1011001101100100111;
		Sin_C0[85] <= 19'b1011010000111000001;
		Sin_C0[86] <= 19'b1011010100001001010;
		Sin_C0[87] <= 19'b1011010111011000011;
		Sin_C0[88] <= 19'b1011011010100101000;
		Sin_C0[89] <= 19'b1011011101101111010;
		Sin_C0[90] <= 19'b1011100000110111000;
		Sin_C0[91] <= 19'b1011100011111011111;
		Sin_C0[92] <= 19'b1011100110111110000;
		Sin_C0[93] <= 19'b1011101001111101001;
		Sin_C0[94] <= 19'b1011101100111001001;
		Sin_C0[95] <= 19'b1011101111110001111;
		Sin_C0[96] <= 19'b1011110010100111001;
		Sin_C0[97] <= 19'b1011110101011000111;
		Sin_C0[98] <= 19'b1011111000000110111;
		Sin_C0[99] <= 19'b1011111010110001001;
		Sin_C0[100] <= 19'b1011111101010111011;
		Sin_C0[101] <= 19'b1011111111111001100;
		Sin_C0[102] <= 19'b1100000010010111011;
		Sin_C0[103] <= 19'b1100000100110000111;
		Sin_C0[104] <= 19'b1100000111000101111;
		Sin_C0[105] <= 19'b1100001001010110001;
		Sin_C0[106] <= 19'b1100001011100001101;
		Sin_C0[107] <= 19'b1100001101101000010;
		Sin_C0[108] <= 19'b1100001111101001110;
		Sin_C0[109] <= 19'b1100010001100110000;
		Sin_C0[110] <= 19'b1100010011011100111;
		Sin_C0[111] <= 19'b1100010101001110011;
		Sin_C0[112] <= 19'b1100010110111010010;
		Sin_C0[113] <= 19'b1100011000100000010;
		Sin_C0[114] <= 19'b1100011010000000011;
		Sin_C0[115] <= 19'b1100011011011010101;
		Sin_C0[116] <= 19'b1100011100101110100;
		Sin_C0[117] <= 19'b1100011101111100010;
		Sin_C0[118] <= 19'b1100011111000011100;
		Sin_C0[119] <= 19'b1100100000000100010;
		Sin_C0[120] <= 19'b1100100000111110010;
		Sin_C0[121] <= 19'b1100100001110001100;
		Sin_C0[122] <= 19'b1100100010011101110;
		Sin_C0[123] <= 19'b1100100011000011000;
		Sin_C0[124] <= 19'b1100100011100001000;
		Sin_C0[125] <= 19'b1100100011110111110;
		Sin_C0[126] <= 19'b1100100100000111000;
		Sin_C0[127] <= 19'b1100100100001110101;

		Sin_C1[0] <= 12'b000000001101;
		Sin_C1[1] <= 12'b000000100110;
		Sin_C1[2] <= 12'b000000111111;
		Sin_C1[3] <= 12'b000001011000;
		Sin_C1[4] <= 12'b000001110001;
		Sin_C1[5] <= 12'b000010001010;
		Sin_C1[6] <= 12'b000010100011;
		Sin_C1[7] <= 12'b000010111100;
		Sin_C1[8] <= 12'b000011010101;
		Sin_C1[9] <= 12'b000011101110;
		Sin_C1[10] <= 12'b000100000111;
		Sin_C1[11] <= 12'b000100100000;
		Sin_C1[12] <= 12'b000100111001;
		Sin_C1[13] <= 12'b000101010010;
		Sin_C1[14] <= 12'b000101101011;
		Sin_C1[15] <= 12'b000110000011;
		Sin_C1[16] <= 12'b000110011100;
		Sin_C1[17] <= 12'b000110110100;
		Sin_C1[18] <= 12'b000111001101;
		Sin_C1[19] <= 12'b000111100101;
		Sin_C1[20] <= 12'b000111111110;
		Sin_C1[21] <= 12'b001000010110;
		Sin_C1[22] <= 12'b001000101110;
		Sin_C1[23] <= 12'b001001000110;
		Sin_C1[24] <= 12'b001001011111;
		Sin_C1[25] <= 12'b001001110110;
		Sin_C1[26] <= 12'b001010001110;
		Sin_C1[27] <= 12'b001010100110;
		Sin_C1[28] <= 12'b001010111110;
		Sin_C1[29] <= 12'b001011010101;
		Sin_C1[30] <= 12'b001011101101;
		Sin_C1[31] <= 12'b001100000100;
		Sin_C1[32] <= 12'b001100011011;
		Sin_C1[33] <= 12'b001100110010;
		Sin_C1[34] <= 12'b001101001001;
		Sin_C1[35] <= 12'b001101100000;
		Sin_C1[36] <= 12'b001101110111;
		Sin_C1[37] <= 12'b001110001110;
		Sin_C1[38] <= 12'b001110100100;
		Sin_C1[39] <= 12'b001110111010;
		Sin_C1[40] <= 12'b001111010000;
		Sin_C1[41] <= 12'b001111100110;
		Sin_C1[42] <= 12'b001111111100;
		Sin_C1[43] <= 12'b010000010010;
		Sin_C1[44] <= 12'b010000101000;
		Sin_C1[45] <= 12'b010000111101;
		Sin_C1[46] <= 12'b010001010010;
		Sin_C1[47] <= 12'b010001100111;
		Sin_C1[48] <= 12'b010001111100;
		Sin_C1[49] <= 12'b010010010001;
		Sin_C1[50] <= 12'b010010100110;
		Sin_C1[51] <= 12'b010010111010;
		Sin_C1[52] <= 12'b010011001110;
		Sin_C1[53] <= 12'b010011100010;
		Sin_C1[54] <= 12'b010011110110;
		Sin_C1[55] <= 12'b010100001001;
		Sin_C1[56] <= 12'b010100011101;
		Sin_C1[57] <= 12'b010100110000;
		Sin_C1[58] <= 12'b010101000011;
		Sin_C1[59] <= 12'b010101010110;
		Sin_C1[60] <= 12'b010101101001;
		Sin_C1[61] <= 12'b010101111011;
		Sin_C1[62] <= 12'b010110001101;
		Sin_C1[63] <= 12'b010110011111;
		Sin_C1[64] <= 12'b010110110001;
		Sin_C1[65] <= 12'b010111000011;
		Sin_C1[66] <= 12'b010111010100;
		Sin_C1[67] <= 12'b010111100101;
		Sin_C1[68] <= 12'b010111110110;
		Sin_C1[69] <= 12'b011000000111;
		Sin_C1[70] <= 12'b011000010111;
		Sin_C1[71] <= 12'b011000100111;
		Sin_C1[72] <= 12'b011000110111;
		Sin_C1[73] <= 12'b011001000111;
		Sin_C1[74] <= 12'b011001010110;
		Sin_C1[75] <= 12'b011001100101;
		Sin_C1[76] <= 12'b011001110100;
		Sin_C1[77] <= 12'b011010000011;
		Sin_C1[78] <= 12'b011010010010;
		Sin_C1[79] <= 12'b011010100000;
		Sin_C1[80] <= 12'b011010101110;
		Sin_C1[81] <= 12'b011010111011;
		Sin_C1[82] <= 12'b011011001001;
		Sin_C1[83] <= 12'b011011010110;
		Sin_C1[84] <= 12'b011011100011;
		Sin_C1[85] <= 12'b011011110000;
		Sin_C1[86] <= 12'b011011111100;
		Sin_C1[87] <= 12'b011100001000;
		Sin_C1[88] <= 12'b011100010100;
		Sin_C1[89] <= 12'b011100100000;
		Sin_C1[90] <= 12'b011100101011;
		Sin_C1[91] <= 12'b011100110110;
		Sin_C1[92] <= 12'b011101000001;
		Sin_C1[93] <= 12'b011101001011;
		Sin_C1[94] <= 12'b011101010101;
		Sin_C1[95] <= 12'b011101011111;
		Sin_C1[96] <= 12'b011101101001;
		Sin_C1[97] <= 12'b011101110010;
		Sin_C1[98] <= 12'b011101111011;
		Sin_C1[99] <= 12'b011110000100;
		Sin_C1[100] <= 12'b011110001100;
		Sin_C1[101] <= 12'b011110010101;
		Sin_C1[102] <= 12'b011110011101;
		Sin_C1[103] <= 12'b011110100100;
		Sin_C1[104] <= 12'b011110101011;
		Sin_C1[105] <= 12'b011110110010;
		Sin_C1[106] <= 12'b011110111001;
		Sin_C1[107] <= 12'b011111000000;
		Sin_C1[108] <= 12'b011111000110;
		Sin_C1[109] <= 12'b011111001011;
		Sin_C1[110] <= 12'b011111010001;
		Sin_C1[111] <= 12'b011111010110;
		Sin_C1[112] <= 12'b011111011011;
		Sin_C1[113] <= 12'b011111100000;
		Sin_C1[114] <= 12'b011111100100;
		Sin_C1[115] <= 12'b011111101000;
		Sin_C1[116] <= 12'b011111101100;
		Sin_C1[117] <= 12'b011111101111;
		Sin_C1[118] <= 12'b011111110010;
		Sin_C1[119] <= 12'b011111110101;
		Sin_C1[120] <= 12'b011111110111;
		Sin_C1[121] <= 12'b011111111001;
		Sin_C1[122] <= 12'b011111111011;
		Sin_C1[123] <= 12'b011111111101;
		Sin_C1[124] <= 12'b011111111110;
		Sin_C1[125] <= 12'b011111111111;
		Sin_C1[126] <= 12'b100000000000;
		Sin_C1[127] <= 12'b100000000000;
	end
end

endmodule

