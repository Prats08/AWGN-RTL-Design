
module SinBlock_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   \A[9] , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59;
  assign SUM[10] = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];

  AO6 U2 ( .A(n16), .B(n3), .C(n17), .Z(n15) );
  OR2P U3 ( .A(B[11]), .B(A[11]), .Z(n1) );
  AN2P U4 ( .A(n1), .B(n59), .Z(SUM[11]) );
  AO6 U5 ( .A(n13), .B(n14), .C(n56), .Z(n53) );
  AO7 U6 ( .A(n52), .B(n53), .C(n54), .Z(n48) );
  AO6 U7 ( .A(n11), .B(n48), .C(n49), .Z(n45) );
  IVP U8 ( .A(n50), .Z(n11) );
  AO7 U9 ( .A(n44), .B(n45), .C(n46), .Z(n40) );
  AO6 U10 ( .A(n9), .B(n40), .C(n41), .Z(n37) );
  IVP U11 ( .A(n42), .Z(n9) );
  AO7 U12 ( .A(n36), .B(n37), .C(n38), .Z(n32) );
  AO6 U13 ( .A(n7), .B(n32), .C(n33), .Z(n29) );
  IVP U14 ( .A(n34), .Z(n7) );
  AO6 U15 ( .A(n5), .B(n24), .C(n25), .Z(n21) );
  IVP U16 ( .A(n26), .Z(n5) );
  IVP U17 ( .A(n59), .Z(n14) );
  IVP U18 ( .A(n22), .Z(n4) );
  IVP U19 ( .A(n30), .Z(n6) );
  IVP U20 ( .A(n38), .Z(n8) );
  IVP U21 ( .A(n46), .Z(n10) );
  IVP U22 ( .A(n54), .Z(n12) );
  IVP U23 ( .A(n18), .Z(n3) );
  NR2 U24 ( .A(B[12]), .B(A[12]), .Z(n57) );
  EN U25 ( .A(B[23]), .B(n15), .Z(SUM[23]) );
  IVP U26 ( .A(n57), .Z(n13) );
  EO U27 ( .A(n16), .B(n19), .Z(SUM[22]) );
  NR2 U28 ( .A(n17), .B(n18), .Z(n19) );
  NR2 U29 ( .A(B[22]), .B(A[22]), .Z(n18) );
  AN2 U30 ( .A(B[22]), .B(A[22]), .Z(n17) );
  AO7 U31 ( .A(n20), .B(n21), .C(n22), .Z(n16) );
  EN U32 ( .A(n21), .B(n23), .Z(SUM[21]) );
  NR2 U33 ( .A(n4), .B(n20), .Z(n23) );
  NR2 U34 ( .A(B[21]), .B(A[21]), .Z(n20) );
  ND2 U35 ( .A(B[21]), .B(A[21]), .Z(n22) );
  EO U36 ( .A(n24), .B(n27), .Z(SUM[20]) );
  NR2 U37 ( .A(n25), .B(n26), .Z(n27) );
  NR2 U38 ( .A(B[20]), .B(A[20]), .Z(n26) );
  AN2 U39 ( .A(B[20]), .B(A[20]), .Z(n25) );
  AO7 U40 ( .A(n28), .B(n29), .C(n30), .Z(n24) );
  EN U41 ( .A(n29), .B(n31), .Z(SUM[19]) );
  NR2 U42 ( .A(n6), .B(n28), .Z(n31) );
  NR2 U43 ( .A(B[19]), .B(A[19]), .Z(n28) );
  ND2 U44 ( .A(B[19]), .B(A[19]), .Z(n30) );
  EO U45 ( .A(n32), .B(n35), .Z(SUM[18]) );
  NR2 U46 ( .A(n33), .B(n34), .Z(n35) );
  NR2 U47 ( .A(B[18]), .B(A[18]), .Z(n34) );
  AN2 U48 ( .A(B[18]), .B(A[18]), .Z(n33) );
  EN U49 ( .A(n37), .B(n39), .Z(SUM[17]) );
  NR2 U50 ( .A(n8), .B(n36), .Z(n39) );
  NR2 U51 ( .A(B[17]), .B(A[17]), .Z(n36) );
  ND2 U52 ( .A(B[17]), .B(A[17]), .Z(n38) );
  EO U53 ( .A(n40), .B(n43), .Z(SUM[16]) );
  NR2 U54 ( .A(n41), .B(n42), .Z(n43) );
  NR2 U55 ( .A(B[16]), .B(A[16]), .Z(n42) );
  AN2 U56 ( .A(B[16]), .B(A[16]), .Z(n41) );
  EN U57 ( .A(n45), .B(n47), .Z(SUM[15]) );
  NR2 U58 ( .A(n10), .B(n44), .Z(n47) );
  NR2 U59 ( .A(B[15]), .B(A[15]), .Z(n44) );
  ND2 U60 ( .A(B[15]), .B(A[15]), .Z(n46) );
  EO U61 ( .A(n48), .B(n51), .Z(SUM[14]) );
  NR2 U62 ( .A(n49), .B(n50), .Z(n51) );
  NR2 U63 ( .A(B[14]), .B(A[14]), .Z(n50) );
  AN2 U64 ( .A(B[14]), .B(A[14]), .Z(n49) );
  EN U65 ( .A(n53), .B(n55), .Z(SUM[13]) );
  NR2 U66 ( .A(n12), .B(n52), .Z(n55) );
  NR2 U67 ( .A(B[13]), .B(A[13]), .Z(n52) );
  ND2 U68 ( .A(B[13]), .B(A[13]), .Z(n54) );
  EO U69 ( .A(n14), .B(n58), .Z(SUM[12]) );
  NR2 U70 ( .A(n56), .B(n57), .Z(n58) );
  AN2 U71 ( .A(B[12]), .B(A[12]), .Z(n56) );
  ND2 U72 ( .A(B[11]), .B(A[11]), .Z(n59) );
endmodule


module SinBlock_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [11:0] A;
  input [13:0] B;
  output [25:0] PRODUCT;
  input TC;
  wire   \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][13] ,
         \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] ,
         \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] ,
         \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][13] , \ab[8][12] , \ab[8][11] ,
         \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] , \ab[8][6] ,
         \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] ,
         \ab[8][0] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][13] ,
         \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] ,
         \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] ,
         \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][13] , \ab[3][12] , \ab[3][11] ,
         \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[0][13] , \ab[0][12] ,
         \ab[0][11] , \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] ,
         \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] ,
         \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] ,
         \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] ,
         \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] ,
         \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] ,
         \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][12] , \CARRYB[1][11] ,
         \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] ,
         \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[11][0] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][12] ,
         \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] ,
         \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] ,
         \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][12] ,
         \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] ,
         \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] ,
         \A2[17] , \A2[16] , \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] ,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8;

  SinBlock_DW01_add_1 FS_1 ( .A({1'b0, \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , 
        \A1[11] , \A1[10] , \SUMB[11][0] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[23] , \A2[22] , 
        \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , 
        \A2[14] , \A2[13] , \A2[12] , \A2[11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[25:11], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8}) );
  FA1A S5_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\ab[10][13] ), .CO(
        \CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S3_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\ab[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S3_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\ab[8][13] ), .CO(
        \CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S3_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\ab[7][13] ), .CO(
        \CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S3_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\ab[6][13] ), .CO(
        \CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S3_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\ab[5][13] ), .CO(
        \CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S3_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\ab[4][13] ), .CO(
        \CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S3_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\ab[3][13] ), .CO(
        \CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S3_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\ab[2][13] ), .CO(
        \CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S3_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\ab[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S4_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(
        \CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S4_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), .CO(
        \CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S4_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(
        \CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S4_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(
        \CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S4_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(
        \CARRYB[11][0] ), .S(\SUMB[11][0] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S4_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(
        \CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S4_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(
        \CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S4_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(
        \CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(
        \CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S4_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(
        \CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  EO U2 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A1[12] ) );
  EO U3 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A1[11] ) );
  EO U4 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A1[13] ) );
  EO U5 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A1[14] ) );
  EO U6 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  EO U7 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A1[15] ) );
  EO U8 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A1[16] ) );
  EO U9 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A1[17] ) );
  EO U10 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A1[18] ) );
  EO U11 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A1[19] ) );
  EO U12 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A1[20] ) );
  EO U13 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A1[21] ) );
  EO U14 ( .A(\CARRYB[11][12] ), .B(\ab[11][13] ), .Z(\A1[22] ) );
  EO U15 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A1[10] ) );
  NR2 U16 ( .A(n11), .B(n27), .Z(\ab[1][1] ) );
  IVP U17 ( .A(A[0]), .Z(n10) );
  NR2 U18 ( .A(n25), .B(n10), .Z(\ab[0][3] ) );
  EO U19 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U20 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U21 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U22 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U23 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U24 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U25 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U26 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U27 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U28 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U29 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  IVP U30 ( .A(A[1]), .Z(n11) );
  IVP U31 ( .A(A[2]), .Z(n12) );
  IVP U32 ( .A(A[3]), .Z(n13) );
  IVP U33 ( .A(A[4]), .Z(n14) );
  IVP U34 ( .A(A[5]), .Z(n15) );
  IVP U35 ( .A(B[3]), .Z(n25) );
  IVP U36 ( .A(B[2]), .Z(n26) );
  IVP U37 ( .A(B[4]), .Z(n24) );
  IVP U38 ( .A(B[1]), .Z(n27) );
  IVP U39 ( .A(B[5]), .Z(n23) );
  IVP U40 ( .A(B[6]), .Z(n22) );
  IVP U41 ( .A(A[6]), .Z(n16) );
  IVP U42 ( .A(B[7]), .Z(n21) );
  IVP U43 ( .A(B[8]), .Z(n3) );
  IVP U44 ( .A(B[9]), .Z(n4) );
  IVP U45 ( .A(B[0]), .Z(n28) );
  IVP U46 ( .A(B[10]), .Z(n5) );
  IVP U47 ( .A(A[7]), .Z(n17) );
  IVP U48 ( .A(B[11]), .Z(n6) );
  IVP U49 ( .A(B[12]), .Z(n7) );
  IVP U50 ( .A(A[8]), .Z(n18) );
  IVP U51 ( .A(B[13]), .Z(n8) );
  IVP U52 ( .A(A[9]), .Z(n19) );
  IVP U53 ( .A(A[10]), .Z(n20) );
  IVP U54 ( .A(A[11]), .Z(n9) );
  AN2P U55 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A2[11] ) );
  AN2P U56 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A2[14] ) );
  AN2P U57 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A2[15] ) );
  AN2P U58 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A2[16] ) );
  AN2P U59 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A2[17] ) );
  AN2P U60 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A2[18] ) );
  AN2P U61 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A2[19] ) );
  AN2P U62 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A2[20] ) );
  AN2P U63 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A2[21] ) );
  AN2P U64 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A2[22] ) );
  AN2P U65 ( .A(\CARRYB[11][12] ), .B(\ab[11][13] ), .Z(\A2[23] ) );
  AN2P U66 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U67 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U68 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U69 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U70 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U71 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U72 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U73 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U74 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U75 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U76 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U77 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U78 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A2[13] ) );
  AN2P U79 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A2[12] ) );
  NR2 U81 ( .A(n19), .B(n4), .Z(\ab[9][9] ) );
  NR2 U82 ( .A(n19), .B(n3), .Z(\ab[9][8] ) );
  NR2 U83 ( .A(n19), .B(n21), .Z(\ab[9][7] ) );
  NR2 U84 ( .A(n19), .B(n22), .Z(\ab[9][6] ) );
  NR2 U85 ( .A(n19), .B(n23), .Z(\ab[9][5] ) );
  NR2 U86 ( .A(n19), .B(n24), .Z(\ab[9][4] ) );
  NR2 U87 ( .A(n19), .B(n25), .Z(\ab[9][3] ) );
  NR2 U88 ( .A(n19), .B(n26), .Z(\ab[9][2] ) );
  NR2 U89 ( .A(n19), .B(n27), .Z(\ab[9][1] ) );
  NR2 U90 ( .A(n19), .B(n8), .Z(\ab[9][13] ) );
  NR2 U91 ( .A(n19), .B(n7), .Z(\ab[9][12] ) );
  NR2 U92 ( .A(n19), .B(n6), .Z(\ab[9][11] ) );
  NR2 U93 ( .A(n19), .B(n5), .Z(\ab[9][10] ) );
  NR2 U94 ( .A(n19), .B(n28), .Z(\ab[9][0] ) );
  NR2 U95 ( .A(n4), .B(n18), .Z(\ab[8][9] ) );
  NR2 U96 ( .A(n3), .B(n18), .Z(\ab[8][8] ) );
  NR2 U97 ( .A(n21), .B(n18), .Z(\ab[8][7] ) );
  NR2 U98 ( .A(n22), .B(n18), .Z(\ab[8][6] ) );
  NR2 U99 ( .A(n23), .B(n18), .Z(\ab[8][5] ) );
  NR2 U100 ( .A(n24), .B(n18), .Z(\ab[8][4] ) );
  NR2 U101 ( .A(n25), .B(n18), .Z(\ab[8][3] ) );
  NR2 U102 ( .A(n26), .B(n18), .Z(\ab[8][2] ) );
  NR2 U103 ( .A(n27), .B(n18), .Z(\ab[8][1] ) );
  NR2 U104 ( .A(n8), .B(n18), .Z(\ab[8][13] ) );
  NR2 U105 ( .A(n7), .B(n18), .Z(\ab[8][12] ) );
  NR2 U106 ( .A(n6), .B(n18), .Z(\ab[8][11] ) );
  NR2 U107 ( .A(n5), .B(n18), .Z(\ab[8][10] ) );
  NR2 U108 ( .A(n28), .B(n18), .Z(\ab[8][0] ) );
  NR2 U109 ( .A(n4), .B(n17), .Z(\ab[7][9] ) );
  NR2 U110 ( .A(n3), .B(n17), .Z(\ab[7][8] ) );
  NR2 U111 ( .A(n21), .B(n17), .Z(\ab[7][7] ) );
  NR2 U112 ( .A(n22), .B(n17), .Z(\ab[7][6] ) );
  NR2 U113 ( .A(n23), .B(n17), .Z(\ab[7][5] ) );
  NR2 U114 ( .A(n24), .B(n17), .Z(\ab[7][4] ) );
  NR2 U115 ( .A(n25), .B(n17), .Z(\ab[7][3] ) );
  NR2 U116 ( .A(n26), .B(n17), .Z(\ab[7][2] ) );
  NR2 U117 ( .A(n27), .B(n17), .Z(\ab[7][1] ) );
  NR2 U118 ( .A(n8), .B(n17), .Z(\ab[7][13] ) );
  NR2 U119 ( .A(n7), .B(n17), .Z(\ab[7][12] ) );
  NR2 U120 ( .A(n6), .B(n17), .Z(\ab[7][11] ) );
  NR2 U121 ( .A(n5), .B(n17), .Z(\ab[7][10] ) );
  NR2 U122 ( .A(n28), .B(n17), .Z(\ab[7][0] ) );
  NR2 U123 ( .A(n4), .B(n16), .Z(\ab[6][9] ) );
  NR2 U124 ( .A(n3), .B(n16), .Z(\ab[6][8] ) );
  NR2 U125 ( .A(n21), .B(n16), .Z(\ab[6][7] ) );
  NR2 U126 ( .A(n22), .B(n16), .Z(\ab[6][6] ) );
  NR2 U127 ( .A(n23), .B(n16), .Z(\ab[6][5] ) );
  NR2 U128 ( .A(n24), .B(n16), .Z(\ab[6][4] ) );
  NR2 U129 ( .A(n25), .B(n16), .Z(\ab[6][3] ) );
  NR2 U130 ( .A(n26), .B(n16), .Z(\ab[6][2] ) );
  NR2 U131 ( .A(n27), .B(n16), .Z(\ab[6][1] ) );
  NR2 U132 ( .A(n8), .B(n16), .Z(\ab[6][13] ) );
  NR2 U133 ( .A(n7), .B(n16), .Z(\ab[6][12] ) );
  NR2 U134 ( .A(n6), .B(n16), .Z(\ab[6][11] ) );
  NR2 U135 ( .A(n5), .B(n16), .Z(\ab[6][10] ) );
  NR2 U136 ( .A(n28), .B(n16), .Z(\ab[6][0] ) );
  NR2 U137 ( .A(n4), .B(n15), .Z(\ab[5][9] ) );
  NR2 U138 ( .A(n3), .B(n15), .Z(\ab[5][8] ) );
  NR2 U139 ( .A(n21), .B(n15), .Z(\ab[5][7] ) );
  NR2 U140 ( .A(n22), .B(n15), .Z(\ab[5][6] ) );
  NR2 U141 ( .A(n23), .B(n15), .Z(\ab[5][5] ) );
  NR2 U142 ( .A(n24), .B(n15), .Z(\ab[5][4] ) );
  NR2 U143 ( .A(n25), .B(n15), .Z(\ab[5][3] ) );
  NR2 U144 ( .A(n26), .B(n15), .Z(\ab[5][2] ) );
  NR2 U145 ( .A(n27), .B(n15), .Z(\ab[5][1] ) );
  NR2 U146 ( .A(n8), .B(n15), .Z(\ab[5][13] ) );
  NR2 U147 ( .A(n7), .B(n15), .Z(\ab[5][12] ) );
  NR2 U148 ( .A(n6), .B(n15), .Z(\ab[5][11] ) );
  NR2 U149 ( .A(n5), .B(n15), .Z(\ab[5][10] ) );
  NR2 U150 ( .A(n28), .B(n15), .Z(\ab[5][0] ) );
  NR2 U151 ( .A(n4), .B(n14), .Z(\ab[4][9] ) );
  NR2 U152 ( .A(n3), .B(n14), .Z(\ab[4][8] ) );
  NR2 U153 ( .A(n21), .B(n14), .Z(\ab[4][7] ) );
  NR2 U154 ( .A(n22), .B(n14), .Z(\ab[4][6] ) );
  NR2 U155 ( .A(n23), .B(n14), .Z(\ab[4][5] ) );
  NR2 U156 ( .A(n24), .B(n14), .Z(\ab[4][4] ) );
  NR2 U157 ( .A(n25), .B(n14), .Z(\ab[4][3] ) );
  NR2 U158 ( .A(n26), .B(n14), .Z(\ab[4][2] ) );
  NR2 U159 ( .A(n27), .B(n14), .Z(\ab[4][1] ) );
  NR2 U160 ( .A(n8), .B(n14), .Z(\ab[4][13] ) );
  NR2 U161 ( .A(n7), .B(n14), .Z(\ab[4][12] ) );
  NR2 U162 ( .A(n6), .B(n14), .Z(\ab[4][11] ) );
  NR2 U163 ( .A(n5), .B(n14), .Z(\ab[4][10] ) );
  NR2 U164 ( .A(n28), .B(n14), .Z(\ab[4][0] ) );
  NR2 U165 ( .A(n4), .B(n13), .Z(\ab[3][9] ) );
  NR2 U166 ( .A(n3), .B(n13), .Z(\ab[3][8] ) );
  NR2 U167 ( .A(n21), .B(n13), .Z(\ab[3][7] ) );
  NR2 U168 ( .A(n22), .B(n13), .Z(\ab[3][6] ) );
  NR2 U169 ( .A(n23), .B(n13), .Z(\ab[3][5] ) );
  NR2 U170 ( .A(n24), .B(n13), .Z(\ab[3][4] ) );
  NR2 U171 ( .A(n25), .B(n13), .Z(\ab[3][3] ) );
  NR2 U172 ( .A(n26), .B(n13), .Z(\ab[3][2] ) );
  NR2 U173 ( .A(n27), .B(n13), .Z(\ab[3][1] ) );
  NR2 U174 ( .A(n8), .B(n13), .Z(\ab[3][13] ) );
  NR2 U175 ( .A(n7), .B(n13), .Z(\ab[3][12] ) );
  NR2 U176 ( .A(n6), .B(n13), .Z(\ab[3][11] ) );
  NR2 U177 ( .A(n5), .B(n13), .Z(\ab[3][10] ) );
  NR2 U178 ( .A(n28), .B(n13), .Z(\ab[3][0] ) );
  NR2 U179 ( .A(n4), .B(n12), .Z(\ab[2][9] ) );
  NR2 U180 ( .A(n3), .B(n12), .Z(\ab[2][8] ) );
  NR2 U181 ( .A(n21), .B(n12), .Z(\ab[2][7] ) );
  NR2 U182 ( .A(n22), .B(n12), .Z(\ab[2][6] ) );
  NR2 U183 ( .A(n23), .B(n12), .Z(\ab[2][5] ) );
  NR2 U184 ( .A(n24), .B(n12), .Z(\ab[2][4] ) );
  NR2 U185 ( .A(n25), .B(n12), .Z(\ab[2][3] ) );
  NR2 U186 ( .A(n26), .B(n12), .Z(\ab[2][2] ) );
  NR2 U187 ( .A(n27), .B(n12), .Z(\ab[2][1] ) );
  NR2 U188 ( .A(n8), .B(n12), .Z(\ab[2][13] ) );
  NR2 U189 ( .A(n7), .B(n12), .Z(\ab[2][12] ) );
  NR2 U190 ( .A(n6), .B(n12), .Z(\ab[2][11] ) );
  NR2 U191 ( .A(n5), .B(n12), .Z(\ab[2][10] ) );
  NR2 U192 ( .A(n28), .B(n12), .Z(\ab[2][0] ) );
  NR2 U193 ( .A(n4), .B(n11), .Z(\ab[1][9] ) );
  NR2 U194 ( .A(n3), .B(n11), .Z(\ab[1][8] ) );
  NR2 U195 ( .A(n21), .B(n11), .Z(\ab[1][7] ) );
  NR2 U196 ( .A(n22), .B(n11), .Z(\ab[1][6] ) );
  NR2 U197 ( .A(n23), .B(n11), .Z(\ab[1][5] ) );
  NR2 U198 ( .A(n24), .B(n11), .Z(\ab[1][4] ) );
  NR2 U199 ( .A(n25), .B(n11), .Z(\ab[1][3] ) );
  NR2 U200 ( .A(n26), .B(n11), .Z(\ab[1][2] ) );
  NR2 U201 ( .A(n8), .B(n11), .Z(\ab[1][13] ) );
  NR2 U202 ( .A(n7), .B(n11), .Z(\ab[1][12] ) );
  NR2 U203 ( .A(n6), .B(n11), .Z(\ab[1][11] ) );
  NR2 U204 ( .A(n5), .B(n11), .Z(\ab[1][10] ) );
  NR2 U205 ( .A(n4), .B(n9), .Z(\ab[11][9] ) );
  NR2 U206 ( .A(n3), .B(n9), .Z(\ab[11][8] ) );
  NR2 U207 ( .A(n21), .B(n9), .Z(\ab[11][7] ) );
  NR2 U208 ( .A(n22), .B(n9), .Z(\ab[11][6] ) );
  NR2 U209 ( .A(n23), .B(n9), .Z(\ab[11][5] ) );
  NR2 U210 ( .A(n24), .B(n9), .Z(\ab[11][4] ) );
  NR2 U211 ( .A(n25), .B(n9), .Z(\ab[11][3] ) );
  NR2 U212 ( .A(n26), .B(n9), .Z(\ab[11][2] ) );
  NR2 U213 ( .A(n27), .B(n9), .Z(\ab[11][1] ) );
  NR2 U214 ( .A(n8), .B(n9), .Z(\ab[11][13] ) );
  NR2 U215 ( .A(n7), .B(n9), .Z(\ab[11][12] ) );
  NR2 U216 ( .A(n6), .B(n9), .Z(\ab[11][11] ) );
  NR2 U217 ( .A(n5), .B(n9), .Z(\ab[11][10] ) );
  NR2 U218 ( .A(n28), .B(n9), .Z(\ab[11][0] ) );
  NR2 U219 ( .A(n4), .B(n20), .Z(\ab[10][9] ) );
  NR2 U220 ( .A(n3), .B(n20), .Z(\ab[10][8] ) );
  NR2 U221 ( .A(n21), .B(n20), .Z(\ab[10][7] ) );
  NR2 U222 ( .A(n22), .B(n20), .Z(\ab[10][6] ) );
  NR2 U223 ( .A(n23), .B(n20), .Z(\ab[10][5] ) );
  NR2 U224 ( .A(n24), .B(n20), .Z(\ab[10][4] ) );
  NR2 U225 ( .A(n25), .B(n20), .Z(\ab[10][3] ) );
  NR2 U226 ( .A(n26), .B(n20), .Z(\ab[10][2] ) );
  NR2 U227 ( .A(n27), .B(n20), .Z(\ab[10][1] ) );
  NR2 U228 ( .A(n8), .B(n20), .Z(\ab[10][13] ) );
  NR2 U229 ( .A(n7), .B(n20), .Z(\ab[10][12] ) );
  NR2 U230 ( .A(n6), .B(n20), .Z(\ab[10][11] ) );
  NR2 U231 ( .A(n5), .B(n20), .Z(\ab[10][10] ) );
  NR2 U232 ( .A(n28), .B(n20), .Z(\ab[10][0] ) );
  NR2 U233 ( .A(n4), .B(n10), .Z(\ab[0][9] ) );
  NR2 U234 ( .A(n3), .B(n10), .Z(\ab[0][8] ) );
  NR2 U235 ( .A(n21), .B(n10), .Z(\ab[0][7] ) );
  NR2 U236 ( .A(n22), .B(n10), .Z(\ab[0][6] ) );
  NR2 U237 ( .A(n23), .B(n10), .Z(\ab[0][5] ) );
  NR2 U238 ( .A(n24), .B(n10), .Z(\ab[0][4] ) );
  NR2 U239 ( .A(n26), .B(n10), .Z(\ab[0][2] ) );
  NR2 U240 ( .A(n8), .B(n10), .Z(\ab[0][13] ) );
  NR2 U241 ( .A(n7), .B(n10), .Z(\ab[0][12] ) );
  NR2 U242 ( .A(n6), .B(n10), .Z(\ab[0][11] ) );
  NR2 U243 ( .A(n5), .B(n10), .Z(\ab[0][10] ) );
  AN3 U244 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
endmodule


module SinBlock ( clk, reset, func, x, sinValue );
  input [15:0] x;
  output [15:0] sinValue;
  input clk, reset, func;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         \Term2[18] , N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, sValue, N57, n35, \add_29/carry[14] ,
         \add_29/carry[13] , \add_29/carry[12] , \add_29/carry[11] ,
         \add_29/carry[10] , \add_29/carry[9] , \add_29/carry[8] ,
         \add_29/carry[7] , \add_29/carry[6] , \add_29/carry[5] ,
         \add_29/carry[4] , \add_29/carry[3] , \add_29/carry[2] ,
         \add_29/carry[1] , n37, n38, n39, n40, n41, n42, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540;
  wire   [25:11] Term1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10;

  SinBlock_DW02_mult_0 mult_25 ( .A({n42, N9, N10, N11, N12, N13, N14, N15, 
        N16, N17, N18, N19}), .B(x[13:0]), .TC(1'b0), .PRODUCT({N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  FDS2L \Term1_reg[25]  ( .CR(1'b1), .D(N34), .LD(n540), .CP(clk), .Q(
        Term1[25]) );
  FDS2L \Term1_reg[24]  ( .CR(1'b1), .D(N33), .LD(n540), .CP(clk), .Q(
        Term1[24]) );
  FDS2L \Term1_reg[23]  ( .CR(1'b1), .D(N32), .LD(n540), .CP(clk), .Q(
        Term1[23]) );
  FDS2L \Term1_reg[22]  ( .CR(1'b1), .D(N31), .LD(n540), .CP(clk), .Q(
        Term1[22]) );
  FDS2L \Term1_reg[21]  ( .CR(1'b1), .D(N30), .LD(n540), .CP(clk), .Q(
        Term1[21]) );
  FDS2L \Term1_reg[20]  ( .CR(1'b1), .D(N29), .LD(n540), .CP(clk), .Q(
        Term1[20]) );
  FDS2L \Term1_reg[19]  ( .CR(1'b1), .D(N28), .LD(n540), .CP(clk), .Q(
        Term1[19]) );
  FDS2L \Term1_reg[18]  ( .CR(1'b1), .D(N27), .LD(n540), .CP(clk), .Q(
        Term1[18]) );
  FDS2L \Term1_reg[17]  ( .CR(1'b1), .D(N26), .LD(n540), .CP(clk), .Q(
        Term1[17]) );
  FDS2L \Term1_reg[16]  ( .CR(1'b1), .D(N25), .LD(n540), .CP(clk), .Q(
        Term1[16]) );
  FDS2L \Term1_reg[15]  ( .CR(1'b1), .D(N24), .LD(n540), .CP(clk), .Q(
        Term1[15]) );
  FDS2L \Term1_reg[14]  ( .CR(1'b1), .D(N23), .LD(n540), .CP(clk), .Q(
        Term1[14]) );
  FDS2L \Term1_reg[13]  ( .CR(1'b1), .D(N22), .LD(n540), .CP(clk), .Q(
        Term1[13]) );
  FDS2L \Term1_reg[12]  ( .CR(1'b1), .D(N21), .LD(n540), .CP(clk), .Q(
        Term1[12]) );
  FDS2L \Term1_reg[11]  ( .CR(1'b1), .D(N20), .LD(n540), .CP(clk), .Q(
        Term1[11]) );
  FDS2L \sinValue_reg[14]  ( .CR(1'b1), .D(N50), .LD(n540), .CP(clk), .Q(
        sinValue[14]) );
  FDS2L \sinValue_reg[13]  ( .CR(1'b1), .D(N49), .LD(n540), .CP(clk), .Q(
        sinValue[13]) );
  FDS2L \sinValue_reg[12]  ( .CR(1'b1), .D(N48), .LD(n540), .CP(clk), .Q(
        sinValue[12]) );
  FDS2L \sinValue_reg[11]  ( .CR(1'b1), .D(N47), .LD(n540), .CP(clk), .Q(
        sinValue[11]) );
  FDS2L \sinValue_reg[10]  ( .CR(1'b1), .D(N46), .LD(n540), .CP(clk), .Q(
        sinValue[10]) );
  FDS2L \sinValue_reg[9]  ( .CR(1'b1), .D(N45), .LD(n540), .CP(clk), .Q(
        sinValue[9]) );
  FDS2L \sinValue_reg[8]  ( .CR(1'b1), .D(N44), .LD(n540), .CP(clk), .Q(
        sinValue[8]) );
  FDS2L \sinValue_reg[7]  ( .CR(1'b1), .D(N43), .LD(n540), .CP(clk), .Q(
        sinValue[7]) );
  FDS2L \sinValue_reg[6]  ( .CR(1'b1), .D(N42), .LD(n540), .CP(clk), .Q(
        sinValue[6]) );
  FDS2L \sinValue_reg[5]  ( .CR(1'b1), .D(N41), .LD(n540), .CP(clk), .Q(
        sinValue[5]) );
  FDS2L \sinValue_reg[4]  ( .CR(1'b1), .D(N40), .LD(n540), .CP(clk), .Q(
        sinValue[4]) );
  FDS2L \sinValue_reg[3]  ( .CR(1'b1), .D(N39), .LD(n540), .CP(clk), .Q(
        sinValue[3]) );
  FDS2L \sinValue_reg[2]  ( .CR(1'b1), .D(N38), .LD(n540), .CP(clk), .Q(
        sinValue[2]) );
  FDS2L \sinValue_reg[1]  ( .CR(1'b1), .D(N37), .LD(n540), .CP(clk), .Q(
        sinValue[1]) );
  FDS2L \sinValue_reg[0]  ( .CR(1'b1), .D(N36), .LD(n540), .CP(clk), .Q(
        sinValue[0]) );
  FDS2L \sinValue_reg[15]  ( .CR(1'b1), .D(sValue), .LD(n540), .CP(clk), .Q(
        sinValue[15]) );
  FDS2L sValue_reg ( .CR(1'b1), .D(N57), .LD(n540), .CP(clk), .Q(sValue) );
  FJK1 \Term2_reg[18]  ( .J(n540), .K(1'b0), .CP(clk), .Q(\Term2[18] ) );
  AN2P U1719 ( .A(n342), .B(n341), .Z(n37) );
  AN2P U1720 ( .A(n303), .B(n302), .Z(n38) );
  AN2P U1721 ( .A(n261), .B(n260), .Z(n39) );
  AN2P U1722 ( .A(n246), .B(n245), .Z(n40) );
  AN2P U1723 ( .A(n327), .B(n326), .Z(n41) );
  AN2P U1724 ( .A(x[14]), .B(n47), .Z(n42) );
  NR2 U1726 ( .A(n530), .B(n498), .Z(n234) );
  EO U1727 ( .A(n525), .B(n493), .Z(n166) );
  ND2 U1728 ( .A(n236), .B(n235), .Z(n173) );
  ND2 U1729 ( .A(n232), .B(n531), .Z(n235) );
  MUX21L U1730 ( .A(n233), .B(n234), .S(n462), .Z(n236) );
  NR2 U1731 ( .A(n498), .B(n463), .Z(n232) );
  AO4 U1732 ( .A(n527), .B(n467), .C(n527), .D(n495), .Z(n179) );
  ND2 U1733 ( .A(n500), .B(n206), .Z(n153) );
  ND2 U1734 ( .A(n532), .B(n460), .Z(n206) );
  ND2 U1735 ( .A(n337), .B(n336), .Z(n165) );
  ND2 U1736 ( .A(n526), .B(n458), .Z(n336) );
  EN U1737 ( .A(n525), .B(n494), .Z(n337) );
  ND2 U1738 ( .A(n495), .B(n305), .Z(n163) );
  ND2 U1739 ( .A(n527), .B(n467), .Z(n305) );
  ND2 U1740 ( .A(n527), .B(n335), .Z(n182) );
  ND2 U1741 ( .A(n494), .B(n459), .Z(n335) );
  ND2 U1742 ( .A(n228), .B(n227), .Z(n142) );
  ND2 U1743 ( .A(n459), .B(n499), .Z(n227) );
  MUX21L U1744 ( .A(n226), .B(n499), .S(n531), .Z(n228) );
  NR2 U1745 ( .A(n499), .B(n460), .Z(n226) );
  MUX21L U1746 ( .A(n267), .B(n497), .S(n529), .Z(n269) );
  NR2 U1747 ( .A(n497), .B(n464), .Z(n267) );
  MUX21L U1748 ( .A(n498), .B(n463), .S(n530), .Z(n156) );
  MUX21L U1749 ( .A(n528), .B(n501), .S(n462), .Z(n151) );
  ND2 U1750 ( .A(n293), .B(n292), .Z(n148) );
  ND2 U1751 ( .A(n466), .B(n528), .Z(n292) );
  MUX21L U1752 ( .A(n528), .B(n291), .S(n495), .Z(n293) );
  NR2 U1753 ( .A(n527), .B(n466), .Z(n291) );
  AO4 U1754 ( .A(n494), .B(n460), .C(n526), .D(n459), .Z(n149) );
  AO7 U1755 ( .A(n526), .B(n494), .C(n468), .Z(n164) );
  AO7 U1756 ( .A(n530), .B(n498), .C(n463), .Z(n144) );
  ND2 U1757 ( .A(n464), .B(n496), .Z(n268) );
  AN2P U1758 ( .A(n528), .B(n466), .Z(n44) );
  EO U1759 ( .A(n493), .B(n463), .Z(n248) );
  EN U1760 ( .A(n525), .B(n496), .Z(n132) );
  EN U1761 ( .A(n525), .B(n467), .Z(n134) );
  EO U1762 ( .A(n524), .B(n499), .Z(n114) );
  ND2 U1763 ( .A(n231), .B(n230), .Z(n115) );
  ND2 U1764 ( .A(n459), .B(n499), .Z(n230) );
  MUX21L U1765 ( .A(n229), .B(n499), .S(n531), .Z(n231) );
  NR2 U1766 ( .A(n499), .B(n459), .Z(n229) );
  ND2 U1767 ( .A(n501), .B(n462), .Z(n111) );
  EN U1768 ( .A(n525), .B(n498), .Z(n99) );
  AO4 U1769 ( .A(n500), .B(n461), .C(n532), .D(n460), .Z(n95) );
  EO U1770 ( .A(n525), .B(n468), .Z(n106) );
  EO U1771 ( .A(n525), .B(n468), .Z(n107) );
  EO U1772 ( .A(n525), .B(n459), .Z(n108) );
  EN U1773 ( .A(n525), .B(n497), .Z(n100) );
  ND2 U1774 ( .A(n310), .B(n309), .Z(n105) );
  ND2 U1775 ( .A(n494), .B(n467), .Z(n309) );
  EN U1776 ( .A(n525), .B(n467), .Z(n310) );
  ND2 U1777 ( .A(n501), .B(n462), .Z(n93) );
  AO4 U1778 ( .A(n499), .B(n460), .C(n531), .D(n460), .Z(n81) );
  ND2 U1779 ( .A(n531), .B(n500), .Z(n212) );
  EO U1780 ( .A(n493), .B(n464), .Z(n84) );
  ND2 U1781 ( .A(n498), .B(n464), .Z(n257) );
  ND2 U1782 ( .A(n283), .B(n282), .Z(n71) );
  EN U1783 ( .A(n525), .B(n465), .Z(n282) );
  EN U1784 ( .A(n493), .B(n465), .Z(n283) );
  ND2 U1785 ( .A(n354), .B(n353), .Z(n77) );
  ND2 U1786 ( .A(n528), .B(n458), .Z(n354) );
  ND2 U1787 ( .A(n501), .B(n458), .Z(n353) );
  AO4 U1788 ( .A(n496), .B(n466), .C(n528), .D(n466), .Z(n72) );
  AO7 U1789 ( .A(n527), .B(n495), .C(n468), .Z(n75) );
  ND2 U1790 ( .A(n530), .B(n463), .Z(n258) );
  ND2 U1791 ( .A(n312), .B(n311), .Z(n73) );
  ND2 U1792 ( .A(n495), .B(n467), .Z(n311) );
  ND2 U1793 ( .A(n527), .B(n467), .Z(n312) );
  AN2P U1794 ( .A(n496), .B(n465), .Z(n45) );
  MUX21L U1795 ( .A(n459), .B(n334), .S(n495), .Z(n76) );
  ND2 U1796 ( .A(n525), .B(n459), .Z(n334) );
  AN3 U1797 ( .A(n493), .B(n458), .C(n524), .Z(n62) );
  ND2 U1798 ( .A(n496), .B(n468), .Z(n326) );
  ND2 U1799 ( .A(n527), .B(n468), .Z(n327) );
  ND2 U1800 ( .A(n529), .B(n464), .Z(n264) );
  AN2P U1801 ( .A(n501), .B(n462), .Z(n46) );
  IVP U1802 ( .A(n439), .Z(n458) );
  IVP U1803 ( .A(n475), .Z(n498) );
  IVP U1804 ( .A(n475), .Z(n500) );
  IVP U1805 ( .A(n475), .Z(n501) );
  ND2 U1806 ( .A(n193), .B(n192), .Z(n152) );
  ND2 U1807 ( .A(n189), .B(n521), .Z(n192) );
  MUX21L U1808 ( .A(n190), .B(n191), .S(n501), .Z(n193) );
  NR2 U1809 ( .A(n461), .B(n501), .Z(n189) );
  ND2 U1810 ( .A(n253), .B(n252), .Z(n157) );
  ND2 U1811 ( .A(n451), .B(n486), .Z(n252) );
  EN U1812 ( .A(n525), .B(n498), .Z(n253) );
  ND2 U1813 ( .A(n271), .B(n270), .Z(n161) );
  ND2 U1814 ( .A(n465), .B(n514), .Z(n270) );
  EN U1815 ( .A(n493), .B(n465), .Z(n271) );
  ND2 U1816 ( .A(n204), .B(n203), .Z(n170) );
  ND2 U1817 ( .A(n500), .B(n520), .Z(n203) );
  MUX21L U1818 ( .A(n520), .B(n202), .S(n461), .Z(n204) );
  NR2 U1819 ( .A(n500), .B(n520), .Z(n202) );
  ND2 U1820 ( .A(n215), .B(n214), .Z(n171) );
  ND2 U1821 ( .A(n500), .B(n518), .Z(n214) );
  MUX21L U1822 ( .A(n519), .B(n213), .S(n461), .Z(n215) );
  NR2 U1823 ( .A(n500), .B(n518), .Z(n213) );
  ND2 U1824 ( .A(n262), .B(n516), .Z(n175) );
  EO U1825 ( .A(n493), .B(n464), .Z(n262) );
  ND2 U1826 ( .A(n317), .B(n316), .Z(n180) );
  ND2 U1827 ( .A(n313), .B(n510), .Z(n316) );
  MUX21L U1828 ( .A(n314), .B(n315), .S(n494), .Z(n317) );
  NR2 U1829 ( .A(n468), .B(n495), .Z(n313) );
  IVP U1830 ( .A(n508), .Z(n531) );
  IVP U1831 ( .A(n440), .Z(n461) );
  IVP U1832 ( .A(n439), .Z(n459) );
  IVP U1833 ( .A(n508), .Z(n529) );
  IVP U1834 ( .A(n440), .Z(n463) );
  IVP U1835 ( .A(n475), .Z(n499) );
  IVP U1836 ( .A(n474), .Z(n495) );
  IVP U1837 ( .A(n441), .Z(n467) );
  IVP U1838 ( .A(n508), .Z(n530) );
  IVP U1839 ( .A(n440), .Z(n462) );
  IVP U1840 ( .A(n507), .Z(n527) );
  IVP U1841 ( .A(n507), .Z(n526) );
  IVP U1842 ( .A(n441), .Z(n468) );
  IVP U1843 ( .A(n439), .Z(n460) );
  IVP U1844 ( .A(n474), .Z(n494) );
  IVP U1845 ( .A(n507), .Z(n525) );
  IVP U1846 ( .A(n508), .Z(n528) );
  IVP U1847 ( .A(n440), .Z(n464) );
  IVP U1848 ( .A(n508), .Z(n532) );
  IVP U1849 ( .A(n440), .Z(n465) );
  AO7 U1850 ( .A(n531), .B(n488), .C(n443), .Z(n172) );
  NR2 U1851 ( .A(n532), .B(n448), .Z(n191) );
  NR2 U1852 ( .A(n531), .B(n487), .Z(n233) );
  NR2 U1853 ( .A(n527), .B(n457), .Z(n315) );
  ND3 U1854 ( .A(n251), .B(n250), .C(n249), .Z(n174) );
  ND2 U1855 ( .A(n450), .B(n486), .Z(n250) );
  ND2 U1856 ( .A(n530), .B(n486), .Z(n251) );
  ND2 U1857 ( .A(n530), .B(n450), .Z(n249) );
  ND2 U1858 ( .A(n241), .B(n240), .Z(n143) );
  ND2 U1859 ( .A(n237), .B(n517), .Z(n240) );
  MUX21L U1860 ( .A(n238), .B(n239), .S(n463), .Z(n241) );
  NR2 U1861 ( .A(n463), .B(n498), .Z(n237) );
  ND2 U1862 ( .A(n442), .B(n509), .Z(n341) );
  MUX21L U1863 ( .A(n476), .B(n340), .S(n459), .Z(n342) );
  MUX21L U1864 ( .A(n217), .B(n216), .S(n500), .Z(n154) );
  ND2 U1865 ( .A(n446), .B(n518), .Z(n216) );
  ND2 U1866 ( .A(n531), .B(n446), .Z(n217) );
  MUX21L U1867 ( .A(n488), .B(n517), .S(n460), .Z(n155) );
  MUX21L U1868 ( .A(n285), .B(n284), .S(n496), .Z(n178) );
  ND2 U1869 ( .A(n529), .B(n455), .Z(n285) );
  ND2 U1870 ( .A(n528), .B(n465), .Z(n284) );
  MUX21L U1871 ( .A(n208), .B(n207), .S(n532), .Z(n140) );
  ND2 U1872 ( .A(n460), .B(n489), .Z(n208) );
  ND2 U1873 ( .A(n500), .B(n460), .Z(n207) );
  IVP U1874 ( .A(n474), .Z(n496) );
  IVP U1875 ( .A(n474), .Z(n497) );
  IVP U1876 ( .A(n440), .Z(n466) );
  AO7 U1877 ( .A(n497), .B(n515), .C(n453), .Z(n158) );
  AO7 U1878 ( .A(n497), .B(n522), .C(n463), .Z(n168) );
  NR2 U1879 ( .A(n530), .B(n487), .Z(n239) );
  NR2 U1880 ( .A(n468), .B(n479), .Z(n181) );
  ND2 U1881 ( .A(n467), .B(n482), .Z(n303) );
  ND2 U1882 ( .A(n467), .B(n511), .Z(n302) );
  ND2 U1883 ( .A(n221), .B(n445), .Z(n141) );
  ND2 U1884 ( .A(n531), .B(n499), .Z(n221) );
  ND2 U1885 ( .A(n186), .B(n185), .Z(n138) );
  ND2 U1886 ( .A(n462), .B(n492), .Z(n185) );
  MUX21L U1887 ( .A(n492), .B(n184), .S(n532), .Z(n186) );
  NR2 U1888 ( .A(n462), .B(n492), .Z(n184) );
  ND2 U1889 ( .A(n200), .B(n199), .Z(n139) );
  ND2 U1890 ( .A(n461), .B(n490), .Z(n199) );
  MUX21L U1891 ( .A(n198), .B(n532), .S(n461), .Z(n200) );
  NR2 U1892 ( .A(n532), .B(n490), .Z(n198) );
  MUX21L U1893 ( .A(n512), .B(n482), .S(n466), .Z(n162) );
  MUX21L U1894 ( .A(n484), .B(n515), .S(n464), .Z(n160) );
  MUX21L U1895 ( .A(n197), .B(n448), .S(n532), .Z(n169) );
  ND2 U1896 ( .A(n448), .B(n490), .Z(n197) );
  ND2 U1897 ( .A(n188), .B(n187), .Z(n125) );
  ND2 U1898 ( .A(n532), .B(n449), .Z(n187) );
  EN U1899 ( .A(n493), .B(n462), .Z(n188) );
  ND2 U1900 ( .A(n499), .B(n444), .Z(n225) );
  ND2 U1901 ( .A(n461), .B(n489), .Z(n205) );
  ND2 U1902 ( .A(n344), .B(n343), .Z(n136) );
  ND2 U1903 ( .A(n494), .B(n442), .Z(n343) );
  EO U1904 ( .A(n524), .B(n458), .Z(n344) );
  ND2 U1905 ( .A(n453), .B(n485), .Z(n145) );
  ND2 U1906 ( .A(n196), .B(n195), .Z(n126) );
  ND2 U1907 ( .A(n461), .B(n491), .Z(n195) );
  MUX21L U1908 ( .A(n491), .B(n194), .S(n532), .Z(n196) );
  NR2 U1909 ( .A(n461), .B(n491), .Z(n194) );
  MUX21L U1910 ( .A(n328), .B(n525), .S(n459), .Z(n135) );
  ND2 U1911 ( .A(n527), .B(n478), .Z(n328) );
  AO7 U1912 ( .A(n529), .B(n496), .C(n454), .Z(n131) );
  ND2 U1913 ( .A(n450), .B(n516), .Z(n247) );
  MUX21L U1914 ( .A(n286), .B(n496), .S(n465), .Z(n133) );
  ND2 U1915 ( .A(n495), .B(n513), .Z(n286) );
  ND2 U1916 ( .A(n308), .B(n307), .Z(n121) );
  ND2 U1917 ( .A(n481), .B(n511), .Z(n307) );
  MUX21L U1918 ( .A(n481), .B(n306), .S(n467), .Z(n308) );
  ND2 U1919 ( .A(n244), .B(n243), .Z(n116) );
  ND2 U1920 ( .A(n530), .B(n487), .Z(n243) );
  MUX21L U1921 ( .A(n242), .B(n449), .S(n530), .Z(n244) );
  ND2 U1922 ( .A(n211), .B(n210), .Z(n113) );
  ND2 U1923 ( .A(n461), .B(n500), .Z(n210) );
  MUX21L U1924 ( .A(n209), .B(n519), .S(n500), .Z(n211) );
  NR2 U1925 ( .A(n460), .B(n519), .Z(n209) );
  ND2 U1926 ( .A(n290), .B(n289), .Z(n120) );
  AO6 U1927 ( .A(n497), .B(n455), .C(n288), .Z(n290) );
  MUX21L U1928 ( .A(n287), .B(n513), .S(n495), .Z(n289) );
  NR2 U1929 ( .A(n528), .B(n465), .Z(n288) );
  ND2 U1930 ( .A(n347), .B(n346), .Z(n123) );
  ND2 U1931 ( .A(n526), .B(n493), .Z(n346) );
  MUX21L U1932 ( .A(n345), .B(n442), .S(n493), .Z(n347) );
  NR2 U1933 ( .A(n526), .B(n441), .Z(n345) );
  MUX21L U1934 ( .A(n201), .B(n447), .S(n500), .Z(n112) );
  ND2 U1935 ( .A(n447), .B(n521), .Z(n201) );
  ND2 U1936 ( .A(n274), .B(n273), .Z(n119) );
  ND2 U1937 ( .A(n529), .B(n454), .Z(n273) );
  MUX21L U1938 ( .A(n484), .B(n272), .S(n465), .Z(n274) );
  NR2 U1939 ( .A(n529), .B(n484), .Z(n272) );
  ND2 U1940 ( .A(n330), .B(n329), .Z(n122) );
  ND2 U1941 ( .A(n478), .B(n510), .Z(n330) );
  ND2 U1942 ( .A(n459), .B(n478), .Z(n329) );
  AO7 U1943 ( .A(n497), .B(n464), .C(n515), .Z(n118) );
  ND2 U1944 ( .A(n220), .B(n219), .Z(n96) );
  ND2 U1945 ( .A(n445), .B(n517), .Z(n219) );
  MUX21L U1946 ( .A(n488), .B(n218), .S(n460), .Z(n220) );
  ND2 U1947 ( .A(n278), .B(n277), .Z(n103) );
  AO6 U1948 ( .A(n496), .B(n455), .C(n276), .Z(n278) );
  MUX21L U1949 ( .A(n275), .B(n514), .S(n496), .Z(n277) );
  NR2 U1950 ( .A(n529), .B(n465), .Z(n276) );
  AO7 U1951 ( .A(n530), .B(n449), .C(n498), .Z(n98) );
  NR2 U1952 ( .A(n458), .B(n509), .Z(n348) );
  NR2 U1953 ( .A(n526), .B(n475), .Z(n349) );
  NR2 U1954 ( .A(n495), .B(n512), .Z(n295) );
  ND2 U1955 ( .A(n298), .B(n297), .Z(n104) );
  NR2 U1956 ( .A(n296), .B(n295), .Z(n298) );
  MUX21L U1957 ( .A(n294), .B(n466), .S(n528), .Z(n297) );
  NR2 U1958 ( .A(n496), .B(n456), .Z(n296) );
  ND2 U1959 ( .A(n224), .B(n223), .Z(n97) );
  ND2 U1960 ( .A(n531), .B(n444), .Z(n224) );
  ND2 U1961 ( .A(n499), .B(n444), .Z(n223) );
  ND2 U1962 ( .A(n352), .B(n351), .Z(n109) );
  NR2 U1963 ( .A(n350), .B(n349), .Z(n352) );
  MUX21L U1964 ( .A(n348), .B(n458), .S(n494), .Z(n351) );
  NR2 U1965 ( .A(n525), .B(n441), .Z(n350) );
  NR2 U1966 ( .A(n466), .B(n483), .Z(n294) );
  NR2 U1967 ( .A(n497), .B(n452), .Z(n259) );
  ND2 U1968 ( .A(n256), .B(n255), .Z(n82) );
  ND2 U1969 ( .A(n498), .B(n451), .Z(n255) );
  MUX21L U1970 ( .A(n254), .B(n452), .S(n530), .Z(n256) );
  NR2 U1971 ( .A(n498), .B(n451), .Z(n254) );
  ND2 U1972 ( .A(n463), .B(n516), .Z(n245) );
  EN U1973 ( .A(n493), .B(n463), .Z(n246) );
  ND2 U1974 ( .A(n266), .B(n265), .Z(n102) );
  ND2 U1975 ( .A(n464), .B(n485), .Z(n265) );
  ND2 U1976 ( .A(n529), .B(n485), .Z(n266) );
  ND2 U1977 ( .A(n497), .B(n452), .Z(n260) );
  MUX21L U1978 ( .A(n259), .B(n453), .S(n529), .Z(n261) );
  ND2 U1979 ( .A(n320), .B(n319), .Z(n88) );
  ND2 U1980 ( .A(n526), .B(n480), .Z(n319) );
  MUX21L U1981 ( .A(n480), .B(n318), .S(n468), .Z(n320) );
  NR2 U1982 ( .A(n527), .B(n479), .Z(n318) );
  ND2 U1983 ( .A(n333), .B(n332), .Z(n90) );
  ND2 U1984 ( .A(n526), .B(n477), .Z(n332) );
  MUX21L U1985 ( .A(n477), .B(n331), .S(n460), .Z(n333) );
  NR2 U1986 ( .A(n526), .B(n477), .Z(n331) );
  ND2 U1987 ( .A(n325), .B(n324), .Z(n89) );
  ND2 U1988 ( .A(n528), .B(n494), .Z(n324) );
  MUX21L U1989 ( .A(n323), .B(n457), .S(n494), .Z(n325) );
  NR2 U1990 ( .A(n526), .B(n457), .Z(n323) );
  ND3 U1991 ( .A(n489), .B(n521), .C(n447), .Z(n94) );
  ND2 U1992 ( .A(n300), .B(n299), .Z(n86) );
  ND2 U1993 ( .A(n456), .B(n512), .Z(n299) );
  EO U1994 ( .A(n493), .B(n467), .Z(n300) );
  MUX21L U1995 ( .A(n339), .B(n338), .S(n459), .Z(n91) );
  ND2 U1996 ( .A(n476), .B(n509), .Z(n338) );
  ND2 U1997 ( .A(n526), .B(n494), .Z(n339) );
  ND3 U1998 ( .A(n281), .B(n280), .C(n279), .Z(n85) );
  ND2 U1999 ( .A(n483), .B(n513), .Z(n280) );
  ND2 U2000 ( .A(n465), .B(n514), .Z(n281) );
  ND2 U2001 ( .A(n465), .B(n483), .Z(n279) );
  MUX21L U2002 ( .A(n481), .B(n304), .S(n467), .Z(n87) );
  ND2 U2003 ( .A(n482), .B(n511), .Z(n304) );
  ND2 U2004 ( .A(n322), .B(n321), .Z(n74) );
  ND2 U2005 ( .A(n468), .B(n510), .Z(n321) );
  EN U2006 ( .A(n493), .B(n468), .Z(n322) );
  ND2 U2007 ( .A(n222), .B(n445), .Z(n67) );
  ND2 U2008 ( .A(n531), .B(n499), .Z(n222) );
  IVP U2009 ( .A(n503), .Z(n474) );
  IVP U2010 ( .A(n534), .Z(n508) );
  IVP U2011 ( .A(n470), .Z(n440) );
  MUX21L U2012 ( .A(n416), .B(n415), .S(n430), .Z(n424) );
  NR3 U2013 ( .A(n436), .B(n38), .C(n432), .Z(n415) );
  NR2 U2014 ( .A(n436), .B(n37), .Z(n416) );
  MUX21L U2015 ( .A(n420), .B(n419), .S(n433), .Z(n422) );
  AN3 U2016 ( .A(n429), .B(n148), .C(n436), .Z(n420) );
  ND2 U2017 ( .A(n269), .B(n268), .Z(n147) );
  MUX21L U2018 ( .A(n418), .B(n417), .S(n436), .Z(n423) );
  NR2 U2019 ( .A(n430), .B(n426), .Z(n417) );
  IVP U2020 ( .A(n149), .Z(n426) );
  MUX21L U2021 ( .A(n370), .B(n369), .S(n429), .Z(n373) );
  AN3 U2022 ( .A(n128), .B(n432), .C(n436), .Z(n370) );
  AN3 U2023 ( .A(n125), .B(n432), .C(n436), .Z(n369) );
  MUX21L U2024 ( .A(n225), .B(n443), .S(n531), .Z(n128) );
  MUX21L U2025 ( .A(n402), .B(n403), .S(n430), .Z(n411) );
  NR2 U2026 ( .A(n437), .B(n425), .Z(n403) );
  NR3 U2027 ( .A(n437), .B(n39), .C(n433), .Z(n402) );
  IVP U2028 ( .A(n81), .Z(n425) );
  MUX21L U2029 ( .A(n407), .B(n406), .S(n430), .Z(n408) );
  AN3 U2030 ( .A(n436), .B(n458), .C(n432), .Z(n407) );
  ND2 U2031 ( .A(n501), .B(n462), .Z(n79) );
  MUX21L U2032 ( .A(n357), .B(n358), .S(n433), .Z(n366) );
  NR2 U2033 ( .A(n437), .B(n62), .Z(n358) );
  MUX21L U2034 ( .A(n359), .B(n360), .S(n433), .Z(n365) );
  ND2 U2035 ( .A(n501), .B(n462), .Z(n66) );
  MUX21L U2036 ( .A(n376), .B(n56), .S(n429), .Z(n381) );
  ND2 U2037 ( .A(n501), .B(n462), .Z(n56) );
  MUX21L U2038 ( .A(n394), .B(n395), .S(n433), .Z(n397) );
  AO4 U2039 ( .A(n496), .B(n466), .C(n528), .D(n466), .Z(n61) );
  MUX21L U2040 ( .A(n384), .B(n385), .S(n433), .Z(n386) );
  NR2 U2041 ( .A(n430), .B(n41), .Z(n385) );
  AO4 U2042 ( .A(n495), .B(n466), .C(n528), .D(n466), .Z(n54) );
  MUX21L U2043 ( .A(n52), .B(n51), .S(n430), .Z(n412) );
  ND2 U2044 ( .A(n264), .B(n263), .Z(n52) );
  ND2 U2045 ( .A(n501), .B(n462), .Z(n51) );
  ND2 U2046 ( .A(n497), .B(n464), .Z(n263) );
  EN U2047 ( .A(n432), .B(n430), .Z(n414) );
  MUX21L U2048 ( .A(n382), .B(n383), .S(n430), .Z(n387) );
  NR2 U2049 ( .A(n437), .B(n433), .Z(n383) );
  EN U2050 ( .A(n436), .B(n430), .Z(n413) );
  ND2 U2051 ( .A(n49), .B(n437), .Z(n389) );
  ND2 U2052 ( .A(n301), .B(n456), .Z(n49) );
  ND2 U2053 ( .A(n527), .B(n495), .Z(n301) );
  ND2 U2054 ( .A(n429), .B(n46), .Z(n356) );
  ND2 U2055 ( .A(n433), .B(n429), .Z(n388) );
  ND2 U2056 ( .A(n438), .B(n433), .Z(n355) );
  IVP U2057 ( .A(n469), .Z(n470) );
  IVP U2058 ( .A(n502), .Z(n503) );
  IVP U2059 ( .A(n533), .Z(n534) );
  IVP U2060 ( .A(n469), .Z(n472) );
  IVP U2061 ( .A(n442), .Z(n473) );
  IVP U2062 ( .A(n476), .Z(n505) );
  IVP U2063 ( .A(n431), .Z(n434) );
  IVP U2064 ( .A(n427), .Z(n429) );
  IVP U2065 ( .A(n431), .Z(n432) );
  IVP U2066 ( .A(n427), .Z(n428) );
  IVP U2067 ( .A(n502), .Z(n504) );
  IVP U2068 ( .A(n477), .Z(n506) );
  IVP U2069 ( .A(n469), .Z(n471) );
  MUX21L U2070 ( .A(n371), .B(n372), .S(n429), .Z(n374) );
  NR3 U2071 ( .A(n437), .B(n532), .C(n433), .Z(n372) );
  AN3 U2072 ( .A(n129), .B(n435), .C(n432), .Z(n371) );
  ND2 U2073 ( .A(n248), .B(n247), .Z(n129) );
  IVP U2074 ( .A(n431), .Z(n433) );
  IVP U2075 ( .A(n435), .Z(n438) );
  IVP U2076 ( .A(n427), .Z(n430) );
  IVP U2077 ( .A(n435), .Z(n436) );
  MUX21L U2078 ( .A(n367), .B(n368), .S(n433), .Z(n375) );
  AN3 U2079 ( .A(n127), .B(n428), .C(n436), .Z(n367) );
  AN3 U2080 ( .A(n126), .B(n435), .C(n428), .Z(n368) );
  MUX21L U2081 ( .A(n461), .B(n205), .S(n532), .Z(n127) );
  ND2 U2082 ( .A(n432), .B(n427), .Z(n421) );
  IVP U2083 ( .A(n435), .Z(n437) );
  AO2 U2084 ( .A(n401), .B(n433), .C(n400), .D(n433), .Z(n409) );
  NR2 U2085 ( .A(n437), .B(n427), .Z(n400) );
  NR2 U2086 ( .A(n437), .B(n40), .Z(n401) );
  MUX21L U2087 ( .A(n405), .B(n404), .S(n430), .Z(n410) );
  AN3 U2088 ( .A(n80), .B(n431), .C(n436), .Z(n404) );
  AN3 U2089 ( .A(n82), .B(n431), .C(n436), .Z(n405) );
  ND2 U2090 ( .A(n212), .B(n446), .Z(n80) );
  MUX21L U2091 ( .A(n361), .B(n362), .S(n433), .Z(n364) );
  NR2 U2092 ( .A(n437), .B(n427), .Z(n362) );
  ND2 U2093 ( .A(n258), .B(n257), .Z(n68) );
  ND4 U2094 ( .A(n69), .B(n427), .C(n431), .D(n435), .Z(n363) );
  AO7 U2095 ( .A(n529), .B(n497), .C(n464), .Z(n69) );
  MUX21L U2096 ( .A(n377), .B(n435), .S(n430), .Z(n380) );
  AN3 U2097 ( .A(n493), .B(n458), .C(n524), .Z(n57) );
  MUX21L U2098 ( .A(n392), .B(n393), .S(n433), .Z(n398) );
  AN3 U2099 ( .A(n64), .B(n427), .C(n436), .Z(n392) );
  ND2 U2100 ( .A(n443), .B(n476), .Z(n64) );
  MUX21L U2101 ( .A(n390), .B(n391), .S(n433), .Z(n399) );
  NR2 U2102 ( .A(n437), .B(n427), .Z(n390) );
  AN3 U2103 ( .A(n493), .B(n458), .C(n525), .Z(n60) );
  ND4 U2104 ( .A(n63), .B(n433), .C(n427), .D(n435), .Z(n396) );
  AO7 U2105 ( .A(n526), .B(n494), .C(n468), .Z(n63) );
  ND3 U2106 ( .A(n58), .B(n435), .C(n431), .Z(n378) );
  AO7 U2107 ( .A(n529), .B(n497), .C(n464), .Z(n58) );
  ND2 U2108 ( .A(n429), .B(n431), .Z(n379) );
  ND2 U2109 ( .A(n529), .B(n454), .Z(n177) );
  ND4 U2110 ( .A(n424), .B(n423), .C(n422), .D(n421), .Z(n150) );
  ND3 U2111 ( .A(n375), .B(n374), .C(n373), .Z(n130) );
  ND4 U2112 ( .A(n411), .B(n410), .C(n409), .D(n408), .Z(n83) );
  ND4 U2113 ( .A(n366), .B(n365), .C(n364), .D(n363), .Z(n70) );
  ND4 U2114 ( .A(n399), .B(n398), .C(n397), .D(n396), .Z(n65) );
  ND4 U2115 ( .A(n381), .B(n380), .C(n379), .D(n378), .Z(n59) );
  ND3 U2116 ( .A(n414), .B(n413), .C(n412), .Z(n53) );
  ND2 U2117 ( .A(n387), .B(n386), .Z(n55) );
  AO7 U2118 ( .A(n427), .B(n389), .C(n388), .Z(n50) );
  ND4 U2119 ( .A(n437), .B(n433), .C(n430), .D(n46), .Z(n48) );
  NR2 U2120 ( .A(n356), .B(n355), .Z(n47) );
  EN U2121 ( .A(n35), .B(x[15]), .Z(N57) );
  ND2 U2122 ( .A(x[14]), .B(func), .Z(n35) );
  IVP U2123 ( .A(reset), .Z(n540) );
  MUX21H U2124 ( .A(n50), .B(n48), .S(x[14]), .Z(N9) );
  MUX21H U2125 ( .A(n55), .B(n53), .S(x[14]), .Z(N10) );
  MUX21H U2126 ( .A(n65), .B(n59), .S(x[14]), .Z(N11) );
  MUX81P U2127 ( .D0(n77), .D1(n73), .D2(n75), .D3(n71), .D4(n76), .D5(n72), 
        .D6(n74), .D7(n45), .A(n429), .B(n434), .C(n437), .Z(n78) );
  MUX21H U2128 ( .A(n78), .B(n70), .S(x[14]), .Z(N12) );
  MUX81P U2129 ( .D0(n91), .D1(n87), .D2(n89), .D3(n85), .D4(n90), .D5(n86), 
        .D6(n88), .D7(n84), .A(n429), .B(n434), .C(n438), .Z(n92) );
  MUX21H U2130 ( .A(n92), .B(n83), .S(x[14]), .Z(N13) );
  MUX81P U2131 ( .D0(n100), .D1(n96), .D2(n98), .D3(n94), .D4(n99), .D5(n95), 
        .D6(n97), .D7(n93), .A(n429), .B(n434), .C(n438), .Z(n101) );
  MUX81P U2132 ( .D0(n109), .D1(n105), .D2(n107), .D3(n103), .D4(n108), .D5(
        n104), .D6(n106), .D7(n102), .A(n429), .B(n434), .C(n438), .Z(n110) );
  MUX21H U2133 ( .A(n110), .B(n101), .S(x[14]), .Z(N14) );
  MUX81P U2134 ( .D0(n522), .D1(n114), .D2(n116), .D3(n112), .D4(n522), .D5(
        n113), .D6(n115), .D7(n111), .A(n429), .B(n434), .C(n438), .Z(n117) );
  MUX81P U2135 ( .D0(n123), .D1(n121), .D2(n479), .D3(n119), .D4(n122), .D5(
        n120), .D6(n480), .D7(n118), .A(n429), .B(n434), .C(n438), .Z(n124) );
  MUX21H U2136 ( .A(n124), .B(n117), .S(x[14]), .Z(N15) );
  MUX81P U2137 ( .D0(n136), .D1(n134), .D2(n523), .D3(n132), .D4(n135), .D5(
        n133), .D6(n523), .D7(n131), .A(n429), .B(n434), .C(n438), .Z(n137) );
  MUX21H U2138 ( .A(n137), .B(n130), .S(x[14]), .Z(N16) );
  MUX81P U2139 ( .D0(n145), .D1(n141), .D2(n143), .D3(n139), .D4(n144), .D5(
        n140), .D6(n142), .D7(n138), .A(n429), .B(n434), .C(n438), .Z(n146) );
  MUX21H U2140 ( .A(n150), .B(n146), .S(x[14]), .Z(N17) );
  MUX81P U2141 ( .D0(n158), .D1(n154), .D2(n156), .D3(n152), .D4(n157), .D5(
        n153), .D6(n155), .D7(n151), .A(n429), .B(n434), .C(n438), .Z(n159) );
  MUX81P U2142 ( .D0(n166), .D1(n163), .D2(n463), .D3(n161), .D4(n165), .D5(
        n162), .D6(n164), .D7(n160), .A(n429), .B(n434), .C(n438), .Z(n167) );
  MUX21H U2143 ( .A(n167), .B(n159), .S(x[14]), .Z(N18) );
  MUX81P U2144 ( .D0(n175), .D1(n171), .D2(n173), .D3(n169), .D4(n174), .D5(
        n170), .D6(n172), .D7(n168), .A(n429), .B(n434), .C(n438), .Z(n176) );
  MUX81P U2145 ( .D0(n523), .D1(n179), .D2(n181), .D3(n178), .D4(n182), .D5(
        n44), .D6(n180), .D7(n177), .A(n428), .B(n434), .C(n438), .Z(n183) );
  AN2P U2146 ( .A(n524), .B(n458), .Z(n190) );
  AN2P U2147 ( .A(n525), .B(n493), .Z(n218) );
  AN2P U2148 ( .A(n525), .B(n493), .Z(n238) );
  AN2P U2149 ( .A(n493), .B(n458), .Z(n242) );
  AN2P U2150 ( .A(n525), .B(n458), .Z(n275) );
  AN2P U2151 ( .A(n525), .B(n458), .Z(n287) );
  AN2P U2152 ( .A(n525), .B(n493), .Z(n306) );
  AN2P U2153 ( .A(n524), .B(n458), .Z(n314) );
  AN2P U2154 ( .A(n524), .B(n493), .Z(n340) );
  AN2P U2155 ( .A(n436), .B(n428), .Z(n357) );
  AN2P U2156 ( .A(n67), .B(n428), .Z(n359) );
  AN2P U2157 ( .A(n66), .B(n428), .Z(n360) );
  AN2P U2158 ( .A(n436), .B(n68), .Z(n361) );
  AN2P U2159 ( .A(n436), .B(n432), .Z(n376) );
  AN2P U2160 ( .A(n432), .B(n57), .Z(n377) );
  AN2P U2161 ( .A(n436), .B(n432), .Z(n382) );
  AN2P U2162 ( .A(n428), .B(n54), .Z(n384) );
  AN2P U2163 ( .A(n60), .B(n428), .Z(n391) );
  AN2P U2164 ( .A(n62), .B(n436), .Z(n393) );
  AN2P U2165 ( .A(n61), .B(n428), .Z(n394) );
  AN2P U2166 ( .A(n436), .B(n428), .Z(n395) );
  AN2P U2167 ( .A(n79), .B(n432), .Z(n406) );
  AN2P U2168 ( .A(n508), .B(n432), .Z(n418) );
  AN2P U2169 ( .A(n147), .B(n436), .Z(n419) );
  IVA U2170 ( .A(x[13]), .Z(n427) );
  IVP U2171 ( .A(x[12]), .Z(n431) );
  IVA U2172 ( .A(x[11]), .Z(n435) );
  IVA U2173 ( .A(n470), .Z(n439) );
  IVA U2174 ( .A(n470), .Z(n441) );
  IVA U2175 ( .A(n470), .Z(n442) );
  IVA U2176 ( .A(n471), .Z(n443) );
  IVA U2177 ( .A(n471), .Z(n444) );
  IVA U2178 ( .A(n471), .Z(n445) );
  IVA U2179 ( .A(n471), .Z(n446) );
  IVA U2180 ( .A(n471), .Z(n447) );
  IVA U2181 ( .A(n472), .Z(n448) );
  IVA U2182 ( .A(n472), .Z(n449) );
  IVA U2183 ( .A(n472), .Z(n450) );
  IVA U2184 ( .A(n472), .Z(n451) );
  IVA U2185 ( .A(n472), .Z(n452) );
  IVA U2186 ( .A(n473), .Z(n453) );
  IVA U2187 ( .A(n473), .Z(n454) );
  IVA U2188 ( .A(n473), .Z(n455) );
  IVA U2189 ( .A(n473), .Z(n456) );
  IVA U2190 ( .A(n473), .Z(n457) );
  IVP U2191 ( .A(x[10]), .Z(n469) );
  IVA U2192 ( .A(n503), .Z(n475) );
  IVA U2193 ( .A(n503), .Z(n476) );
  IVA U2194 ( .A(n503), .Z(n477) );
  IVA U2195 ( .A(n504), .Z(n478) );
  IVA U2196 ( .A(n504), .Z(n479) );
  IVA U2197 ( .A(n504), .Z(n480) );
  IVA U2198 ( .A(n504), .Z(n481) );
  IVA U2199 ( .A(n504), .Z(n482) );
  IVA U2200 ( .A(n505), .Z(n483) );
  IVA U2201 ( .A(n505), .Z(n484) );
  IVA U2202 ( .A(n505), .Z(n485) );
  IVA U2203 ( .A(n505), .Z(n486) );
  IVA U2204 ( .A(n505), .Z(n487) );
  IVA U2205 ( .A(n506), .Z(n488) );
  IVA U2206 ( .A(n506), .Z(n489) );
  IVA U2207 ( .A(n506), .Z(n490) );
  IVA U2208 ( .A(n506), .Z(n491) );
  IVA U2209 ( .A(n506), .Z(n492) );
  IVP U2210 ( .A(x[9]), .Z(n502) );
  IVA U2211 ( .A(n534), .Z(n507) );
  IVA U2212 ( .A(n535), .Z(n509) );
  IVA U2213 ( .A(n535), .Z(n510) );
  IVA U2214 ( .A(n535), .Z(n511) );
  IVA U2215 ( .A(n536), .Z(n512) );
  IVA U2216 ( .A(n536), .Z(n513) );
  IVA U2217 ( .A(n536), .Z(n514) );
  IVA U2218 ( .A(n537), .Z(n515) );
  IVA U2219 ( .A(n537), .Z(n516) );
  IVA U2220 ( .A(n537), .Z(n517) );
  IVA U2221 ( .A(n538), .Z(n518) );
  IVA U2222 ( .A(n538), .Z(n519) );
  IVA U2223 ( .A(n538), .Z(n520) );
  IVA U2224 ( .A(n539), .Z(n521) );
  IVA U2225 ( .A(n539), .Z(n522) );
  IVA U2226 ( .A(n539), .Z(n523) );
  IV U2227 ( .A(n507), .Z(n524) );
  IVA U2228 ( .A(x[8]), .Z(n533) );
  IVA U2229 ( .A(n533), .Z(n535) );
  IVA U2230 ( .A(n533), .Z(n536) );
  IVA U2231 ( .A(n509), .Z(n537) );
  IVA U2232 ( .A(n511), .Z(n538) );
  IVA U2233 ( .A(n510), .Z(n539) );
  IVP U2234 ( .A(n474), .Z(n493) );
  MUX21H U2235 ( .A(n183), .B(n176), .S(x[14]), .Z(N19) );
  EO U2236 ( .A(Term1[25]), .B(\add_29/carry[14] ), .Z(N50) );
  AN2 U2237 ( .A(\add_29/carry[13] ), .B(Term1[24]), .Z(\add_29/carry[14] ) );
  EO U2238 ( .A(Term1[24]), .B(\add_29/carry[13] ), .Z(N49) );
  AN2 U2239 ( .A(\add_29/carry[12] ), .B(Term1[23]), .Z(\add_29/carry[13] ) );
  EO U2240 ( .A(Term1[23]), .B(\add_29/carry[12] ), .Z(N48) );
  AN2 U2241 ( .A(\add_29/carry[11] ), .B(Term1[22]), .Z(\add_29/carry[12] ) );
  EO U2242 ( .A(Term1[22]), .B(\add_29/carry[11] ), .Z(N47) );
  AN2 U2243 ( .A(\add_29/carry[10] ), .B(Term1[21]), .Z(\add_29/carry[11] ) );
  EO U2244 ( .A(Term1[21]), .B(\add_29/carry[10] ), .Z(N46) );
  AN2 U2245 ( .A(\add_29/carry[9] ), .B(Term1[20]), .Z(\add_29/carry[10] ) );
  EO U2246 ( .A(Term1[20]), .B(\add_29/carry[9] ), .Z(N45) );
  AN2 U2247 ( .A(\add_29/carry[8] ), .B(Term1[19]), .Z(\add_29/carry[9] ) );
  EO U2248 ( .A(Term1[19]), .B(\add_29/carry[8] ), .Z(N44) );
  AN2 U2249 ( .A(\add_29/carry[7] ), .B(Term1[18]), .Z(\add_29/carry[8] ) );
  EO U2250 ( .A(Term1[18]), .B(\add_29/carry[7] ), .Z(N43) );
  AN2 U2251 ( .A(\add_29/carry[6] ), .B(Term1[17]), .Z(\add_29/carry[7] ) );
  EO U2252 ( .A(Term1[17]), .B(\add_29/carry[6] ), .Z(N42) );
  AN2 U2253 ( .A(\add_29/carry[5] ), .B(Term1[16]), .Z(\add_29/carry[6] ) );
  EO U2254 ( .A(Term1[16]), .B(\add_29/carry[5] ), .Z(N41) );
  AN2 U2255 ( .A(\add_29/carry[4] ), .B(Term1[15]), .Z(\add_29/carry[5] ) );
  EO U2256 ( .A(Term1[15]), .B(\add_29/carry[4] ), .Z(N40) );
  AN2 U2257 ( .A(\add_29/carry[3] ), .B(Term1[14]), .Z(\add_29/carry[4] ) );
  EO U2258 ( .A(Term1[14]), .B(\add_29/carry[3] ), .Z(N39) );
  AN2 U2259 ( .A(\add_29/carry[2] ), .B(Term1[13]), .Z(\add_29/carry[3] ) );
  EO U2260 ( .A(Term1[13]), .B(\add_29/carry[2] ), .Z(N38) );
  AN2 U2261 ( .A(\add_29/carry[1] ), .B(Term1[12]), .Z(\add_29/carry[2] ) );
  EO U2262 ( .A(Term1[12]), .B(\add_29/carry[1] ), .Z(N37) );
  AN2 U2263 ( .A(\Term2[18] ), .B(Term1[11]), .Z(\add_29/carry[1] ) );
  EO U2264 ( .A(Term1[11]), .B(\Term2[18] ), .Z(N36) );
endmodule

