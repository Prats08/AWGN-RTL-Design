
module Taus_0 ( clk, reset, Tout );
  output [31:0] Tout;
  input clk, reset;
  wire   N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N145, N183,
         N184, N185, N236, N238, n75, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n8, n14, n15, n21, n22, n37, n38, n39, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92;
  wire   [31:0] s0;
  wire   [31:0] b0;
  wire   [31:0] s1;
  wire   [31:0] b1;
  wire   [31:0] s2;
  wire   [31:0] b2;

  OR2 U182 ( .A(b2[2]), .B(reset), .Z(N238) );
  OR2 U183 ( .A(b2[0]), .B(reset), .Z(N236) );
  OR2 U184 ( .A(b1[2]), .B(reset), .Z(N185) );
  OR2 U185 ( .A(b1[1]), .B(reset), .Z(N184) );
  OR2 U186 ( .A(b1[0]), .B(reset), .Z(N183) );
  OR2 U187 ( .A(b0[1]), .B(reset), .Z(N145) );
  FDS2 \b0_reg[1]  ( .CR(n85), .D(n61), .CP(clk), .Q(b0[1]) );
  FDS2 \b1_reg[1]  ( .CR(n82), .D(n41), .CP(clk), .Q(b1[1]) );
  FDS2 \b1_reg[2]  ( .CR(n82), .D(n39), .CP(clk), .Q(b1[2]) );
  FDS2 \b1_reg[0]  ( .CR(n81), .D(n38), .CP(clk), .Q(b1[0]) );
  FDS2 \b2_reg[0]  ( .CR(n76), .D(n44), .CP(clk), .Q(b2[0]) );
  FDS2 \b2_reg[2]  ( .CR(n74), .D(n8), .CP(clk), .Q(b2[2]) );
  FDS2L \Tout_reg[11]  ( .CR(1'b1), .D(N119), .LD(n76), .CP(clk), .Q(Tout[11])
         );
  FDS2L \Tout_reg[4]  ( .CR(1'b1), .D(N126), .LD(n74), .CP(clk), .Q(Tout[4])
         );
  FDS2L \Tout_reg[2]  ( .CR(1'b1), .D(N128), .LD(n74), .CP(clk), .Q(Tout[2])
         );
  FDS2 \s0_reg[0]  ( .CR(b0[0]), .D(n84), .CP(clk), .Q(s0[0]) );
  FD1 \s0_reg[1]  ( .D(N145), .CP(clk), .Q(s0[1]) );
  FDS2 \s0_reg[5]  ( .CR(b0[5]), .D(n87), .CP(clk), .Q(s0[5]) );
  FDS2 \s0_reg[22]  ( .CR(n86), .D(s0[10]), .CP(clk), .Q(s0[22]) );
  FDS2 \s0_reg[4]  ( .CR(b0[4]), .D(n86), .CP(clk), .Q(s0[4]) );
  FDS2 \s0_reg[21]  ( .CR(n86), .D(s0[9]), .CP(clk), .Q(s0[21]) );
  FDS2 \s0_reg[3]  ( .CR(b0[3]), .D(n85), .CP(clk), .Q(s0[3]) );
  FDS2 \s0_reg[20]  ( .CR(n85), .D(s0[8]), .CP(clk), .Q(s0[20]) );
  FDS2 \s0_reg[2]  ( .CR(b0[2]), .D(n85), .CP(clk), .Q(s0[2]) );
  FDS2 \s0_reg[13]  ( .CR(n88), .D(s0[1]), .CP(clk), .Q(s0[13]) );
  FDS2 \s0_reg[25]  ( .CR(n88), .D(s0[13]), .CP(clk), .Q(s0[25]) );
  FDS2 \s0_reg[19]  ( .CR(n88), .D(s0[7]), .CP(clk), .Q(s0[19]) );
  FDS2 \s0_reg[31]  ( .CR(n88), .D(s0[19]), .CP(clk), .Q(s0[31]) );
  FDS2 \s0_reg[12]  ( .CR(b0[12]), .D(n87), .CP(clk), .Q(s0[12]) );
  FDS2 \s0_reg[24]  ( .CR(n87), .D(s0[12]), .CP(clk), .Q(s0[24]) );
  FDS2 \s0_reg[18]  ( .CR(n87), .D(s0[6]), .CP(clk), .Q(s0[18]) );
  FDS2 \s0_reg[30]  ( .CR(n87), .D(s0[18]), .CP(clk), .Q(s0[30]) );
  FDS2 \s0_reg[11]  ( .CR(b0[11]), .D(n87), .CP(clk), .Q(s0[11]) );
  FDS2 \s0_reg[23]  ( .CR(n87), .D(s0[11]), .CP(clk), .Q(s0[23]) );
  FDS2 \s0_reg[17]  ( .CR(n87), .D(s0[5]), .CP(clk), .Q(s0[17]) );
  FDS2 \s0_reg[29]  ( .CR(n86), .D(s0[17]), .CP(clk), .Q(s0[29]) );
  FDS2 \s0_reg[10]  ( .CR(b0[10]), .D(n86), .CP(clk), .Q(s0[10]) );
  FDS2 \s0_reg[16]  ( .CR(n86), .D(s0[4]), .CP(clk), .Q(s0[16]) );
  FDS2 \s0_reg[28]  ( .CR(n86), .D(s0[16]), .CP(clk), .Q(s0[28]) );
  FDS2 \s0_reg[15]  ( .CR(n85), .D(s0[3]), .CP(clk), .Q(s0[15]) );
  FDS2 \s0_reg[27]  ( .CR(n85), .D(s0[15]), .CP(clk), .Q(s0[27]) );
  FDS2 \s0_reg[14]  ( .CR(n85), .D(s0[2]), .CP(clk), .Q(s0[14]) );
  FDS2 \s0_reg[26]  ( .CR(n85), .D(s0[14]), .CP(clk), .Q(s0[26]) );
  FDS2 \s0_reg[7]  ( .CR(b0[7]), .D(n88), .CP(clk), .Q(s0[7]) );
  FDS2 \s0_reg[6]  ( .CR(b0[6]), .D(n87), .CP(clk), .Q(s0[6]) );
  FDS2 \s0_reg[9]  ( .CR(b0[9]), .D(n86), .CP(clk), .Q(s0[9]) );
  FDS2 \s0_reg[8]  ( .CR(b0[8]), .D(n85), .CP(clk), .Q(s0[8]) );
  FDS2 \s2_reg[3]  ( .CR(b2[3]), .D(n74), .CP(clk), .Q(s2[3]) );
  FD1 \s2_reg[2]  ( .D(N238), .CP(clk), .Q(s2[2]) );
  FDS2 \s2_reg[1]  ( .CR(b2[1]), .D(n74), .CP(clk), .Q(s2[1]) );
  FD1 \s2_reg[0]  ( .D(N236), .CP(clk), .Q(s2[0]) );
  FD1 \s1_reg[2]  ( .D(N185), .CP(clk), .Q(s1[2]) );
  FD1 \s1_reg[1]  ( .D(N184), .CP(clk), .Q(s1[1]) );
  FD1 \s1_reg[0]  ( .D(N183), .CP(clk), .Q(s1[0]) );
  FDS2 \s2_reg[4]  ( .CR(b2[4]), .D(n81), .CP(clk), .Q(s2[4]) );
  FDS2 \s2_reg[5]  ( .CR(b2[5]), .D(n81), .CP(clk), .Q(s2[5]) );
  FDS2 \s2_reg[6]  ( .CR(b2[6]), .D(n80), .CP(clk), .Q(s2[6]) );
  FDS2 \s2_reg[7]  ( .CR(b2[7]), .D(n79), .CP(clk), .Q(s2[7]) );
  FDS2 \s1_reg[3]  ( .CR(b1[3]), .D(n84), .CP(clk), .Q(s1[3]) );
  FDS2 \s1_reg[7]  ( .CR(n84), .D(s1[3]), .CP(clk), .Q(s1[7]) );
  FDS2 \s1_reg[11]  ( .CR(n84), .D(s1[7]), .CP(clk), .Q(s1[11]) );
  FDS2 \s1_reg[15]  ( .CR(n84), .D(s1[11]), .CP(clk), .Q(s1[15]) );
  FDS2 \s1_reg[19]  ( .CR(n84), .D(s1[15]), .CP(clk), .Q(s1[19]) );
  FDS2 \s1_reg[4]  ( .CR(b1[4]), .D(n84), .CP(clk), .Q(s1[4]) );
  FDS2 \s1_reg[8]  ( .CR(n84), .D(s1[4]), .CP(clk), .Q(s1[8]) );
  FDS2 \s1_reg[12]  ( .CR(n83), .D(s1[8]), .CP(clk), .Q(s1[12]) );
  FDS2 \s1_reg[16]  ( .CR(n83), .D(s1[12]), .CP(clk), .Q(s1[16]) );
  FDS2 \s1_reg[20]  ( .CR(n83), .D(s1[16]), .CP(clk), .Q(s1[20]) );
  FDS2 \s1_reg[5]  ( .CR(b1[5]), .D(n83), .CP(clk), .Q(s1[5]) );
  FDS2 \s1_reg[9]  ( .CR(n83), .D(s1[5]), .CP(clk), .Q(s1[9]) );
  FDS2 \s1_reg[13]  ( .CR(n83), .D(s1[9]), .CP(clk), .Q(s1[13]) );
  FDS2 \s1_reg[17]  ( .CR(n83), .D(s1[13]), .CP(clk), .Q(s1[17]) );
  FDS2 \s1_reg[21]  ( .CR(n83), .D(s1[17]), .CP(clk), .Q(s1[21]) );
  FDS2 \s1_reg[6]  ( .CR(b1[6]), .D(n82), .CP(clk), .Q(s1[6]) );
  FDS2 \s1_reg[10]  ( .CR(n82), .D(s1[6]), .CP(clk), .Q(s1[10]) );
  FDS2 \s1_reg[14]  ( .CR(n82), .D(s1[10]), .CP(clk), .Q(s1[14]) );
  FDS2 \s1_reg[18]  ( .CR(n82), .D(s1[14]), .CP(clk), .Q(s1[18]) );
  FDS2 \s1_reg[22]  ( .CR(n82), .D(s1[18]), .CP(clk), .Q(s1[22]) );
  FDS2 \s2_reg[10]  ( .CR(b2[10]), .D(n81), .CP(clk), .Q(s2[10]) );
  FDS2 \s2_reg[16]  ( .CR(b2[16]), .D(n81), .CP(clk), .Q(s2[16]) );
  FDS2 \s2_reg[17]  ( .CR(b2[17]), .D(n80), .CP(clk), .Q(s2[17]) );
  FDS2 \s2_reg[29]  ( .CR(n80), .D(s2[12]), .CP(clk), .Q(s2[29]) );
  FDS2 \s2_reg[30]  ( .CR(n79), .D(s2[13]), .CP(clk), .Q(s2[30]) );
  FDS2 \s2_reg[8]  ( .CR(b2[8]), .D(n79), .CP(clk), .Q(s2[8]) );
  FDS2 \s2_reg[31]  ( .CR(n78), .D(s2[14]), .CP(clk), .Q(s2[31]) );
  FDS2 \s2_reg[9]  ( .CR(b2[9]), .D(n78), .CP(clk), .Q(s2[9]) );
  FDS2 \s2_reg[15]  ( .CR(b2[15]), .D(n78), .CP(clk), .Q(s2[15]) );
  FDS2 \s1_reg[23]  ( .CR(n84), .D(s1[19]), .CP(clk), .Q(s1[23]) );
  FDS2 \s1_reg[31]  ( .CR(n84), .D(s1[27]), .CP(clk), .Q(s1[31]) );
  FDS2 \s1_reg[24]  ( .CR(n83), .D(s1[20]), .CP(clk), .Q(s1[24]) );
  FDS2 \s1_reg[28]  ( .CR(n83), .D(s1[24]), .CP(clk), .Q(s1[28]) );
  FDS2 \s1_reg[29]  ( .CR(n82), .D(s1[25]), .CP(clk), .Q(s1[29]) );
  FDS2 \s1_reg[30]  ( .CR(n82), .D(s1[26]), .CP(clk), .Q(s1[30]) );
  FDS2 \s2_reg[21]  ( .CR(n81), .D(s2[4]), .CP(clk), .Q(s2[21]) );
  FDS2 \s2_reg[27]  ( .CR(n81), .D(s2[10]), .CP(clk), .Q(s2[27]) );
  FDS2 \s2_reg[22]  ( .CR(n81), .D(s2[5]), .CP(clk), .Q(s2[22]) );
  FDS2 \s2_reg[28]  ( .CR(n80), .D(s2[11]), .CP(clk), .Q(s2[28]) );
  FDS2 \s2_reg[23]  ( .CR(n80), .D(s2[6]), .CP(clk), .Q(s2[23]) );
  FDS2 \s2_reg[18]  ( .CR(b2[18]), .D(n80), .CP(clk), .Q(s2[18]) );
  FDS2 \s2_reg[24]  ( .CR(n79), .D(s2[7]), .CP(clk), .Q(s2[24]) );
  FDS2 \s2_reg[19]  ( .CR(b2[19]), .D(n79), .CP(clk), .Q(s2[19]) );
  FDS2 \s2_reg[25]  ( .CR(n79), .D(s2[8]), .CP(clk), .Q(s2[25]) );
  FDS2 \s2_reg[20]  ( .CR(b2[20]), .D(n78), .CP(clk), .Q(s2[20]) );
  FDS2 \s2_reg[26]  ( .CR(n78), .D(s2[9]), .CP(clk), .Q(s2[26]) );
  FDS2 \s2_reg[11]  ( .CR(b2[11]), .D(n80), .CP(clk), .Q(s2[11]) );
  FDS2 \s1_reg[25]  ( .CR(n83), .D(s1[21]), .CP(clk), .Q(s1[25]) );
  FDS2 \s2_reg[12]  ( .CR(b2[12]), .D(n80), .CP(clk), .Q(s2[12]) );
  FDS2 \s2_reg[13]  ( .CR(b2[13]), .D(n79), .CP(clk), .Q(s2[13]) );
  FDS2 \s2_reg[14]  ( .CR(b2[14]), .D(n78), .CP(clk), .Q(s2[14]) );
  FDS2 \s1_reg[27]  ( .CR(n84), .D(s1[23]), .CP(clk), .Q(s1[27]) );
  FDS2 \s1_reg[26]  ( .CR(n82), .D(s1[22]), .CP(clk), .Q(s1[26]) );
  FDS2 \b0_reg[7]  ( .CR(n88), .D(n73), .CP(clk), .Q(b0[7]) );
  FDS2 \b0_reg[12]  ( .CR(n88), .D(n72), .CP(clk), .Q(b0[12]) );
  FDS2 \b0_reg[6]  ( .CR(n87), .D(n71), .CP(clk), .Q(b0[6]) );
  FDS2 \b0_reg[11]  ( .CR(n87), .D(n70), .CP(clk), .Q(b0[11]) );
  FDS2 \b0_reg[5]  ( .CR(n87), .D(n69), .CP(clk), .Q(b0[5]) );
  FDS2 \b0_reg[10]  ( .CR(n86), .D(n68), .CP(clk), .Q(b0[10]) );
  FDS2 \b0_reg[4]  ( .CR(n86), .D(n67), .CP(clk), .Q(b0[4]) );
  FDS2 \b0_reg[9]  ( .CR(n86), .D(n66), .CP(clk), .Q(b0[9]) );
  FDS2 \b0_reg[3]  ( .CR(n86), .D(n65), .CP(clk), .Q(b0[3]) );
  FDS2 \b0_reg[8]  ( .CR(n85), .D(n64), .CP(clk), .Q(b0[8]) );
  FDS2 \b0_reg[2]  ( .CR(n85), .D(n63), .CP(clk), .Q(b0[2]) );
  FDS2 \b0_reg[0]  ( .CR(n85), .D(n62), .CP(clk), .Q(b0[0]) );
  FDS2 \b1_reg[4]  ( .CR(n84), .D(n43), .CP(clk), .Q(b1[4]) );
  FDS2 \b1_reg[5]  ( .CR(n83), .D(n60), .CP(clk), .Q(b1[5]) );
  FDS2 \b1_reg[6]  ( .CR(n82), .D(n59), .CP(clk), .Q(b1[6]) );
  FDS2 \b1_reg[3]  ( .CR(n82), .D(n42), .CP(clk), .Q(b1[3]) );
  FDS2 \b2_reg[10]  ( .CR(n81), .D(n58), .CP(clk), .Q(b2[10]) );
  FDS2 \b2_reg[16]  ( .CR(n81), .D(n57), .CP(clk), .Q(b2[16]) );
  FDS2 \b2_reg[5]  ( .CR(n81), .D(n37), .CP(clk), .Q(b2[5]) );
  FDS2 \b2_reg[11]  ( .CR(n81), .D(n56), .CP(clk), .Q(b2[11]) );
  FDS2 \b2_reg[17]  ( .CR(n80), .D(n55), .CP(clk), .Q(b2[17]) );
  FDS2 \b2_reg[6]  ( .CR(n80), .D(n22), .CP(clk), .Q(b2[6]) );
  FDS2 \b2_reg[12]  ( .CR(n80), .D(n54), .CP(clk), .Q(b2[12]) );
  FDS2 \b2_reg[18]  ( .CR(n80), .D(n53), .CP(clk), .Q(b2[18]) );
  FDS2 \b2_reg[7]  ( .CR(n79), .D(n52), .CP(clk), .Q(b2[7]) );
  FDS2 \b2_reg[13]  ( .CR(n79), .D(n51), .CP(clk), .Q(b2[13]) );
  FDS2 \b2_reg[19]  ( .CR(n79), .D(n50), .CP(clk), .Q(b2[19]) );
  FDS2 \b2_reg[8]  ( .CR(n79), .D(n49), .CP(clk), .Q(b2[8]) );
  FDS2 \b2_reg[14]  ( .CR(n79), .D(n48), .CP(clk), .Q(b2[14]) );
  FDS2L \Tout_reg[31]  ( .CR(1'b1), .D(N99), .LD(n78), .CP(clk), .Q(Tout[31])
         );
  FDS2 \b2_reg[20]  ( .CR(n78), .D(n47), .CP(clk), .Q(b2[20]) );
  FDS2 \b2_reg[9]  ( .CR(n78), .D(n46), .CP(clk), .Q(b2[9]) );
  FDS2 \b2_reg[15]  ( .CR(n78), .D(n45), .CP(clk), .Q(b2[15]) );
  FDS2L \Tout_reg[15]  ( .CR(1'b1), .D(N115), .LD(n78), .CP(clk), .Q(Tout[15])
         );
  FDS2L \Tout_reg[26]  ( .CR(1'b1), .D(N104), .LD(n78), .CP(clk), .Q(Tout[26])
         );
  FDS2L \Tout_reg[9]  ( .CR(1'b1), .D(N121), .LD(n77), .CP(clk), .Q(Tout[9])
         );
  FDS2L \Tout_reg[20]  ( .CR(1'b1), .D(N110), .LD(n77), .CP(clk), .Q(Tout[20])
         );
  FDS2L \Tout_reg[14]  ( .CR(1'b1), .D(N116), .LD(n77), .CP(clk), .Q(Tout[14])
         );
  FDS2L \Tout_reg[25]  ( .CR(1'b1), .D(N105), .LD(n77), .CP(clk), .Q(Tout[25])
         );
  FDS2L \Tout_reg[8]  ( .CR(1'b1), .D(N122), .LD(n77), .CP(clk), .Q(Tout[8])
         );
  FDS2L \Tout_reg[19]  ( .CR(1'b1), .D(N111), .LD(n77), .CP(clk), .Q(Tout[19])
         );
  FDS2L \Tout_reg[30]  ( .CR(1'b1), .D(N100), .LD(n77), .CP(clk), .Q(Tout[30])
         );
  FDS2L \Tout_reg[13]  ( .CR(1'b1), .D(N117), .LD(n77), .CP(clk), .Q(Tout[13])
         );
  FDS2L \Tout_reg[24]  ( .CR(1'b1), .D(N106), .LD(n77), .CP(clk), .Q(Tout[24])
         );
  FDS2L \Tout_reg[7]  ( .CR(1'b1), .D(N123), .LD(n77), .CP(clk), .Q(Tout[7])
         );
  FDS2L \Tout_reg[18]  ( .CR(1'b1), .D(N112), .LD(n77), .CP(clk), .Q(Tout[18])
         );
  FDS2L \Tout_reg[29]  ( .CR(1'b1), .D(N101), .LD(n77), .CP(clk), .Q(Tout[29])
         );
  FDS2 \b2_reg[4]  ( .CR(n76), .D(n21), .CP(clk), .Q(b2[4]) );
  FDS2 \b2_reg[1]  ( .CR(n76), .D(n15), .CP(clk), .Q(b2[1]) );
  FDS2L \Tout_reg[12]  ( .CR(1'b1), .D(N118), .LD(n76), .CP(clk), .Q(Tout[12])
         );
  FDS2L \Tout_reg[23]  ( .CR(1'b1), .D(N107), .LD(n76), .CP(clk), .Q(Tout[23])
         );
  FDS2L \Tout_reg[6]  ( .CR(1'b1), .D(N124), .LD(n76), .CP(clk), .Q(Tout[6])
         );
  FDS2L \Tout_reg[17]  ( .CR(1'b1), .D(N113), .LD(n76), .CP(clk), .Q(Tout[17])
         );
  FDS2L \Tout_reg[28]  ( .CR(1'b1), .D(N102), .LD(n76), .CP(clk), .Q(Tout[28])
         );
  FDS2 \b2_reg[3]  ( .CR(n76), .D(n14), .CP(clk), .Q(b2[3]) );
  FDS2L \Tout_reg[22]  ( .CR(1'b1), .D(N108), .LD(n76), .CP(clk), .Q(Tout[22])
         );
  FDS2L \Tout_reg[5]  ( .CR(1'b1), .D(N125), .LD(n76), .CP(clk), .Q(Tout[5])
         );
  FDS2L \Tout_reg[16]  ( .CR(1'b1), .D(N114), .LD(n74), .CP(clk), .Q(Tout[16])
         );
  FDS2L \Tout_reg[27]  ( .CR(1'b1), .D(N103), .LD(n74), .CP(clk), .Q(Tout[27])
         );
  FDS2L \Tout_reg[10]  ( .CR(1'b1), .D(N120), .LD(n74), .CP(clk), .Q(Tout[10])
         );
  FDS2L \Tout_reg[21]  ( .CR(1'b1), .D(N109), .LD(n74), .CP(clk), .Q(Tout[21])
         );
  FDS2L \Tout_reg[3]  ( .CR(1'b1), .D(N127), .LD(n74), .CP(clk), .Q(Tout[3])
         );
  FDS2L \Tout_reg[1]  ( .CR(1'b1), .D(N129), .LD(n74), .CP(clk), .Q(Tout[1])
         );
  FDS2L \Tout_reg[0]  ( .CR(1'b1), .D(N130), .LD(n74), .CP(clk), .Q(Tout[0])
         );
  IVP U10 ( .A(n91), .Z(n74) );
  IVP U16 ( .A(n91), .Z(n76) );
  IVP U17 ( .A(n91), .Z(n77) );
  IVP U23 ( .A(n91), .Z(n78) );
  IVP U24 ( .A(n90), .Z(n79) );
  IVP U39 ( .A(n90), .Z(n80) );
  IVP U40 ( .A(n90), .Z(n81) );
  IVP U41 ( .A(n90), .Z(n82) );
  IVP U43 ( .A(n90), .Z(n83) );
  IVP U44 ( .A(n89), .Z(n84) );
  IVP U45 ( .A(n89), .Z(n85) );
  IVP U46 ( .A(n89), .Z(n86) );
  IVP U47 ( .A(n89), .Z(n87) );
  EO U48 ( .A(s0[0]), .B(n117), .Z(N130) );
  EO U49 ( .A(s2[0]), .B(s1[0]), .Z(n117) );
  EO U50 ( .A(s0[1]), .B(n118), .Z(N129) );
  EO U51 ( .A(s2[1]), .B(s1[1]), .Z(n118) );
  EO U52 ( .A(s0[2]), .B(n119), .Z(N128) );
  EO U53 ( .A(s2[2]), .B(s1[2]), .Z(n119) );
  EO U54 ( .A(s0[27]), .B(n144), .Z(N103) );
  EO U55 ( .A(s2[27]), .B(s1[27]), .Z(n144) );
  EO U56 ( .A(s0[12]), .B(n129), .Z(N118) );
  EO U57 ( .A(s2[12]), .B(s1[12]), .Z(n129) );
  EO U58 ( .A(s0[13]), .B(n130), .Z(N117) );
  EO U59 ( .A(s2[13]), .B(s1[13]), .Z(n130) );
  EO U60 ( .A(s0[25]), .B(n142), .Z(N105) );
  EO U61 ( .A(s2[25]), .B(s1[25]), .Z(n142) );
  EO U62 ( .A(s0[14]), .B(n131), .Z(N116) );
  EO U63 ( .A(s2[14]), .B(s1[14]), .Z(n131) );
  EO U64 ( .A(s0[26]), .B(n143), .Z(N104) );
  EO U65 ( .A(s2[26]), .B(s1[26]), .Z(n143) );
  EO U66 ( .A(s0[3]), .B(n120), .Z(N127) );
  EO U67 ( .A(s2[3]), .B(s1[3]), .Z(n120) );
  EO U68 ( .A(s0[4]), .B(n121), .Z(N126) );
  EO U69 ( .A(s2[4]), .B(s1[4]), .Z(n121) );
  EO U70 ( .A(s0[21]), .B(n138), .Z(N109) );
  EO U71 ( .A(s2[21]), .B(s1[21]), .Z(n138) );
  EO U72 ( .A(s0[10]), .B(n127), .Z(N120) );
  EO U73 ( .A(s2[10]), .B(s1[10]), .Z(n127) );
  EO U74 ( .A(s0[16]), .B(n133), .Z(N114) );
  EO U75 ( .A(s2[16]), .B(s1[16]), .Z(n133) );
  EO U76 ( .A(s0[5]), .B(n122), .Z(N125) );
  EO U77 ( .A(s2[5]), .B(s1[5]), .Z(n122) );
  EO U78 ( .A(s0[22]), .B(n139), .Z(N108) );
  EO U79 ( .A(s2[22]), .B(s1[22]), .Z(n139) );
  EO U80 ( .A(s0[11]), .B(n128), .Z(N119) );
  EO U81 ( .A(s2[11]), .B(s1[11]), .Z(n128) );
  EO U82 ( .A(s0[28]), .B(n145), .Z(N102) );
  EO U83 ( .A(s2[28]), .B(s1[28]), .Z(n145) );
  EO U84 ( .A(s0[17]), .B(n134), .Z(N113) );
  EO U85 ( .A(s2[17]), .B(s1[17]), .Z(n134) );
  EO U86 ( .A(s0[6]), .B(n123), .Z(N124) );
  EO U87 ( .A(s2[6]), .B(s1[6]), .Z(n123) );
  EO U88 ( .A(s0[23]), .B(n140), .Z(N107) );
  EO U89 ( .A(s2[23]), .B(s1[23]), .Z(n140) );
  EO U90 ( .A(s0[29]), .B(n146), .Z(N101) );
  EO U91 ( .A(s2[29]), .B(s1[29]), .Z(n146) );
  EO U92 ( .A(s0[18]), .B(n135), .Z(N112) );
  EO U93 ( .A(s2[18]), .B(s1[18]), .Z(n135) );
  EO U94 ( .A(s0[7]), .B(n124), .Z(N123) );
  EO U95 ( .A(s2[7]), .B(s1[7]), .Z(n124) );
  EO U96 ( .A(s0[24]), .B(n141), .Z(N106) );
  EO U97 ( .A(s2[24]), .B(s1[24]), .Z(n141) );
  EO U98 ( .A(s0[30]), .B(n147), .Z(N100) );
  EO U99 ( .A(s2[30]), .B(s1[30]), .Z(n147) );
  EO U100 ( .A(s0[19]), .B(n136), .Z(N111) );
  EO U101 ( .A(s2[19]), .B(s1[19]), .Z(n136) );
  EO U102 ( .A(s0[8]), .B(n125), .Z(N122) );
  EO U103 ( .A(s2[8]), .B(s1[8]), .Z(n125) );
  EO U104 ( .A(s0[20]), .B(n137), .Z(N110) );
  EO U105 ( .A(s2[20]), .B(s1[20]), .Z(n137) );
  EO U106 ( .A(s0[9]), .B(n126), .Z(N121) );
  EO U107 ( .A(s2[9]), .B(s1[9]), .Z(n126) );
  EO U108 ( .A(s0[15]), .B(n132), .Z(N115) );
  EO U109 ( .A(s2[15]), .B(s1[15]), .Z(n132) );
  EO U110 ( .A(s0[31]), .B(n75), .Z(N99) );
  EO U111 ( .A(s2[31]), .B(s1[31]), .Z(n75) );
  EO U112 ( .A(s2[10]), .B(s2[13]), .Z(n8) );
  EO U113 ( .A(s2[11]), .B(s2[14]), .Z(n14) );
  EO U114 ( .A(s2[9]), .B(s2[12]), .Z(n15) );
  EO U115 ( .A(s2[15]), .B(s2[12]), .Z(n21) );
  EO U116 ( .A(s2[17]), .B(s2[14]), .Z(n22) );
  EO U117 ( .A(s2[16]), .B(s2[13]), .Z(n37) );
  EO U118 ( .A(s1[23]), .B(s1[25]), .Z(n38) );
  EO U119 ( .A(s1[25]), .B(s1[27]), .Z(n39) );
  EO U120 ( .A(s1[24]), .B(s1[26]), .Z(n41) );
  EO U121 ( .A(s1[28]), .B(s1[26]), .Z(n42) );
  EO U122 ( .A(s1[29]), .B(s1[27]), .Z(n43) );
  IVP U123 ( .A(reset), .Z(n92) );
  EO U124 ( .A(s2[8]), .B(s2[11]), .Z(n44) );
  EO U125 ( .A(s2[23]), .B(s2[26]), .Z(n45) );
  EO U126 ( .A(s2[17]), .B(s2[20]), .Z(n46) );
  EO U127 ( .A(s2[28]), .B(s2[31]), .Z(n47) );
  EO U128 ( .A(s2[22]), .B(s2[25]), .Z(n48) );
  EO U129 ( .A(s2[16]), .B(s2[19]), .Z(n49) );
  EO U130 ( .A(s2[27]), .B(s2[30]), .Z(n50) );
  EO U131 ( .A(s2[21]), .B(s2[24]), .Z(n51) );
  EO U132 ( .A(s2[15]), .B(s2[18]), .Z(n52) );
  EO U133 ( .A(s2[26]), .B(s2[29]), .Z(n53) );
  EO U134 ( .A(s2[20]), .B(s2[23]), .Z(n54) );
  EO U135 ( .A(s2[25]), .B(s2[28]), .Z(n55) );
  EO U136 ( .A(s2[19]), .B(s2[22]), .Z(n56) );
  EO U137 ( .A(s2[24]), .B(s2[27]), .Z(n57) );
  EO U138 ( .A(s2[18]), .B(s2[21]), .Z(n58) );
  EO U139 ( .A(s1[29]), .B(s1[31]), .Z(n59) );
  EO U140 ( .A(s1[28]), .B(s1[30]), .Z(n60) );
  EO U141 ( .A(s0[20]), .B(s0[7]), .Z(n61) );
  EO U142 ( .A(s0[19]), .B(s0[6]), .Z(n62) );
  EO U143 ( .A(s0[21]), .B(s0[8]), .Z(n63) );
  EO U144 ( .A(s0[14]), .B(s0[27]), .Z(n64) );
  EO U145 ( .A(s0[22]), .B(s0[9]), .Z(n65) );
  EO U146 ( .A(s0[15]), .B(s0[28]), .Z(n66) );
  EO U147 ( .A(s0[10]), .B(s0[23]), .Z(n67) );
  EO U148 ( .A(s0[16]), .B(s0[29]), .Z(n68) );
  EO U149 ( .A(s0[11]), .B(s0[24]), .Z(n69) );
  EO U150 ( .A(s0[17]), .B(s0[30]), .Z(n70) );
  EO U151 ( .A(s0[12]), .B(s0[25]), .Z(n71) );
  EO U152 ( .A(s0[18]), .B(s0[31]), .Z(n72) );
  EO U153 ( .A(s0[13]), .B(s0[26]), .Z(n73) );
  IV U154 ( .A(n89), .Z(n88) );
  IVA U155 ( .A(n92), .Z(n89) );
  IVA U156 ( .A(n92), .Z(n90) );
  IVA U157 ( .A(n92), .Z(n91) );
endmodule


module Taus_1 ( clk, reset, Tout );
  output [31:0] Tout;
  input clk, reset;
  wire   N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N145, N183,
         N184, N185, N236, N238, n8, n14, n15, n21, n22, n37, n38, n39, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n124, n125, n126, n127, n128,
         n129, n130, n131;
  wire   [31:0] s0;
  wire   [31:0] b0;
  wire   [31:0] s1;
  wire   [31:0] b1;
  wire   [31:0] s2;
  wire   [31:0] b2;

  OR2 U182 ( .A(b2[2]), .B(reset), .Z(N238) );
  OR2 U183 ( .A(b2[0]), .B(reset), .Z(N236) );
  OR2 U184 ( .A(b1[2]), .B(reset), .Z(N185) );
  OR2 U185 ( .A(b1[1]), .B(reset), .Z(N184) );
  OR2 U186 ( .A(b1[0]), .B(reset), .Z(N183) );
  OR2 U187 ( .A(b0[1]), .B(reset), .Z(N145) );
  FDS2 \b0_reg[1]  ( .CR(n85), .D(n61), .CP(clk), .Q(b0[1]) );
  FDS2 \b1_reg[1]  ( .CR(n82), .D(n41), .CP(clk), .Q(b1[1]) );
  FDS2 \b1_reg[2]  ( .CR(n82), .D(n39), .CP(clk), .Q(b1[2]) );
  FDS2 \b1_reg[0]  ( .CR(n81), .D(n38), .CP(clk), .Q(b1[0]) );
  FDS2 \b2_reg[0]  ( .CR(n76), .D(n44), .CP(clk), .Q(b2[0]) );
  FDS2 \b2_reg[2]  ( .CR(n74), .D(n8), .CP(clk), .Q(b2[2]) );
  FDS2L \Tout_reg[18]  ( .CR(1'b1), .D(N112), .LD(n77), .CP(clk), .Q(Tout[18])
         );
  FDS2L \Tout_reg[28]  ( .CR(1'b1), .D(N102), .LD(n76), .CP(clk), .Q(Tout[28])
         );
  FDS2L \Tout_reg[27]  ( .CR(1'b1), .D(N103), .LD(n74), .CP(clk), .Q(Tout[27])
         );
  FDS2 \s0_reg[0]  ( .CR(b0[0]), .D(n84), .CP(clk), .Q(s0[0]) );
  FD1 \s0_reg[1]  ( .D(N145), .CP(clk), .Q(s0[1]) );
  FDS2 \s0_reg[5]  ( .CR(b0[5]), .D(n87), .CP(clk), .Q(s0[5]) );
  FDS2 \s0_reg[22]  ( .CR(n86), .D(s0[10]), .CP(clk), .Q(s0[22]) );
  FDS2 \s0_reg[4]  ( .CR(b0[4]), .D(n86), .CP(clk), .Q(s0[4]) );
  FDS2 \s0_reg[21]  ( .CR(n86), .D(s0[9]), .CP(clk), .Q(s0[21]) );
  FDS2 \s0_reg[3]  ( .CR(b0[3]), .D(n85), .CP(clk), .Q(s0[3]) );
  FDS2 \s0_reg[20]  ( .CR(n85), .D(s0[8]), .CP(clk), .Q(s0[20]) );
  FDS2 \s0_reg[2]  ( .CR(b0[2]), .D(n85), .CP(clk), .Q(s0[2]) );
  FDS2 \s0_reg[13]  ( .CR(n88), .D(s0[1]), .CP(clk), .Q(s0[13]) );
  FDS2 \s0_reg[25]  ( .CR(n88), .D(s0[13]), .CP(clk), .Q(s0[25]) );
  FDS2 \s0_reg[19]  ( .CR(n88), .D(s0[7]), .CP(clk), .Q(s0[19]) );
  FDS2 \s0_reg[31]  ( .CR(n88), .D(s0[19]), .CP(clk), .Q(s0[31]) );
  FDS2 \s0_reg[12]  ( .CR(b0[12]), .D(n87), .CP(clk), .Q(s0[12]) );
  FDS2 \s0_reg[24]  ( .CR(n87), .D(s0[12]), .CP(clk), .Q(s0[24]) );
  FDS2 \s0_reg[18]  ( .CR(n87), .D(s0[6]), .CP(clk), .Q(s0[18]) );
  FDS2 \s0_reg[30]  ( .CR(n87), .D(s0[18]), .CP(clk), .Q(s0[30]) );
  FDS2 \s0_reg[11]  ( .CR(b0[11]), .D(n87), .CP(clk), .Q(s0[11]) );
  FDS2 \s0_reg[23]  ( .CR(n87), .D(s0[11]), .CP(clk), .Q(s0[23]) );
  FDS2 \s0_reg[17]  ( .CR(n87), .D(s0[5]), .CP(clk), .Q(s0[17]) );
  FDS2 \s0_reg[29]  ( .CR(n86), .D(s0[17]), .CP(clk), .Q(s0[29]) );
  FDS2 \s0_reg[10]  ( .CR(b0[10]), .D(n86), .CP(clk), .Q(s0[10]) );
  FDS2 \s0_reg[16]  ( .CR(n86), .D(s0[4]), .CP(clk), .Q(s0[16]) );
  FDS2 \s0_reg[28]  ( .CR(n86), .D(s0[16]), .CP(clk), .Q(s0[28]) );
  FDS2 \s0_reg[15]  ( .CR(n85), .D(s0[3]), .CP(clk), .Q(s0[15]) );
  FDS2 \s0_reg[27]  ( .CR(n85), .D(s0[15]), .CP(clk), .Q(s0[27]) );
  FDS2 \s0_reg[14]  ( .CR(n85), .D(s0[2]), .CP(clk), .Q(s0[14]) );
  FDS2 \s0_reg[26]  ( .CR(n85), .D(s0[14]), .CP(clk), .Q(s0[26]) );
  FDS2 \s0_reg[7]  ( .CR(b0[7]), .D(n88), .CP(clk), .Q(s0[7]) );
  FDS2 \s0_reg[6]  ( .CR(b0[6]), .D(n87), .CP(clk), .Q(s0[6]) );
  FDS2 \s0_reg[9]  ( .CR(b0[9]), .D(n86), .CP(clk), .Q(s0[9]) );
  FDS2 \s0_reg[8]  ( .CR(b0[8]), .D(n85), .CP(clk), .Q(s0[8]) );
  FDS2 \s2_reg[3]  ( .CR(b2[3]), .D(n74), .CP(clk), .Q(s2[3]) );
  FD1 \s2_reg[2]  ( .D(N238), .CP(clk), .Q(s2[2]) );
  FDS2 \s2_reg[1]  ( .CR(b2[1]), .D(n74), .CP(clk), .Q(s2[1]) );
  FD1 \s2_reg[0]  ( .D(N236), .CP(clk), .Q(s2[0]) );
  FD1 \s1_reg[2]  ( .D(N185), .CP(clk), .Q(s1[2]) );
  FD1 \s1_reg[1]  ( .D(N184), .CP(clk), .Q(s1[1]) );
  FD1 \s1_reg[0]  ( .D(N183), .CP(clk), .Q(s1[0]) );
  FDS2 \s2_reg[4]  ( .CR(b2[4]), .D(n81), .CP(clk), .Q(s2[4]) );
  FDS2 \s2_reg[5]  ( .CR(b2[5]), .D(n81), .CP(clk), .Q(s2[5]) );
  FDS2 \s2_reg[6]  ( .CR(b2[6]), .D(n80), .CP(clk), .Q(s2[6]) );
  FDS2 \s2_reg[7]  ( .CR(b2[7]), .D(n79), .CP(clk), .Q(s2[7]) );
  FDS2 \s1_reg[3]  ( .CR(b1[3]), .D(n84), .CP(clk), .Q(s1[3]) );
  FDS2 \s1_reg[7]  ( .CR(n84), .D(s1[3]), .CP(clk), .Q(s1[7]) );
  FDS2 \s1_reg[11]  ( .CR(n84), .D(s1[7]), .CP(clk), .Q(s1[11]) );
  FDS2 \s1_reg[15]  ( .CR(n84), .D(s1[11]), .CP(clk), .Q(s1[15]) );
  FDS2 \s1_reg[19]  ( .CR(n84), .D(s1[15]), .CP(clk), .Q(s1[19]) );
  FDS2 \s1_reg[4]  ( .CR(b1[4]), .D(n84), .CP(clk), .Q(s1[4]) );
  FDS2 \s1_reg[8]  ( .CR(n84), .D(s1[4]), .CP(clk), .Q(s1[8]) );
  FDS2 \s1_reg[12]  ( .CR(n83), .D(s1[8]), .CP(clk), .Q(s1[12]) );
  FDS2 \s1_reg[16]  ( .CR(n83), .D(s1[12]), .CP(clk), .Q(s1[16]) );
  FDS2 \s1_reg[20]  ( .CR(n83), .D(s1[16]), .CP(clk), .Q(s1[20]) );
  FDS2 \s1_reg[5]  ( .CR(b1[5]), .D(n83), .CP(clk), .Q(s1[5]) );
  FDS2 \s1_reg[9]  ( .CR(n83), .D(s1[5]), .CP(clk), .Q(s1[9]) );
  FDS2 \s1_reg[13]  ( .CR(n83), .D(s1[9]), .CP(clk), .Q(s1[13]) );
  FDS2 \s1_reg[17]  ( .CR(n83), .D(s1[13]), .CP(clk), .Q(s1[17]) );
  FDS2 \s1_reg[21]  ( .CR(n83), .D(s1[17]), .CP(clk), .Q(s1[21]) );
  FDS2 \s1_reg[6]  ( .CR(b1[6]), .D(n82), .CP(clk), .Q(s1[6]) );
  FDS2 \s1_reg[10]  ( .CR(n82), .D(s1[6]), .CP(clk), .Q(s1[10]) );
  FDS2 \s1_reg[14]  ( .CR(n82), .D(s1[10]), .CP(clk), .Q(s1[14]) );
  FDS2 \s1_reg[18]  ( .CR(n82), .D(s1[14]), .CP(clk), .Q(s1[18]) );
  FDS2 \s1_reg[22]  ( .CR(n82), .D(s1[18]), .CP(clk), .Q(s1[22]) );
  FDS2 \s2_reg[10]  ( .CR(b2[10]), .D(n81), .CP(clk), .Q(s2[10]) );
  FDS2 \s2_reg[16]  ( .CR(b2[16]), .D(n81), .CP(clk), .Q(s2[16]) );
  FDS2 \s2_reg[17]  ( .CR(b2[17]), .D(n80), .CP(clk), .Q(s2[17]) );
  FDS2 \s2_reg[29]  ( .CR(n80), .D(s2[12]), .CP(clk), .Q(s2[29]) );
  FDS2 \s2_reg[30]  ( .CR(n79), .D(s2[13]), .CP(clk), .Q(s2[30]) );
  FDS2 \s2_reg[8]  ( .CR(b2[8]), .D(n79), .CP(clk), .Q(s2[8]) );
  FDS2 \s2_reg[31]  ( .CR(n78), .D(s2[14]), .CP(clk), .Q(s2[31]) );
  FDS2 \s2_reg[9]  ( .CR(b2[9]), .D(n78), .CP(clk), .Q(s2[9]) );
  FDS2 \s2_reg[15]  ( .CR(b2[15]), .D(n78), .CP(clk), .Q(s2[15]) );
  FDS2 \s1_reg[23]  ( .CR(n84), .D(s1[19]), .CP(clk), .Q(s1[23]) );
  FDS2 \s1_reg[31]  ( .CR(n84), .D(s1[27]), .CP(clk), .Q(s1[31]) );
  FDS2 \s1_reg[24]  ( .CR(n83), .D(s1[20]), .CP(clk), .Q(s1[24]) );
  FDS2 \s1_reg[28]  ( .CR(n83), .D(s1[24]), .CP(clk), .Q(s1[28]) );
  FDS2 \s1_reg[29]  ( .CR(n82), .D(s1[25]), .CP(clk), .Q(s1[29]) );
  FDS2 \s1_reg[30]  ( .CR(n82), .D(s1[26]), .CP(clk), .Q(s1[30]) );
  FDS2 \s2_reg[21]  ( .CR(n81), .D(s2[4]), .CP(clk), .Q(s2[21]) );
  FDS2 \s2_reg[27]  ( .CR(n81), .D(s2[10]), .CP(clk), .Q(s2[27]) );
  FDS2 \s2_reg[22]  ( .CR(n81), .D(s2[5]), .CP(clk), .Q(s2[22]) );
  FDS2 \s2_reg[28]  ( .CR(n80), .D(s2[11]), .CP(clk), .Q(s2[28]) );
  FDS2 \s2_reg[23]  ( .CR(n80), .D(s2[6]), .CP(clk), .Q(s2[23]) );
  FDS2 \s2_reg[18]  ( .CR(b2[18]), .D(n80), .CP(clk), .Q(s2[18]) );
  FDS2 \s2_reg[24]  ( .CR(n79), .D(s2[7]), .CP(clk), .Q(s2[24]) );
  FDS2 \s2_reg[19]  ( .CR(b2[19]), .D(n79), .CP(clk), .Q(s2[19]) );
  FDS2 \s2_reg[25]  ( .CR(n79), .D(s2[8]), .CP(clk), .Q(s2[25]) );
  FDS2 \s2_reg[20]  ( .CR(b2[20]), .D(n78), .CP(clk), .Q(s2[20]) );
  FDS2 \s2_reg[26]  ( .CR(n78), .D(s2[9]), .CP(clk), .Q(s2[26]) );
  FDS2 \s2_reg[11]  ( .CR(b2[11]), .D(n80), .CP(clk), .Q(s2[11]) );
  FDS2 \s1_reg[25]  ( .CR(n83), .D(s1[21]), .CP(clk), .Q(s1[25]) );
  FDS2 \s2_reg[12]  ( .CR(b2[12]), .D(n80), .CP(clk), .Q(s2[12]) );
  FDS2 \s2_reg[13]  ( .CR(b2[13]), .D(n79), .CP(clk), .Q(s2[13]) );
  FDS2 \s2_reg[14]  ( .CR(b2[14]), .D(n78), .CP(clk), .Q(s2[14]) );
  FDS2 \s1_reg[27]  ( .CR(n84), .D(s1[23]), .CP(clk), .Q(s1[27]) );
  FDS2 \s1_reg[26]  ( .CR(n82), .D(s1[22]), .CP(clk), .Q(s1[26]) );
  FDS2 \b0_reg[7]  ( .CR(n88), .D(n73), .CP(clk), .Q(b0[7]) );
  FDS2 \b0_reg[12]  ( .CR(n88), .D(n72), .CP(clk), .Q(b0[12]) );
  FDS2 \b0_reg[6]  ( .CR(n87), .D(n71), .CP(clk), .Q(b0[6]) );
  FDS2 \b0_reg[11]  ( .CR(n87), .D(n70), .CP(clk), .Q(b0[11]) );
  FDS2 \b0_reg[5]  ( .CR(n87), .D(n69), .CP(clk), .Q(b0[5]) );
  FDS2 \b0_reg[10]  ( .CR(n86), .D(n68), .CP(clk), .Q(b0[10]) );
  FDS2 \b0_reg[4]  ( .CR(n86), .D(n67), .CP(clk), .Q(b0[4]) );
  FDS2 \b0_reg[9]  ( .CR(n86), .D(n66), .CP(clk), .Q(b0[9]) );
  FDS2 \b0_reg[3]  ( .CR(n86), .D(n65), .CP(clk), .Q(b0[3]) );
  FDS2 \b0_reg[8]  ( .CR(n85), .D(n64), .CP(clk), .Q(b0[8]) );
  FDS2 \b0_reg[2]  ( .CR(n85), .D(n63), .CP(clk), .Q(b0[2]) );
  FDS2 \b0_reg[0]  ( .CR(n85), .D(n62), .CP(clk), .Q(b0[0]) );
  FDS2 \b1_reg[4]  ( .CR(n84), .D(n43), .CP(clk), .Q(b1[4]) );
  FDS2 \b1_reg[5]  ( .CR(n83), .D(n60), .CP(clk), .Q(b1[5]) );
  FDS2 \b1_reg[6]  ( .CR(n82), .D(n59), .CP(clk), .Q(b1[6]) );
  FDS2 \b1_reg[3]  ( .CR(n82), .D(n42), .CP(clk), .Q(b1[3]) );
  FDS2 \b2_reg[10]  ( .CR(n81), .D(n58), .CP(clk), .Q(b2[10]) );
  FDS2 \b2_reg[16]  ( .CR(n81), .D(n57), .CP(clk), .Q(b2[16]) );
  FDS2 \b2_reg[5]  ( .CR(n81), .D(n37), .CP(clk), .Q(b2[5]) );
  FDS2 \b2_reg[11]  ( .CR(n81), .D(n56), .CP(clk), .Q(b2[11]) );
  FDS2 \b2_reg[17]  ( .CR(n80), .D(n55), .CP(clk), .Q(b2[17]) );
  FDS2 \b2_reg[6]  ( .CR(n80), .D(n22), .CP(clk), .Q(b2[6]) );
  FDS2 \b2_reg[12]  ( .CR(n80), .D(n54), .CP(clk), .Q(b2[12]) );
  FDS2 \b2_reg[18]  ( .CR(n80), .D(n53), .CP(clk), .Q(b2[18]) );
  FDS2 \b2_reg[7]  ( .CR(n79), .D(n52), .CP(clk), .Q(b2[7]) );
  FDS2 \b2_reg[13]  ( .CR(n79), .D(n51), .CP(clk), .Q(b2[13]) );
  FDS2 \b2_reg[19]  ( .CR(n79), .D(n50), .CP(clk), .Q(b2[19]) );
  FDS2 \b2_reg[8]  ( .CR(n79), .D(n49), .CP(clk), .Q(b2[8]) );
  FDS2 \b2_reg[14]  ( .CR(n79), .D(n48), .CP(clk), .Q(b2[14]) );
  FDS2L \Tout_reg[31]  ( .CR(1'b1), .D(N99), .LD(n78), .CP(clk), .Q(Tout[31])
         );
  FDS2 \b2_reg[20]  ( .CR(n78), .D(n47), .CP(clk), .Q(b2[20]) );
  FDS2 \b2_reg[9]  ( .CR(n78), .D(n46), .CP(clk), .Q(b2[9]) );
  FDS2 \b2_reg[15]  ( .CR(n78), .D(n45), .CP(clk), .Q(b2[15]) );
  FDS2L \Tout_reg[15]  ( .CR(1'b1), .D(N115), .LD(n78), .CP(clk), .Q(Tout[15])
         );
  FDS2L \Tout_reg[26]  ( .CR(1'b1), .D(N104), .LD(n78), .CP(clk), .Q(Tout[26])
         );
  FDS2L \Tout_reg[9]  ( .CR(1'b1), .D(N121), .LD(n77), .CP(clk), .Q(Tout[9])
         );
  FDS2L \Tout_reg[20]  ( .CR(1'b1), .D(N110), .LD(n77), .CP(clk), .Q(Tout[20])
         );
  FDS2L \Tout_reg[14]  ( .CR(1'b1), .D(N116), .LD(n77), .CP(clk), .Q(Tout[14])
         );
  FDS2L \Tout_reg[25]  ( .CR(1'b1), .D(N105), .LD(n77), .CP(clk), .Q(Tout[25])
         );
  FDS2L \Tout_reg[8]  ( .CR(1'b1), .D(N122), .LD(n77), .CP(clk), .Q(Tout[8])
         );
  FDS2L \Tout_reg[19]  ( .CR(1'b1), .D(N111), .LD(n77), .CP(clk), .Q(Tout[19])
         );
  FDS2L \Tout_reg[30]  ( .CR(1'b1), .D(N100), .LD(n77), .CP(clk), .Q(Tout[30])
         );
  FDS2L \Tout_reg[13]  ( .CR(1'b1), .D(N117), .LD(n77), .CP(clk), .Q(Tout[13])
         );
  FDS2L \Tout_reg[24]  ( .CR(1'b1), .D(N106), .LD(n77), .CP(clk), .Q(Tout[24])
         );
  FDS2L \Tout_reg[7]  ( .CR(1'b1), .D(N123), .LD(n77), .CP(clk), .Q(Tout[7])
         );
  FDS2L \Tout_reg[29]  ( .CR(1'b1), .D(N101), .LD(n77), .CP(clk), .Q(Tout[29])
         );
  FDS2 \b2_reg[4]  ( .CR(n76), .D(n21), .CP(clk), .Q(b2[4]) );
  FDS2 \b2_reg[1]  ( .CR(n76), .D(n15), .CP(clk), .Q(b2[1]) );
  FDS2L \Tout_reg[12]  ( .CR(1'b1), .D(N118), .LD(n76), .CP(clk), .Q(Tout[12])
         );
  FDS2L \Tout_reg[23]  ( .CR(1'b1), .D(N107), .LD(n76), .CP(clk), .Q(Tout[23])
         );
  FDS2L \Tout_reg[6]  ( .CR(1'b1), .D(N124), .LD(n76), .CP(clk), .Q(Tout[6])
         );
  FDS2L \Tout_reg[17]  ( .CR(1'b1), .D(N113), .LD(n76), .CP(clk), .Q(Tout[17])
         );
  FDS2 \b2_reg[3]  ( .CR(n76), .D(n14), .CP(clk), .Q(b2[3]) );
  FDS2L \Tout_reg[11]  ( .CR(1'b1), .D(N119), .LD(n76), .CP(clk), .Q(Tout[11])
         );
  FDS2L \Tout_reg[22]  ( .CR(1'b1), .D(N108), .LD(n76), .CP(clk), .Q(Tout[22])
         );
  FDS2L \Tout_reg[5]  ( .CR(1'b1), .D(N125), .LD(n76), .CP(clk), .Q(Tout[5])
         );
  FDS2L \Tout_reg[16]  ( .CR(1'b1), .D(N114), .LD(n74), .CP(clk), .Q(Tout[16])
         );
  FDS2L \Tout_reg[10]  ( .CR(1'b1), .D(N120), .LD(n74), .CP(clk), .Q(Tout[10])
         );
  FDS2L \Tout_reg[21]  ( .CR(1'b1), .D(N109), .LD(n74), .CP(clk), .Q(Tout[21])
         );
  FDS2L \Tout_reg[4]  ( .CR(1'b1), .D(N126), .LD(n74), .CP(clk), .Q(Tout[4])
         );
  FDS2L \Tout_reg[3]  ( .CR(1'b1), .D(N127), .LD(n74), .CP(clk), .Q(Tout[3])
         );
  FDS2L \Tout_reg[2]  ( .CR(1'b1), .D(N128), .LD(n74), .CP(clk), .Q(Tout[2])
         );
  FDS2L \Tout_reg[1]  ( .CR(1'b1), .D(N129), .LD(n74), .CP(clk), .Q(Tout[1])
         );
  FDS2L \Tout_reg[0]  ( .CR(1'b1), .D(N130), .LD(n74), .CP(clk), .Q(Tout[0])
         );
  IVP U10 ( .A(n91), .Z(n74) );
  IVP U16 ( .A(n91), .Z(n76) );
  IVP U17 ( .A(n91), .Z(n77) );
  IVP U23 ( .A(n91), .Z(n78) );
  IVP U24 ( .A(n90), .Z(n79) );
  IVP U39 ( .A(n90), .Z(n80) );
  IVP U40 ( .A(n90), .Z(n81) );
  IVP U41 ( .A(n90), .Z(n82) );
  IVP U43 ( .A(n90), .Z(n83) );
  IVP U44 ( .A(n89), .Z(n84) );
  IVP U45 ( .A(n89), .Z(n85) );
  IVP U46 ( .A(n89), .Z(n86) );
  IVP U47 ( .A(n89), .Z(n87) );
  EO U48 ( .A(s0[0]), .B(n130), .Z(N130) );
  EO U49 ( .A(s2[0]), .B(s1[0]), .Z(n130) );
  EO U50 ( .A(s0[1]), .B(n129), .Z(N129) );
  EO U51 ( .A(s2[1]), .B(s1[1]), .Z(n129) );
  EO U52 ( .A(s0[2]), .B(n128), .Z(N128) );
  EO U53 ( .A(s2[2]), .B(s1[2]), .Z(n128) );
  EO U54 ( .A(s0[27]), .B(n96), .Z(N103) );
  EO U55 ( .A(s2[27]), .B(s1[27]), .Z(n96) );
  EO U56 ( .A(s0[12]), .B(n111), .Z(N118) );
  EO U57 ( .A(s2[12]), .B(s1[12]), .Z(n111) );
  EO U58 ( .A(s0[13]), .B(n110), .Z(N117) );
  EO U59 ( .A(s2[13]), .B(s1[13]), .Z(n110) );
  EO U60 ( .A(s0[25]), .B(n98), .Z(N105) );
  EO U61 ( .A(s2[25]), .B(s1[25]), .Z(n98) );
  EO U62 ( .A(s0[14]), .B(n109), .Z(N116) );
  EO U63 ( .A(s2[14]), .B(s1[14]), .Z(n109) );
  EO U64 ( .A(s0[26]), .B(n97), .Z(N104) );
  EO U65 ( .A(s2[26]), .B(s1[26]), .Z(n97) );
  EO U66 ( .A(s0[3]), .B(n127), .Z(N127) );
  EO U67 ( .A(s2[3]), .B(s1[3]), .Z(n127) );
  EO U68 ( .A(s0[4]), .B(n126), .Z(N126) );
  EO U69 ( .A(s2[4]), .B(s1[4]), .Z(n126) );
  EO U70 ( .A(s0[21]), .B(n102), .Z(N109) );
  EO U71 ( .A(s2[21]), .B(s1[21]), .Z(n102) );
  EO U72 ( .A(s0[10]), .B(n113), .Z(N120) );
  EO U73 ( .A(s2[10]), .B(s1[10]), .Z(n113) );
  EO U74 ( .A(s0[16]), .B(n107), .Z(N114) );
  EO U75 ( .A(s2[16]), .B(s1[16]), .Z(n107) );
  EO U76 ( .A(s0[5]), .B(n125), .Z(N125) );
  EO U77 ( .A(s2[5]), .B(s1[5]), .Z(n125) );
  EO U78 ( .A(s0[22]), .B(n101), .Z(N108) );
  EO U79 ( .A(s2[22]), .B(s1[22]), .Z(n101) );
  EO U80 ( .A(s0[11]), .B(n112), .Z(N119) );
  EO U81 ( .A(s2[11]), .B(s1[11]), .Z(n112) );
  EO U82 ( .A(s0[28]), .B(n95), .Z(N102) );
  EO U83 ( .A(s2[28]), .B(s1[28]), .Z(n95) );
  EO U84 ( .A(s0[17]), .B(n106), .Z(N113) );
  EO U85 ( .A(s2[17]), .B(s1[17]), .Z(n106) );
  EO U86 ( .A(s0[6]), .B(n124), .Z(N124) );
  EO U87 ( .A(s2[6]), .B(s1[6]), .Z(n124) );
  EO U88 ( .A(s0[23]), .B(n100), .Z(N107) );
  EO U89 ( .A(s2[23]), .B(s1[23]), .Z(n100) );
  EO U90 ( .A(s0[29]), .B(n94), .Z(N101) );
  EO U91 ( .A(s2[29]), .B(s1[29]), .Z(n94) );
  EO U92 ( .A(s0[18]), .B(n105), .Z(N112) );
  EO U93 ( .A(s2[18]), .B(s1[18]), .Z(n105) );
  EO U94 ( .A(s0[7]), .B(n116), .Z(N123) );
  EO U95 ( .A(s2[7]), .B(s1[7]), .Z(n116) );
  EO U96 ( .A(s0[24]), .B(n99), .Z(N106) );
  EO U97 ( .A(s2[24]), .B(s1[24]), .Z(n99) );
  EO U98 ( .A(s0[30]), .B(n93), .Z(N100) );
  EO U99 ( .A(s2[30]), .B(s1[30]), .Z(n93) );
  EO U100 ( .A(s0[19]), .B(n104), .Z(N111) );
  EO U101 ( .A(s2[19]), .B(s1[19]), .Z(n104) );
  EO U102 ( .A(s0[8]), .B(n115), .Z(N122) );
  EO U103 ( .A(s2[8]), .B(s1[8]), .Z(n115) );
  EO U104 ( .A(s0[20]), .B(n103), .Z(N110) );
  EO U105 ( .A(s2[20]), .B(s1[20]), .Z(n103) );
  EO U106 ( .A(s0[9]), .B(n114), .Z(N121) );
  EO U107 ( .A(s2[9]), .B(s1[9]), .Z(n114) );
  EO U108 ( .A(s0[15]), .B(n108), .Z(N115) );
  EO U109 ( .A(s2[15]), .B(s1[15]), .Z(n108) );
  EO U110 ( .A(s0[31]), .B(n131), .Z(N99) );
  EO U111 ( .A(s2[31]), .B(s1[31]), .Z(n131) );
  EO U112 ( .A(s2[10]), .B(s2[13]), .Z(n8) );
  EO U113 ( .A(s2[11]), .B(s2[14]), .Z(n14) );
  EO U114 ( .A(s2[9]), .B(s2[12]), .Z(n15) );
  EO U115 ( .A(s2[15]), .B(s2[12]), .Z(n21) );
  EO U116 ( .A(s2[17]), .B(s2[14]), .Z(n22) );
  EO U117 ( .A(s2[16]), .B(s2[13]), .Z(n37) );
  EO U118 ( .A(s1[23]), .B(s1[25]), .Z(n38) );
  EO U119 ( .A(s1[25]), .B(s1[27]), .Z(n39) );
  EO U120 ( .A(s1[24]), .B(s1[26]), .Z(n41) );
  EO U121 ( .A(s1[28]), .B(s1[26]), .Z(n42) );
  EO U122 ( .A(s1[29]), .B(s1[27]), .Z(n43) );
  IVP U123 ( .A(reset), .Z(n92) );
  EO U124 ( .A(s2[8]), .B(s2[11]), .Z(n44) );
  EO U125 ( .A(s2[23]), .B(s2[26]), .Z(n45) );
  EO U126 ( .A(s2[17]), .B(s2[20]), .Z(n46) );
  EO U127 ( .A(s2[28]), .B(s2[31]), .Z(n47) );
  EO U128 ( .A(s2[22]), .B(s2[25]), .Z(n48) );
  EO U129 ( .A(s2[16]), .B(s2[19]), .Z(n49) );
  EO U130 ( .A(s2[27]), .B(s2[30]), .Z(n50) );
  EO U131 ( .A(s2[21]), .B(s2[24]), .Z(n51) );
  EO U132 ( .A(s2[15]), .B(s2[18]), .Z(n52) );
  EO U133 ( .A(s2[26]), .B(s2[29]), .Z(n53) );
  EO U134 ( .A(s2[20]), .B(s2[23]), .Z(n54) );
  EO U135 ( .A(s2[25]), .B(s2[28]), .Z(n55) );
  EO U136 ( .A(s2[19]), .B(s2[22]), .Z(n56) );
  EO U137 ( .A(s2[24]), .B(s2[27]), .Z(n57) );
  EO U138 ( .A(s2[18]), .B(s2[21]), .Z(n58) );
  EO U139 ( .A(s1[29]), .B(s1[31]), .Z(n59) );
  EO U140 ( .A(s1[28]), .B(s1[30]), .Z(n60) );
  EO U141 ( .A(s0[20]), .B(s0[7]), .Z(n61) );
  EO U142 ( .A(s0[19]), .B(s0[6]), .Z(n62) );
  EO U143 ( .A(s0[21]), .B(s0[8]), .Z(n63) );
  EO U144 ( .A(s0[14]), .B(s0[27]), .Z(n64) );
  EO U145 ( .A(s0[22]), .B(s0[9]), .Z(n65) );
  EO U146 ( .A(s0[15]), .B(s0[28]), .Z(n66) );
  EO U147 ( .A(s0[10]), .B(s0[23]), .Z(n67) );
  EO U148 ( .A(s0[16]), .B(s0[29]), .Z(n68) );
  EO U149 ( .A(s0[11]), .B(s0[24]), .Z(n69) );
  EO U150 ( .A(s0[17]), .B(s0[30]), .Z(n70) );
  EO U151 ( .A(s0[12]), .B(s0[25]), .Z(n71) );
  EO U152 ( .A(s0[18]), .B(s0[31]), .Z(n72) );
  EO U153 ( .A(s0[13]), .B(s0[26]), .Z(n73) );
  IV U154 ( .A(n89), .Z(n88) );
  IVA U155 ( .A(n92), .Z(n89) );
  IVA U156 ( .A(n92), .Z(n90) );
  IVA U157 ( .A(n92), .Z(n91) );
endmodule


module LOG_POLY_DW01_add_4 ( A, B, CI, SUM, CO );
  input [67:0] A;
  input [67:0] B;
  output [67:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230;

  IVP U2 ( .A(n55), .Z(n2) );
  IVP U3 ( .A(n160), .Z(n24) );
  IVP U4 ( .A(n59), .Z(n3) );
  IVP U5 ( .A(n100), .Z(n11) );
  IVP U6 ( .A(n64), .Z(n5) );
  IVP U7 ( .A(n54), .Z(n1) );
  IVP U8 ( .A(n113), .Z(n16) );
  IVP U9 ( .A(n106), .Z(n13) );
  IVP U10 ( .A(n109), .Z(n15) );
  IVP U11 ( .A(n121), .Z(n21) );
  IVP U12 ( .A(n125), .Z(n18) );
  IVP U13 ( .A(n180), .Z(n31) );
  IVP U14 ( .A(n171), .Z(n28) );
  IVP U15 ( .A(n143), .Z(n25) );
  IVP U16 ( .A(n122), .Z(n23) );
  IVP U17 ( .A(n176), .Z(n30) );
  IVP U18 ( .A(n148), .Z(n27) );
  IVP U19 ( .A(n194), .Z(n36) );
  IVP U20 ( .A(n201), .Z(n35) );
  IVP U21 ( .A(n195), .Z(n33) );
  IVP U22 ( .A(n191), .Z(n34) );
  IVP U23 ( .A(n203), .Z(n37) );
  IVP U24 ( .A(n179), .Z(n29) );
  IVP U25 ( .A(n166), .Z(n26) );
  IVP U26 ( .A(n130), .Z(n19) );
  IVP U27 ( .A(n123), .Z(n20) );
  IVP U28 ( .A(n112), .Z(n14) );
  IVP U29 ( .A(n85), .Z(n7) );
  IVP U30 ( .A(n97), .Z(n9) );
  IVP U31 ( .A(n91), .Z(n10) );
  IVP U32 ( .A(n101), .Z(n12) );
  IVP U33 ( .A(n86), .Z(n8) );
  IVP U34 ( .A(n82), .Z(n6) );
  IVP U35 ( .A(n177), .Z(n32) );
  IVP U36 ( .A(n110), .Z(n17) );
  IVP U37 ( .A(n77), .Z(n4) );
  IVP U38 ( .A(n132), .Z(n22) );
  IVP U39 ( .A(n225), .Z(n48) );
  IVP U40 ( .A(n222), .Z(n45) );
  IVP U41 ( .A(n224), .Z(n46) );
  IVP U42 ( .A(n216), .Z(n43) );
  IVP U43 ( .A(A[22]), .Z(n49) );
  IVP U44 ( .A(n205), .Z(n38) );
  IVP U45 ( .A(n154), .Z(n39) );
  IVP U46 ( .A(n211), .Z(n40) );
  IVP U47 ( .A(A[32]), .Z(n41) );
  IVP U48 ( .A(n219), .Z(n44) );
  IVP U49 ( .A(A[24]), .Z(n47) );
  IVP U50 ( .A(n229), .Z(n50) );
  IVP U51 ( .A(A[29]), .Z(n42) );
  ND2 U52 ( .A(A[21]), .B(B[21]), .Z(n229) );
  EO U53 ( .A(n51), .B(n52), .Z(SUM[65]) );
  EO U54 ( .A(B[65]), .B(A[65]), .Z(n52) );
  AO7 U55 ( .A(n53), .B(n2), .C(n54), .Z(n51) );
  EO U56 ( .A(n55), .B(n56), .Z(SUM[64]) );
  NR2 U57 ( .A(n1), .B(n53), .Z(n56) );
  NR2 U58 ( .A(B[64]), .B(A[64]), .Z(n53) );
  ND2 U59 ( .A(B[64]), .B(A[64]), .Z(n54) );
  AO7 U60 ( .A(n57), .B(n58), .C(n59), .Z(n55) );
  AO6 U61 ( .A(n60), .B(n61), .C(n4), .Z(n58) );
  AO7 U62 ( .A(n62), .B(n63), .C(n64), .Z(n60) );
  AO6 U63 ( .A(n65), .B(n6), .C(n66), .Z(n63) );
  AO7 U64 ( .A(n67), .B(n68), .C(n7), .Z(n65) );
  AO1 U65 ( .A(n69), .B(n70), .C(n71), .D(n72), .Z(n67) );
  AN2 U66 ( .A(n73), .B(n70), .Z(n72) );
  EN U67 ( .A(n74), .B(n75), .Z(SUM[63]) );
  NR2 U68 ( .A(n3), .B(n57), .Z(n75) );
  NR2 U69 ( .A(B[63]), .B(A[63]), .Z(n57) );
  ND2 U70 ( .A(B[63]), .B(A[63]), .Z(n59) );
  AO6 U71 ( .A(n61), .B(n76), .C(n4), .Z(n74) );
  EN U72 ( .A(n78), .B(n76), .Z(SUM[62]) );
  AO7 U73 ( .A(n62), .B(n79), .C(n64), .Z(n76) );
  ND2 U74 ( .A(n61), .B(n77), .Z(n78) );
  ND2 U75 ( .A(B[62]), .B(A[62]), .Z(n77) );
  OR2 U76 ( .A(B[62]), .B(A[62]), .Z(n61) );
  EN U77 ( .A(n79), .B(n80), .Z(SUM[61]) );
  NR2 U78 ( .A(n5), .B(n62), .Z(n80) );
  NR2 U79 ( .A(B[61]), .B(A[61]), .Z(n62) );
  ND2 U80 ( .A(B[61]), .B(A[61]), .Z(n64) );
  AO6 U81 ( .A(n6), .B(n81), .C(n66), .Z(n79) );
  EO U82 ( .A(n81), .B(n83), .Z(SUM[60]) );
  NR2 U83 ( .A(n66), .B(n82), .Z(n83) );
  NR2 U84 ( .A(B[60]), .B(A[60]), .Z(n82) );
  AN2 U85 ( .A(B[60]), .B(A[60]), .Z(n66) );
  AO7 U86 ( .A(n84), .B(n68), .C(n7), .Z(n81) );
  AO7 U87 ( .A(n86), .B(n87), .C(n88), .Z(n85) );
  AO6 U88 ( .A(n89), .B(n9), .C(n90), .Z(n87) );
  AO7 U89 ( .A(n91), .B(n92), .C(n93), .Z(n89) );
  ND4 U90 ( .A(n8), .B(n9), .C(n10), .D(n12), .Z(n68) );
  EO U91 ( .A(n94), .B(n95), .Z(SUM[59]) );
  AO6 U92 ( .A(n96), .B(n9), .C(n90), .Z(n95) );
  ND2 U93 ( .A(n8), .B(n88), .Z(n94) );
  ND2 U94 ( .A(B[59]), .B(A[59]), .Z(n88) );
  NR2 U95 ( .A(B[59]), .B(A[59]), .Z(n86) );
  EO U96 ( .A(n96), .B(n98), .Z(SUM[58]) );
  NR2 U97 ( .A(n90), .B(n97), .Z(n98) );
  NR2 U98 ( .A(B[58]), .B(A[58]), .Z(n97) );
  AN2 U99 ( .A(B[58]), .B(A[58]), .Z(n90) );
  AO7 U100 ( .A(n91), .B(n11), .C(n93), .Z(n96) );
  EO U101 ( .A(n11), .B(n99), .Z(SUM[57]) );
  ND2 U102 ( .A(n93), .B(n10), .Z(n99) );
  NR2 U103 ( .A(B[57]), .B(A[57]), .Z(n91) );
  ND2 U104 ( .A(B[57]), .B(A[57]), .Z(n93) );
  AO7 U105 ( .A(n101), .B(n84), .C(n92), .Z(n100) );
  EO U106 ( .A(n102), .B(n84), .Z(SUM[56]) );
  AO6 U107 ( .A(n103), .B(n70), .C(n71), .Z(n84) );
  AO7 U108 ( .A(n104), .B(n105), .C(n106), .Z(n71) );
  AO6 U109 ( .A(n107), .B(n14), .C(n108), .Z(n105) );
  AO7 U110 ( .A(n109), .B(n110), .C(n111), .Z(n107) );
  NR4 U111 ( .A(n104), .B(n112), .C(n109), .D(n113), .Z(n70) );
  ND2 U112 ( .A(n12), .B(n92), .Z(n102) );
  ND2 U113 ( .A(B[56]), .B(A[56]), .Z(n92) );
  NR2 U114 ( .A(B[56]), .B(A[56]), .Z(n101) );
  EN U115 ( .A(n114), .B(n115), .Z(SUM[55]) );
  NR2 U116 ( .A(n13), .B(n104), .Z(n115) );
  NR2 U117 ( .A(B[55]), .B(A[55]), .Z(n104) );
  ND2 U118 ( .A(B[55]), .B(A[55]), .Z(n106) );
  AO6 U119 ( .A(n14), .B(n116), .C(n108), .Z(n114) );
  EO U120 ( .A(n116), .B(n117), .Z(SUM[54]) );
  NR2 U121 ( .A(n108), .B(n112), .Z(n117) );
  NR2 U122 ( .A(B[54]), .B(A[54]), .Z(n112) );
  AN2 U123 ( .A(B[54]), .B(A[54]), .Z(n108) );
  AO7 U124 ( .A(n109), .B(n118), .C(n111), .Z(n116) );
  EO U125 ( .A(n119), .B(n118), .Z(SUM[53]) );
  AO6 U126 ( .A(n16), .B(n103), .C(n17), .Z(n118) );
  ND2 U127 ( .A(n15), .B(n111), .Z(n119) );
  ND2 U128 ( .A(B[53]), .B(A[53]), .Z(n111) );
  NR2 U129 ( .A(B[53]), .B(A[53]), .Z(n109) );
  EO U130 ( .A(n103), .B(n120), .Z(SUM[52]) );
  NR2 U131 ( .A(n17), .B(n113), .Z(n120) );
  NR2 U132 ( .A(B[52]), .B(A[52]), .Z(n113) );
  ND2 U133 ( .A(B[52]), .B(A[52]), .Z(n110) );
  OR2 U134 ( .A(n73), .B(n69), .Z(n103) );
  NR4 U135 ( .A(n121), .B(n122), .C(n123), .D(n124), .Z(n69) );
  OR2 U136 ( .A(n125), .B(n126), .Z(n124) );
  AO7 U137 ( .A(n125), .B(n127), .C(n128), .Z(n73) );
  AO6 U138 ( .A(n129), .B(n20), .C(n19), .Z(n127) );
  AO7 U139 ( .A(n121), .B(n131), .C(n132), .Z(n129) );
  EN U140 ( .A(n133), .B(n134), .Z(SUM[51]) );
  ND2 U141 ( .A(n128), .B(n18), .Z(n134) );
  NR2 U142 ( .A(B[51]), .B(A[51]), .Z(n125) );
  ND2 U143 ( .A(B[51]), .B(A[51]), .Z(n128) );
  AO7 U144 ( .A(n123), .B(n135), .C(n130), .Z(n133) );
  EO U145 ( .A(n136), .B(n135), .Z(SUM[50]) );
  AO6 U146 ( .A(n21), .B(n137), .C(n22), .Z(n135) );
  ND2 U147 ( .A(n20), .B(n130), .Z(n136) );
  ND2 U148 ( .A(B[50]), .B(A[50]), .Z(n130) );
  NR2 U149 ( .A(B[50]), .B(A[50]), .Z(n123) );
  EO U150 ( .A(n137), .B(n138), .Z(SUM[49]) );
  NR2 U151 ( .A(n22), .B(n121), .Z(n138) );
  NR2 U152 ( .A(B[49]), .B(A[49]), .Z(n121) );
  ND2 U153 ( .A(B[49]), .B(A[49]), .Z(n132) );
  AO7 U154 ( .A(n122), .B(n126), .C(n131), .Z(n137) );
  EO U155 ( .A(n139), .B(n126), .Z(SUM[48]) );
  AO6 U156 ( .A(n24), .B(n140), .C(n141), .Z(n126) );
  AO7 U157 ( .A(n142), .B(n143), .C(n144), .Z(n140) );
  AO6 U158 ( .A(n26), .B(n145), .C(n146), .Z(n142) );
  AO3 U159 ( .A(n147), .B(n148), .C(n149), .D(n150), .Z(n145) );
  OR4 U160 ( .A(n151), .B(n152), .C(n153), .D(n148), .Z(n149) );
  ND2 U161 ( .A(n154), .B(n155), .Z(n151) );
  AO6 U162 ( .A(n156), .B(n155), .C(n157), .Z(n147) );
  AO7 U163 ( .A(n152), .B(n158), .C(n159), .Z(n156) );
  ND2 U164 ( .A(n23), .B(n131), .Z(n139) );
  ND2 U165 ( .A(B[48]), .B(A[48]), .Z(n131) );
  NR2 U166 ( .A(B[48]), .B(A[48]), .Z(n122) );
  EO U167 ( .A(n161), .B(n162), .Z(SUM[47]) );
  NR2 U168 ( .A(n141), .B(n160), .Z(n162) );
  NR2 U169 ( .A(B[47]), .B(A[47]), .Z(n160) );
  AN2 U170 ( .A(B[47]), .B(A[47]), .Z(n141) );
  AO7 U171 ( .A(n143), .B(n163), .C(n144), .Z(n161) );
  EO U172 ( .A(n164), .B(n163), .Z(SUM[46]) );
  AO6 U173 ( .A(n26), .B(n165), .C(n146), .Z(n163) );
  ND2 U174 ( .A(n25), .B(n144), .Z(n164) );
  ND2 U175 ( .A(B[46]), .B(A[46]), .Z(n144) );
  NR2 U176 ( .A(B[46]), .B(A[46]), .Z(n143) );
  EO U177 ( .A(n165), .B(n167), .Z(SUM[45]) );
  NR2 U178 ( .A(n146), .B(n166), .Z(n167) );
  NR2 U179 ( .A(B[45]), .B(A[45]), .Z(n166) );
  AN2 U180 ( .A(B[45]), .B(A[45]), .Z(n146) );
  AO7 U181 ( .A(n148), .B(n168), .C(n150), .Z(n165) );
  EO U182 ( .A(n169), .B(n168), .Z(SUM[44]) );
  AO6 U183 ( .A(n170), .B(n155), .C(n157), .Z(n168) );
  AO7 U184 ( .A(n171), .B(n172), .C(n173), .Z(n157) );
  AO6 U185 ( .A(n174), .B(n29), .C(n175), .Z(n172) );
  AO7 U186 ( .A(n176), .B(n177), .C(n178), .Z(n174) );
  NR4 U187 ( .A(n171), .B(n179), .C(n176), .D(n180), .Z(n155) );
  ND2 U188 ( .A(n27), .B(n150), .Z(n169) );
  ND2 U189 ( .A(B[44]), .B(A[44]), .Z(n150) );
  NR2 U190 ( .A(B[44]), .B(A[44]), .Z(n148) );
  EO U191 ( .A(n181), .B(n182), .Z(SUM[43]) );
  AO6 U192 ( .A(n183), .B(n29), .C(n175), .Z(n182) );
  ND2 U193 ( .A(n28), .B(n173), .Z(n181) );
  ND2 U194 ( .A(B[43]), .B(A[43]), .Z(n173) );
  NR2 U195 ( .A(B[43]), .B(A[43]), .Z(n171) );
  EO U196 ( .A(n183), .B(n184), .Z(SUM[42]) );
  NR2 U197 ( .A(n175), .B(n179), .Z(n184) );
  NR2 U198 ( .A(B[42]), .B(A[42]), .Z(n179) );
  AN2 U199 ( .A(B[42]), .B(A[42]), .Z(n175) );
  AO7 U200 ( .A(n176), .B(n185), .C(n178), .Z(n183) );
  EO U201 ( .A(n186), .B(n185), .Z(SUM[41]) );
  AO6 U202 ( .A(n31), .B(n170), .C(n32), .Z(n185) );
  ND2 U203 ( .A(n30), .B(n178), .Z(n186) );
  ND2 U204 ( .A(B[41]), .B(A[41]), .Z(n178) );
  NR2 U205 ( .A(B[41]), .B(A[41]), .Z(n176) );
  EO U206 ( .A(n170), .B(n187), .Z(SUM[40]) );
  NR2 U207 ( .A(n32), .B(n180), .Z(n187) );
  NR2 U208 ( .A(B[40]), .B(A[40]), .Z(n180) );
  ND2 U209 ( .A(B[40]), .B(A[40]), .Z(n177) );
  AO7 U210 ( .A(n38), .B(n152), .C(n159), .Z(n170) );
  AO6 U211 ( .A(n33), .B(n188), .C(n189), .Z(n159) );
  AO7 U212 ( .A(n190), .B(n191), .C(n192), .Z(n188) );
  AO6 U213 ( .A(n35), .B(n36), .C(n193), .Z(n190) );
  ND4 U214 ( .A(n33), .B(n34), .C(n35), .D(n37), .Z(n152) );
  EO U215 ( .A(n196), .B(n197), .Z(SUM[39]) );
  NR2 U216 ( .A(n189), .B(n195), .Z(n197) );
  NR2 U217 ( .A(B[39]), .B(A[39]), .Z(n195) );
  AN2 U218 ( .A(B[39]), .B(A[39]), .Z(n189) );
  AO7 U219 ( .A(n191), .B(n198), .C(n192), .Z(n196) );
  EO U220 ( .A(n199), .B(n198), .Z(SUM[38]) );
  AO6 U221 ( .A(n35), .B(n200), .C(n193), .Z(n198) );
  ND2 U222 ( .A(n34), .B(n192), .Z(n199) );
  ND2 U223 ( .A(B[38]), .B(A[38]), .Z(n192) );
  NR2 U224 ( .A(B[38]), .B(A[38]), .Z(n191) );
  EO U225 ( .A(n200), .B(n202), .Z(SUM[37]) );
  NR2 U226 ( .A(n193), .B(n201), .Z(n202) );
  NR2 U227 ( .A(B[37]), .B(A[37]), .Z(n201) );
  AN2 U228 ( .A(B[37]), .B(A[37]), .Z(n193) );
  AO7 U229 ( .A(n203), .B(n38), .C(n194), .Z(n200) );
  EO U230 ( .A(n204), .B(n38), .Z(SUM[36]) );
  AO7 U231 ( .A(n153), .B(n39), .C(n158), .Z(n205) );
  AO2 U232 ( .A(A[35]), .B(B[35]), .C(n40), .D(n206), .Z(n158) );
  EON1 U233 ( .A(n207), .B(n208), .C(B[34]), .D(A[34]), .Z(n206) );
  AO2 U234 ( .A(A[33]), .B(B[33]), .C(B[32]), .D(n209), .Z(n207) );
  NR2 U235 ( .A(n41), .B(n210), .Z(n209) );
  NR4 U236 ( .A(n212), .B(n211), .C(n208), .D(n210), .Z(n154) );
  NR2 U237 ( .A(B[33]), .B(A[33]), .Z(n210) );
  NR2 U238 ( .A(B[34]), .B(A[34]), .Z(n208) );
  NR2 U239 ( .A(B[35]), .B(A[35]), .Z(n211) );
  NR2 U240 ( .A(B[32]), .B(A[32]), .Z(n212) );
  EO1 U241 ( .A(A[31]), .B(B[31]), .C(n213), .D(n214), .Z(n153) );
  AO5 U242 ( .A(A[30]), .B(B[30]), .C(n215), .Z(n214) );
  AO7 U243 ( .A(n216), .B(n42), .C(n217), .Z(n215) );
  AO7 U244 ( .A(A[29]), .B(n43), .C(B[29]), .Z(n217) );
  AO6 U245 ( .A(n218), .B(A[28]), .C(n44), .Z(n216) );
  AO7 U246 ( .A(A[28]), .B(n218), .C(B[28]), .Z(n219) );
  EON1 U247 ( .A(n220), .B(n221), .C(A[27]), .D(B[27]), .Z(n218) );
  AO5 U248 ( .A(A[26]), .B(B[26]), .C(n45), .Z(n221) );
  AO6 U249 ( .A(n223), .B(A[25]), .C(n46), .Z(n222) );
  AO7 U250 ( .A(A[25]), .B(n223), .C(B[25]), .Z(n224) );
  AO7 U251 ( .A(n225), .B(n47), .C(n226), .Z(n223) );
  AO7 U252 ( .A(A[24]), .B(n48), .C(B[24]), .Z(n226) );
  AO2 U253 ( .A(n227), .B(A[23]), .C(B[23]), .D(n228), .Z(n225) );
  OR2 U254 ( .A(n227), .B(A[23]), .Z(n228) );
  AO7 U255 ( .A(n229), .B(n49), .C(n230), .Z(n227) );
  AO7 U256 ( .A(A[22]), .B(n50), .C(B[22]), .Z(n230) );
  NR2 U257 ( .A(A[27]), .B(B[27]), .Z(n220) );
  NR2 U258 ( .A(A[31]), .B(B[31]), .Z(n213) );
  ND2 U259 ( .A(n37), .B(n194), .Z(n204) );
  ND2 U260 ( .A(B[36]), .B(A[36]), .Z(n194) );
  NR2 U261 ( .A(B[36]), .B(A[36]), .Z(n203) );
endmodule


module LOG_POLY_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [21:0] A;
  input [47:0] B;
  output [69:0] PRODUCT;
  input TC;
  wire   \ab[21][47] , \ab[21][46] , \ab[21][45] , \ab[21][44] , \ab[21][43] ,
         \ab[21][42] , \ab[21][41] , \ab[21][40] , \ab[21][39] , \ab[21][38] ,
         \ab[21][37] , \ab[21][36] , \ab[21][35] , \ab[21][34] , \ab[21][33] ,
         \ab[21][32] , \ab[21][31] , \ab[21][30] , \ab[21][29] , \ab[21][28] ,
         \ab[21][27] , \ab[21][26] , \ab[21][25] , \ab[21][24] , \ab[21][23] ,
         \ab[21][22] , \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] ,
         \ab[21][17] , \ab[21][16] , \ab[21][15] , \ab[21][14] , \ab[21][13] ,
         \ab[21][12] , \ab[21][11] , \ab[21][10] , \ab[21][9] , \ab[21][8] ,
         \ab[21][7] , \ab[21][6] , \ab[21][5] , \ab[21][4] , \ab[21][3] ,
         \ab[21][2] , \ab[21][1] , \ab[21][0] , \ab[20][47] , \ab[20][46] ,
         \ab[20][45] , \ab[20][44] , \ab[20][43] , \ab[20][42] , \ab[20][41] ,
         \ab[20][40] , \ab[20][39] , \ab[20][38] , \ab[20][37] , \ab[20][36] ,
         \ab[20][35] , \ab[20][34] , \ab[20][33] , \ab[20][32] , \ab[20][31] ,
         \ab[20][30] , \ab[20][29] , \ab[20][28] , \ab[20][27] , \ab[20][26] ,
         \ab[20][25] , \ab[20][24] , \ab[20][23] , \ab[20][22] , \ab[20][21] ,
         \ab[20][20] , \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] ,
         \ab[20][15] , \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] ,
         \ab[20][10] , \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] ,
         \ab[20][5] , \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] ,
         \ab[20][0] , \ab[19][47] , \ab[19][46] , \ab[19][45] , \ab[19][44] ,
         \ab[19][43] , \ab[19][42] , \ab[19][41] , \ab[19][40] , \ab[19][39] ,
         \ab[19][38] , \ab[19][37] , \ab[19][36] , \ab[19][35] , \ab[19][34] ,
         \ab[19][33] , \ab[19][32] , \ab[19][31] , \ab[19][30] , \ab[19][29] ,
         \ab[19][28] , \ab[19][27] , \ab[19][26] , \ab[19][25] , \ab[19][24] ,
         \ab[19][23] , \ab[19][22] , \ab[19][21] , \ab[19][20] , \ab[19][19] ,
         \ab[19][18] , \ab[19][17] , \ab[19][16] , \ab[19][15] , \ab[19][14] ,
         \ab[19][13] , \ab[19][12] , \ab[19][11] , \ab[19][10] , \ab[19][9] ,
         \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] , \ab[19][4] ,
         \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] , \ab[18][47] ,
         \ab[18][46] , \ab[18][45] , \ab[18][44] , \ab[18][43] , \ab[18][42] ,
         \ab[18][41] , \ab[18][40] , \ab[18][39] , \ab[18][38] , \ab[18][37] ,
         \ab[18][36] , \ab[18][35] , \ab[18][34] , \ab[18][33] , \ab[18][32] ,
         \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] , \ab[18][27] ,
         \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] , \ab[18][22] ,
         \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] , \ab[18][17] ,
         \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] , \ab[18][12] ,
         \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] , \ab[18][7] ,
         \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] , \ab[18][2] ,
         \ab[18][1] , \ab[18][0] , \ab[17][47] , \ab[17][46] , \ab[17][45] ,
         \ab[17][44] , \ab[17][43] , \ab[17][42] , \ab[17][41] , \ab[17][40] ,
         \ab[17][39] , \ab[17][38] , \ab[17][37] , \ab[17][36] , \ab[17][35] ,
         \ab[17][34] , \ab[17][33] , \ab[17][32] , \ab[17][31] , \ab[17][30] ,
         \ab[17][29] , \ab[17][28] , \ab[17][27] , \ab[17][26] , \ab[17][25] ,
         \ab[17][24] , \ab[17][23] , \ab[17][22] , \ab[17][21] , \ab[17][20] ,
         \ab[17][19] , \ab[17][18] , \ab[17][17] , \ab[17][16] , \ab[17][15] ,
         \ab[17][14] , \ab[17][13] , \ab[17][12] , \ab[17][11] , \ab[17][10] ,
         \ab[17][9] , \ab[17][8] , \ab[17][7] , \ab[17][6] , \ab[17][5] ,
         \ab[17][4] , \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] ,
         \ab[16][47] , \ab[16][46] , \ab[16][45] , \ab[16][44] , \ab[16][43] ,
         \ab[16][42] , \ab[16][41] , \ab[16][40] , \ab[16][39] , \ab[16][38] ,
         \ab[16][37] , \ab[16][36] , \ab[16][35] , \ab[16][34] , \ab[16][33] ,
         \ab[16][32] , \ab[16][31] , \ab[16][30] , \ab[16][29] , \ab[16][28] ,
         \ab[16][27] , \ab[16][26] , \ab[16][25] , \ab[16][24] , \ab[16][23] ,
         \ab[16][22] , \ab[16][21] , \ab[16][20] , \ab[16][19] , \ab[16][18] ,
         \ab[16][17] , \ab[16][16] , \ab[16][15] , \ab[16][14] , \ab[16][13] ,
         \ab[16][12] , \ab[16][11] , \ab[16][10] , \ab[16][9] , \ab[16][8] ,
         \ab[16][7] , \ab[16][6] , \ab[16][5] , \ab[16][4] , \ab[16][3] ,
         \ab[16][2] , \ab[16][1] , \ab[16][0] , \ab[15][47] , \ab[15][46] ,
         \ab[15][45] , \ab[15][44] , \ab[15][43] , \ab[15][42] , \ab[15][41] ,
         \ab[15][40] , \ab[15][39] , \ab[15][38] , \ab[15][37] , \ab[15][36] ,
         \ab[15][35] , \ab[15][34] , \ab[15][33] , \ab[15][32] , \ab[15][31] ,
         \ab[15][30] , \ab[15][29] , \ab[15][28] , \ab[15][27] , \ab[15][26] ,
         \ab[15][25] , \ab[15][24] , \ab[15][23] , \ab[15][22] , \ab[15][21] ,
         \ab[15][20] , \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] ,
         \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][47] , \ab[14][46] , \ab[14][45] , \ab[14][44] ,
         \ab[14][43] , \ab[14][42] , \ab[14][41] , \ab[14][40] , \ab[14][39] ,
         \ab[14][38] , \ab[14][37] , \ab[14][36] , \ab[14][35] , \ab[14][34] ,
         \ab[14][33] , \ab[14][32] , \ab[14][31] , \ab[14][30] , \ab[14][29] ,
         \ab[14][28] , \ab[14][27] , \ab[14][26] , \ab[14][25] , \ab[14][24] ,
         \ab[14][23] , \ab[14][22] , \ab[14][21] , \ab[14][20] , \ab[14][19] ,
         \ab[14][18] , \ab[14][17] , \ab[14][16] , \ab[14][15] , \ab[14][14] ,
         \ab[14][13] , \ab[14][12] , \ab[14][11] , \ab[14][10] , \ab[14][9] ,
         \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] ,
         \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][47] ,
         \ab[13][46] , \ab[13][45] , \ab[13][44] , \ab[13][43] , \ab[13][42] ,
         \ab[13][41] , \ab[13][40] , \ab[13][39] , \ab[13][38] , \ab[13][37] ,
         \ab[13][36] , \ab[13][35] , \ab[13][34] , \ab[13][33] , \ab[13][32] ,
         \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] , \ab[13][27] ,
         \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] , \ab[13][22] ,
         \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] , \ab[13][17] ,
         \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] , \ab[13][12] ,
         \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] , \ab[13][7] ,
         \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] , \ab[13][2] ,
         \ab[13][1] , \ab[13][0] , \ab[12][47] , \ab[12][46] , \ab[12][45] ,
         \ab[12][44] , \ab[12][43] , \ab[12][42] , \ab[12][41] , \ab[12][40] ,
         \ab[12][39] , \ab[12][38] , \ab[12][37] , \ab[12][36] , \ab[12][35] ,
         \ab[12][34] , \ab[12][33] , \ab[12][32] , \ab[12][31] , \ab[12][30] ,
         \ab[12][29] , \ab[12][28] , \ab[12][27] , \ab[12][26] , \ab[12][25] ,
         \ab[12][24] , \ab[12][23] , \ab[12][22] , \ab[12][21] , \ab[12][20] ,
         \ab[12][19] , \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][47] , \ab[11][46] , \ab[11][45] , \ab[11][44] , \ab[11][43] ,
         \ab[11][42] , \ab[11][41] , \ab[11][40] , \ab[11][39] , \ab[11][38] ,
         \ab[11][37] , \ab[11][36] , \ab[11][35] , \ab[11][34] , \ab[11][33] ,
         \ab[11][32] , \ab[11][31] , \ab[11][30] , \ab[11][29] , \ab[11][28] ,
         \ab[11][27] , \ab[11][26] , \ab[11][25] , \ab[11][24] , \ab[11][23] ,
         \ab[11][22] , \ab[11][21] , \ab[11][20] , \ab[11][19] , \ab[11][18] ,
         \ab[11][17] , \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] ,
         \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] ,
         \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] ,
         \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][47] , \ab[10][46] ,
         \ab[10][45] , \ab[10][44] , \ab[10][43] , \ab[10][42] , \ab[10][41] ,
         \ab[10][40] , \ab[10][39] , \ab[10][38] , \ab[10][37] , \ab[10][36] ,
         \ab[10][35] , \ab[10][34] , \ab[10][33] , \ab[10][32] , \ab[10][31] ,
         \ab[10][30] , \ab[10][29] , \ab[10][28] , \ab[10][27] , \ab[10][26] ,
         \ab[10][25] , \ab[10][24] , \ab[10][23] , \ab[10][22] , \ab[10][21] ,
         \ab[10][20] , \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][47] , \ab[9][46] , \ab[9][45] , \ab[9][44] ,
         \ab[9][43] , \ab[9][42] , \ab[9][41] , \ab[9][40] , \ab[9][39] ,
         \ab[9][38] , \ab[9][37] , \ab[9][36] , \ab[9][35] , \ab[9][34] ,
         \ab[9][33] , \ab[9][32] , \ab[9][31] , \ab[9][30] , \ab[9][29] ,
         \ab[9][28] , \ab[9][27] , \ab[9][26] , \ab[9][25] , \ab[9][24] ,
         \ab[9][23] , \ab[9][22] , \ab[9][21] , \ab[9][20] , \ab[9][19] ,
         \ab[9][18] , \ab[9][17] , \ab[9][16] , \ab[9][15] , \ab[9][14] ,
         \ab[9][13] , \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] ,
         \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] ,
         \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][47] ,
         \ab[8][46] , \ab[8][45] , \ab[8][44] , \ab[8][43] , \ab[8][42] ,
         \ab[8][41] , \ab[8][40] , \ab[8][39] , \ab[8][38] , \ab[8][37] ,
         \ab[8][36] , \ab[8][35] , \ab[8][34] , \ab[8][33] , \ab[8][32] ,
         \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] , \ab[8][27] ,
         \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] , \ab[8][22] ,
         \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] , \ab[8][17] ,
         \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] , \ab[8][12] ,
         \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] ,
         \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] ,
         \ab[8][1] , \ab[8][0] , \ab[7][47] , \ab[7][46] , \ab[7][45] ,
         \ab[7][44] , \ab[7][43] , \ab[7][42] , \ab[7][41] , \ab[7][40] ,
         \ab[7][39] , \ab[7][38] , \ab[7][37] , \ab[7][36] , \ab[7][35] ,
         \ab[7][34] , \ab[7][33] , \ab[7][32] , \ab[7][31] , \ab[7][30] ,
         \ab[7][29] , \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][47] , \ab[6][46] , \ab[6][45] , \ab[6][44] , \ab[6][43] ,
         \ab[6][42] , \ab[6][41] , \ab[6][40] , \ab[6][39] , \ab[6][38] ,
         \ab[6][37] , \ab[6][36] , \ab[6][35] , \ab[6][34] , \ab[6][33] ,
         \ab[6][32] , \ab[6][31] , \ab[6][30] , \ab[6][29] , \ab[6][28] ,
         \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] , \ab[6][23] ,
         \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] , \ab[6][18] ,
         \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] ,
         \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] ,
         \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] ,
         \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][47] , \ab[5][46] ,
         \ab[5][45] , \ab[5][44] , \ab[5][43] , \ab[5][42] , \ab[5][41] ,
         \ab[5][40] , \ab[5][39] , \ab[5][38] , \ab[5][37] , \ab[5][36] ,
         \ab[5][35] , \ab[5][34] , \ab[5][33] , \ab[5][32] , \ab[5][31] ,
         \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] ,
         \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][47] , \ab[4][46] , \ab[4][45] , \ab[4][44] ,
         \ab[4][43] , \ab[4][42] , \ab[4][41] , \ab[4][40] , \ab[4][39] ,
         \ab[4][38] , \ab[4][37] , \ab[4][36] , \ab[4][35] , \ab[4][34] ,
         \ab[4][33] , \ab[4][32] , \ab[4][31] , \ab[4][30] , \ab[4][29] ,
         \ab[4][28] , \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] ,
         \ab[4][23] , \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] ,
         \ab[4][18] , \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] ,
         \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] ,
         \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] ,
         \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][47] ,
         \ab[3][46] , \ab[3][45] , \ab[3][44] , \ab[3][43] , \ab[3][42] ,
         \ab[3][41] , \ab[3][40] , \ab[3][39] , \ab[3][38] , \ab[3][37] ,
         \ab[3][36] , \ab[3][35] , \ab[3][34] , \ab[3][33] , \ab[3][32] ,
         \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] , \ab[3][27] ,
         \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] , \ab[3][22] ,
         \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] , \ab[3][17] ,
         \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] , \ab[3][12] ,
         \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] ,
         \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] ,
         \ab[3][1] , \ab[3][0] , \ab[2][47] , \ab[2][46] , \ab[2][45] ,
         \ab[2][44] , \ab[2][43] , \ab[2][42] , \ab[2][41] , \ab[2][40] ,
         \ab[2][39] , \ab[2][38] , \ab[2][37] , \ab[2][36] , \ab[2][35] ,
         \ab[2][34] , \ab[2][33] , \ab[2][32] , \ab[2][31] , \ab[2][30] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][47] , \ab[1][46] , \ab[1][45] , \ab[1][44] , \ab[1][43] ,
         \ab[1][42] , \ab[1][41] , \ab[1][40] , \ab[1][39] , \ab[1][38] ,
         \ab[1][37] , \ab[1][36] , \ab[1][35] , \ab[1][34] , \ab[1][33] ,
         \ab[1][32] , \ab[1][31] , \ab[1][30] , \ab[1][29] , \ab[1][28] ,
         \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] , \ab[1][23] ,
         \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] ,
         \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[0][47] , \ab[0][46] , \ab[0][45] ,
         \ab[0][44] , \ab[0][43] , \ab[0][42] , \ab[0][41] , \ab[0][40] ,
         \ab[0][39] , \ab[0][38] , \ab[0][37] , \ab[0][36] , \ab[0][35] ,
         \ab[0][34] , \ab[0][33] , \ab[0][32] , \ab[0][31] , \ab[0][30] ,
         \ab[0][29] , \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] ,
         \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] ,
         \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] ,
         \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \CARRYB[11][15] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][46] , \CARRYB[10][45] , \CARRYB[10][44] ,
         \CARRYB[10][43] , \CARRYB[10][42] , \CARRYB[10][41] ,
         \CARRYB[10][40] , \CARRYB[10][39] , \CARRYB[10][38] ,
         \CARRYB[10][37] , \CARRYB[10][36] , \CARRYB[10][35] ,
         \CARRYB[10][34] , \CARRYB[10][33] , \CARRYB[10][32] ,
         \CARRYB[10][31] , \CARRYB[10][30] , \CARRYB[10][29] ,
         \CARRYB[10][28] , \CARRYB[10][27] , \CARRYB[10][26] ,
         \CARRYB[10][25] , \CARRYB[10][24] , \CARRYB[10][23] ,
         \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][46] ,
         \CARRYB[9][45] , \CARRYB[9][44] , \CARRYB[9][43] , \CARRYB[9][42] ,
         \CARRYB[9][41] , \CARRYB[9][40] , \CARRYB[9][39] , \CARRYB[9][38] ,
         \CARRYB[9][37] , \CARRYB[9][36] , \CARRYB[9][35] , \CARRYB[9][34] ,
         \CARRYB[9][33] , \CARRYB[9][32] , \CARRYB[9][31] , \CARRYB[9][30] ,
         \CARRYB[9][29] , \CARRYB[9][28] , \CARRYB[9][27] , \CARRYB[9][26] ,
         \CARRYB[9][25] , \CARRYB[9][24] , \CARRYB[9][23] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][46] , \CARRYB[8][45] ,
         \CARRYB[8][44] , \CARRYB[8][43] , \CARRYB[8][42] , \CARRYB[8][41] ,
         \CARRYB[8][40] , \CARRYB[8][39] , \CARRYB[8][38] , \CARRYB[8][37] ,
         \CARRYB[8][36] , \CARRYB[8][35] , \CARRYB[8][34] , \CARRYB[8][33] ,
         \CARRYB[8][32] , \CARRYB[8][31] , \CARRYB[8][30] , \CARRYB[8][29] ,
         \CARRYB[8][28] , \CARRYB[8][27] , \CARRYB[8][26] , \CARRYB[8][25] ,
         \CARRYB[8][24] , \CARRYB[8][23] , \CARRYB[8][22] , \CARRYB[8][21] ,
         \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] ,
         \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][46] , \CARRYB[7][45] , \CARRYB[7][44] ,
         \CARRYB[7][43] , \CARRYB[7][42] , \CARRYB[7][41] , \CARRYB[7][40] ,
         \CARRYB[7][39] , \CARRYB[7][38] , \CARRYB[7][37] , \CARRYB[7][36] ,
         \CARRYB[7][35] , \CARRYB[7][34] , \CARRYB[7][33] , \CARRYB[7][32] ,
         \CARRYB[7][31] , \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] ,
         \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] ,
         \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][46] , \CARRYB[6][45] , \CARRYB[6][44] , \CARRYB[6][43] ,
         \CARRYB[6][42] , \CARRYB[6][41] , \CARRYB[6][40] , \CARRYB[6][39] ,
         \CARRYB[6][38] , \CARRYB[6][37] , \CARRYB[6][36] , \CARRYB[6][35] ,
         \CARRYB[6][34] , \CARRYB[6][33] , \CARRYB[6][32] , \CARRYB[6][31] ,
         \CARRYB[6][30] , \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] ,
         \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][46] ,
         \CARRYB[5][45] , \CARRYB[5][44] , \CARRYB[5][43] , \CARRYB[5][42] ,
         \CARRYB[5][41] , \CARRYB[5][40] , \CARRYB[5][39] , \CARRYB[5][38] ,
         \CARRYB[5][37] , \CARRYB[5][36] , \CARRYB[5][35] , \CARRYB[5][34] ,
         \CARRYB[5][33] , \CARRYB[5][32] , \CARRYB[5][31] , \CARRYB[5][30] ,
         \CARRYB[5][29] , \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][46] , \CARRYB[4][45] ,
         \CARRYB[4][44] , \CARRYB[4][43] , \CARRYB[4][42] , \CARRYB[4][41] ,
         \CARRYB[4][40] , \CARRYB[4][39] , \CARRYB[4][38] , \CARRYB[4][37] ,
         \CARRYB[4][36] , \CARRYB[4][35] , \CARRYB[4][34] , \CARRYB[4][33] ,
         \CARRYB[4][32] , \CARRYB[4][31] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][46] , \CARRYB[3][45] , \CARRYB[3][44] ,
         \CARRYB[3][43] , \CARRYB[3][42] , \CARRYB[3][41] , \CARRYB[3][40] ,
         \CARRYB[3][39] , \CARRYB[3][38] , \CARRYB[3][37] , \CARRYB[3][36] ,
         \CARRYB[3][35] , \CARRYB[3][34] , \CARRYB[3][33] , \CARRYB[3][32] ,
         \CARRYB[3][31] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][46] , \CARRYB[2][45] , \CARRYB[2][44] , \CARRYB[2][43] ,
         \CARRYB[2][42] , \CARRYB[2][41] , \CARRYB[2][40] , \CARRYB[2][39] ,
         \CARRYB[2][38] , \CARRYB[2][37] , \CARRYB[2][36] , \CARRYB[2][35] ,
         \CARRYB[2][34] , \CARRYB[2][33] , \CARRYB[2][32] , \CARRYB[2][31] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][46] ,
         \CARRYB[1][45] , \CARRYB[1][44] , \CARRYB[1][43] , \CARRYB[1][42] ,
         \CARRYB[1][41] , \CARRYB[1][40] , \CARRYB[1][39] , \CARRYB[1][38] ,
         \CARRYB[1][37] , \CARRYB[1][36] , \CARRYB[1][35] , \CARRYB[1][34] ,
         \CARRYB[1][33] , \CARRYB[1][32] , \CARRYB[1][31] , \CARRYB[1][30] ,
         \CARRYB[1][29] , \CARRYB[1][28] , \CARRYB[1][27] , \CARRYB[1][26] ,
         \CARRYB[1][25] , \CARRYB[1][24] , \CARRYB[1][23] , \CARRYB[1][22] ,
         \CARRYB[1][21] , \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] ,
         \CARRYB[1][17] , \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] ,
         \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] ,
         \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] ,
         \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] ,
         \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[11][15] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][46] , \SUMB[10][45] , \SUMB[10][44] ,
         \SUMB[10][43] , \SUMB[10][42] , \SUMB[10][41] , \SUMB[10][40] ,
         \SUMB[10][39] , \SUMB[10][38] , \SUMB[10][37] , \SUMB[10][36] ,
         \SUMB[10][35] , \SUMB[10][34] , \SUMB[10][33] , \SUMB[10][32] ,
         \SUMB[10][31] , \SUMB[10][30] , \SUMB[10][29] , \SUMB[10][28] ,
         \SUMB[10][27] , \SUMB[10][26] , \SUMB[10][25] , \SUMB[10][24] ,
         \SUMB[10][23] , \SUMB[10][22] , \SUMB[10][21] , \SUMB[10][20] ,
         \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] , \SUMB[10][16] ,
         \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] , \SUMB[10][12] ,
         \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] , \SUMB[10][8] ,
         \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] ,
         \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][46] ,
         \SUMB[9][45] , \SUMB[9][44] , \SUMB[9][43] , \SUMB[9][42] ,
         \SUMB[9][41] , \SUMB[9][40] , \SUMB[9][39] , \SUMB[9][38] ,
         \SUMB[9][37] , \SUMB[9][36] , \SUMB[9][35] , \SUMB[9][34] ,
         \SUMB[9][33] , \SUMB[9][32] , \SUMB[9][31] , \SUMB[9][30] ,
         \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] , \SUMB[9][26] ,
         \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] , \SUMB[9][22] ,
         \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] ,
         \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][46] ,
         \SUMB[8][45] , \SUMB[8][44] , \SUMB[8][43] , \SUMB[8][42] ,
         \SUMB[8][41] , \SUMB[8][40] , \SUMB[8][39] , \SUMB[8][38] ,
         \SUMB[8][37] , \SUMB[8][36] , \SUMB[8][35] , \SUMB[8][34] ,
         \SUMB[8][33] , \SUMB[8][32] , \SUMB[8][31] , \SUMB[8][30] ,
         \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] , \SUMB[8][26] ,
         \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] , \SUMB[8][22] ,
         \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] ,
         \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][46] ,
         \SUMB[7][45] , \SUMB[7][44] , \SUMB[7][43] , \SUMB[7][42] ,
         \SUMB[7][41] , \SUMB[7][40] , \SUMB[7][39] , \SUMB[7][38] ,
         \SUMB[7][37] , \SUMB[7][36] , \SUMB[7][35] , \SUMB[7][34] ,
         \SUMB[7][33] , \SUMB[7][32] , \SUMB[7][31] , \SUMB[7][30] ,
         \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] ,
         \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][46] ,
         \SUMB[6][45] , \SUMB[6][44] , \SUMB[6][43] , \SUMB[6][42] ,
         \SUMB[6][41] , \SUMB[6][40] , \SUMB[6][39] , \SUMB[6][38] ,
         \SUMB[6][37] , \SUMB[6][36] , \SUMB[6][35] , \SUMB[6][34] ,
         \SUMB[6][33] , \SUMB[6][32] , \SUMB[6][31] , \SUMB[6][30] ,
         \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][46] ,
         \SUMB[5][45] , \SUMB[5][44] , \SUMB[5][43] , \SUMB[5][42] ,
         \SUMB[5][41] , \SUMB[5][40] , \SUMB[5][39] , \SUMB[5][38] ,
         \SUMB[5][37] , \SUMB[5][36] , \SUMB[5][35] , \SUMB[5][34] ,
         \SUMB[5][33] , \SUMB[5][32] , \SUMB[5][31] , \SUMB[5][30] ,
         \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] ,
         \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][46] ,
         \SUMB[4][45] , \SUMB[4][44] , \SUMB[4][43] , \SUMB[4][42] ,
         \SUMB[4][41] , \SUMB[4][40] , \SUMB[4][39] , \SUMB[4][38] ,
         \SUMB[4][37] , \SUMB[4][36] , \SUMB[4][35] , \SUMB[4][34] ,
         \SUMB[4][33] , \SUMB[4][32] , \SUMB[4][31] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][46] ,
         \SUMB[3][45] , \SUMB[3][44] , \SUMB[3][43] , \SUMB[3][42] ,
         \SUMB[3][41] , \SUMB[3][40] , \SUMB[3][39] , \SUMB[3][38] ,
         \SUMB[3][37] , \SUMB[3][36] , \SUMB[3][35] , \SUMB[3][34] ,
         \SUMB[3][33] , \SUMB[3][32] , \SUMB[3][31] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][46] ,
         \SUMB[2][45] , \SUMB[2][44] , \SUMB[2][43] , \SUMB[2][42] ,
         \SUMB[2][41] , \SUMB[2][40] , \SUMB[2][39] , \SUMB[2][38] ,
         \SUMB[2][37] , \SUMB[2][36] , \SUMB[2][35] , \SUMB[2][34] ,
         \SUMB[2][33] , \SUMB[2][32] , \SUMB[2][31] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][46] ,
         \SUMB[1][45] , \SUMB[1][44] , \SUMB[1][43] , \SUMB[1][42] ,
         \SUMB[1][41] , \SUMB[1][40] , \SUMB[1][39] , \SUMB[1][38] ,
         \SUMB[1][37] , \SUMB[1][36] , \SUMB[1][35] , \SUMB[1][34] ,
         \SUMB[1][33] , \SUMB[1][32] , \SUMB[1][31] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[21][46] , \CARRYB[21][45] , \CARRYB[21][44] ,
         \CARRYB[21][43] , \CARRYB[21][42] , \CARRYB[21][41] ,
         \CARRYB[21][40] , \CARRYB[21][39] , \CARRYB[21][38] ,
         \CARRYB[21][37] , \CARRYB[21][36] , \CARRYB[21][35] ,
         \CARRYB[21][34] , \CARRYB[21][33] , \CARRYB[21][32] ,
         \CARRYB[21][31] , \CARRYB[21][30] , \CARRYB[21][29] ,
         \CARRYB[21][28] , \CARRYB[21][27] , \CARRYB[21][26] ,
         \CARRYB[21][25] , \CARRYB[21][24] , \CARRYB[21][23] ,
         \CARRYB[21][22] , \CARRYB[21][21] , \CARRYB[21][20] ,
         \CARRYB[21][19] , \CARRYB[21][18] , \CARRYB[21][17] ,
         \CARRYB[21][16] , \CARRYB[21][15] , \CARRYB[21][14] ,
         \CARRYB[21][13] , \CARRYB[21][12] , \CARRYB[21][11] ,
         \CARRYB[21][10] , \CARRYB[21][9] , \CARRYB[21][8] , \CARRYB[21][7] ,
         \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] , \CARRYB[21][3] ,
         \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] , \CARRYB[20][46] ,
         \CARRYB[20][45] , \CARRYB[20][44] , \CARRYB[20][43] ,
         \CARRYB[20][42] , \CARRYB[20][41] , \CARRYB[20][40] ,
         \CARRYB[20][39] , \CARRYB[20][38] , \CARRYB[20][37] ,
         \CARRYB[20][36] , \CARRYB[20][35] , \CARRYB[20][34] ,
         \CARRYB[20][33] , \CARRYB[20][32] , \CARRYB[20][31] ,
         \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][46] , \CARRYB[19][45] , \CARRYB[19][44] ,
         \CARRYB[19][43] , \CARRYB[19][42] , \CARRYB[19][41] ,
         \CARRYB[19][40] , \CARRYB[19][39] , \CARRYB[19][38] ,
         \CARRYB[19][37] , \CARRYB[19][36] , \CARRYB[19][35] ,
         \CARRYB[19][34] , \CARRYB[19][33] , \CARRYB[19][32] ,
         \CARRYB[19][31] , \CARRYB[19][30] , \CARRYB[19][29] ,
         \CARRYB[19][28] , \CARRYB[19][27] , \CARRYB[19][26] ,
         \CARRYB[19][25] , \CARRYB[19][24] , \CARRYB[19][23] ,
         \CARRYB[19][22] , \CARRYB[19][21] , \CARRYB[19][20] ,
         \CARRYB[19][19] , \CARRYB[19][18] , \CARRYB[19][17] ,
         \CARRYB[19][16] , \CARRYB[19][15] , \CARRYB[19][14] ,
         \CARRYB[19][13] , \CARRYB[19][12] , \CARRYB[19][11] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][46] ,
         \CARRYB[18][45] , \CARRYB[18][44] , \CARRYB[18][43] ,
         \CARRYB[18][42] , \CARRYB[18][41] , \CARRYB[18][40] ,
         \CARRYB[18][39] , \CARRYB[18][38] , \CARRYB[18][37] ,
         \CARRYB[18][36] , \CARRYB[18][35] , \CARRYB[18][34] ,
         \CARRYB[18][33] , \CARRYB[18][32] , \CARRYB[18][31] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][46] , \CARRYB[17][45] , \CARRYB[17][44] ,
         \CARRYB[17][43] , \CARRYB[17][42] , \CARRYB[17][41] ,
         \CARRYB[17][40] , \CARRYB[17][39] , \CARRYB[17][38] ,
         \CARRYB[17][37] , \CARRYB[17][36] , \CARRYB[17][35] ,
         \CARRYB[17][34] , \CARRYB[17][33] , \CARRYB[17][32] ,
         \CARRYB[17][31] , \CARRYB[17][30] , \CARRYB[17][29] ,
         \CARRYB[17][28] , \CARRYB[17][27] , \CARRYB[17][26] ,
         \CARRYB[17][25] , \CARRYB[17][24] , \CARRYB[17][23] ,
         \CARRYB[17][22] , \CARRYB[17][21] , \CARRYB[17][20] ,
         \CARRYB[17][19] , \CARRYB[17][18] , \CARRYB[17][17] ,
         \CARRYB[17][16] , \CARRYB[17][15] , \CARRYB[17][14] ,
         \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][46] ,
         \CARRYB[16][45] , \CARRYB[16][44] , \CARRYB[16][43] ,
         \CARRYB[16][42] , \CARRYB[16][41] , \CARRYB[16][40] ,
         \CARRYB[16][39] , \CARRYB[16][38] , \CARRYB[16][37] ,
         \CARRYB[16][36] , \CARRYB[16][35] , \CARRYB[16][34] ,
         \CARRYB[16][33] , \CARRYB[16][32] , \CARRYB[16][31] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \CARRYB[15][46] , \CARRYB[15][45] , \CARRYB[15][44] ,
         \CARRYB[15][43] , \CARRYB[15][42] , \CARRYB[15][41] ,
         \CARRYB[15][40] , \CARRYB[15][39] , \CARRYB[15][38] ,
         \CARRYB[15][37] , \CARRYB[15][36] , \CARRYB[15][35] ,
         \CARRYB[15][34] , \CARRYB[15][33] , \CARRYB[15][32] ,
         \CARRYB[15][31] , \CARRYB[15][30] , \CARRYB[15][29] ,
         \CARRYB[15][28] , \CARRYB[15][27] , \CARRYB[15][26] ,
         \CARRYB[15][25] , \CARRYB[15][24] , \CARRYB[15][23] ,
         \CARRYB[15][22] , \CARRYB[15][21] , \CARRYB[15][20] ,
         \CARRYB[15][19] , \CARRYB[15][18] , \CARRYB[15][17] ,
         \CARRYB[15][16] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][46] ,
         \CARRYB[14][45] , \CARRYB[14][44] , \CARRYB[14][43] ,
         \CARRYB[14][42] , \CARRYB[14][41] , \CARRYB[14][40] ,
         \CARRYB[14][39] , \CARRYB[14][38] , \CARRYB[14][37] ,
         \CARRYB[14][36] , \CARRYB[14][35] , \CARRYB[14][34] ,
         \CARRYB[14][33] , \CARRYB[14][32] , \CARRYB[14][31] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][46] , \CARRYB[13][45] , \CARRYB[13][44] ,
         \CARRYB[13][43] , \CARRYB[13][42] , \CARRYB[13][41] ,
         \CARRYB[13][40] , \CARRYB[13][39] , \CARRYB[13][38] ,
         \CARRYB[13][37] , \CARRYB[13][36] , \CARRYB[13][35] ,
         \CARRYB[13][34] , \CARRYB[13][33] , \CARRYB[13][32] ,
         \CARRYB[13][31] , \CARRYB[13][30] , \CARRYB[13][29] ,
         \CARRYB[13][28] , \CARRYB[13][27] , \CARRYB[13][26] ,
         \CARRYB[13][25] , \CARRYB[13][24] , \CARRYB[13][23] ,
         \CARRYB[13][22] , \CARRYB[13][21] , \CARRYB[13][20] ,
         \CARRYB[13][19] , \CARRYB[13][18] , \CARRYB[13][17] ,
         \CARRYB[13][16] , \CARRYB[13][15] , \CARRYB[13][14] ,
         \CARRYB[13][13] , \CARRYB[13][12] , \CARRYB[13][11] ,
         \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] , \CARRYB[13][7] ,
         \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] , \CARRYB[13][3] ,
         \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] , \CARRYB[12][46] ,
         \CARRYB[12][45] , \CARRYB[12][44] , \CARRYB[12][43] ,
         \CARRYB[12][42] , \CARRYB[12][41] , \CARRYB[12][40] ,
         \CARRYB[12][39] , \CARRYB[12][38] , \CARRYB[12][37] ,
         \CARRYB[12][36] , \CARRYB[12][35] , \CARRYB[12][34] ,
         \CARRYB[12][33] , \CARRYB[12][32] , \CARRYB[12][31] ,
         \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][46] , \CARRYB[11][45] , \CARRYB[11][44] ,
         \CARRYB[11][43] , \CARRYB[11][42] , \CARRYB[11][41] ,
         \CARRYB[11][40] , \CARRYB[11][39] , \CARRYB[11][38] ,
         \CARRYB[11][37] , \CARRYB[11][36] , \CARRYB[11][35] ,
         \CARRYB[11][34] , \CARRYB[11][33] , \CARRYB[11][32] ,
         \CARRYB[11][31] , \CARRYB[11][30] , \CARRYB[11][29] ,
         \CARRYB[11][28] , \CARRYB[11][27] , \CARRYB[11][26] ,
         \CARRYB[11][25] , \CARRYB[11][24] , \CARRYB[11][23] ,
         \CARRYB[11][22] , \CARRYB[11][21] , \CARRYB[11][20] ,
         \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \SUMB[21][46] , \SUMB[21][45] , \SUMB[21][44] ,
         \SUMB[21][43] , \SUMB[21][42] , \SUMB[21][41] , \SUMB[21][40] ,
         \SUMB[21][39] , \SUMB[21][38] , \SUMB[21][37] , \SUMB[21][36] ,
         \SUMB[21][35] , \SUMB[21][34] , \SUMB[21][33] , \SUMB[21][32] ,
         \SUMB[21][31] , \SUMB[21][30] , \SUMB[21][29] , \SUMB[21][28] ,
         \SUMB[21][27] , \SUMB[21][26] , \SUMB[21][25] , \SUMB[21][24] ,
         \SUMB[21][23] , \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] ,
         \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] ,
         \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] ,
         \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] ,
         \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] ,
         \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] , \SUMB[21][0] ,
         \SUMB[20][46] , \SUMB[20][45] , \SUMB[20][44] , \SUMB[20][43] ,
         \SUMB[20][42] , \SUMB[20][41] , \SUMB[20][40] , \SUMB[20][39] ,
         \SUMB[20][38] , \SUMB[20][37] , \SUMB[20][36] , \SUMB[20][35] ,
         \SUMB[20][34] , \SUMB[20][33] , \SUMB[20][32] , \SUMB[20][31] ,
         \SUMB[20][30] , \SUMB[20][29] , \SUMB[20][28] , \SUMB[20][27] ,
         \SUMB[20][26] , \SUMB[20][25] , \SUMB[20][24] , \SUMB[20][23] ,
         \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] , \SUMB[20][19] ,
         \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] , \SUMB[20][15] ,
         \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] ,
         \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] ,
         \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] ,
         \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][46] , \SUMB[19][45] ,
         \SUMB[19][44] , \SUMB[19][43] , \SUMB[19][42] , \SUMB[19][41] ,
         \SUMB[19][40] , \SUMB[19][39] , \SUMB[19][38] , \SUMB[19][37] ,
         \SUMB[19][36] , \SUMB[19][35] , \SUMB[19][34] , \SUMB[19][33] ,
         \SUMB[19][32] , \SUMB[19][31] , \SUMB[19][30] , \SUMB[19][29] ,
         \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] , \SUMB[19][25] ,
         \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] , \SUMB[19][21] ,
         \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] ,
         \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] ,
         \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] ,
         \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] ,
         \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] ,
         \SUMB[18][46] , \SUMB[18][45] , \SUMB[18][44] , \SUMB[18][43] ,
         \SUMB[18][42] , \SUMB[18][41] , \SUMB[18][40] , \SUMB[18][39] ,
         \SUMB[18][38] , \SUMB[18][37] , \SUMB[18][36] , \SUMB[18][35] ,
         \SUMB[18][34] , \SUMB[18][33] , \SUMB[18][32] , \SUMB[18][31] ,
         \SUMB[18][30] , \SUMB[18][29] , \SUMB[18][28] , \SUMB[18][27] ,
         \SUMB[18][26] , \SUMB[18][25] , \SUMB[18][24] , \SUMB[18][23] ,
         \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] ,
         \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] ,
         \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] ,
         \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] ,
         \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][46] , \SUMB[17][45] ,
         \SUMB[17][44] , \SUMB[17][43] , \SUMB[17][42] , \SUMB[17][41] ,
         \SUMB[17][40] , \SUMB[17][39] , \SUMB[17][38] , \SUMB[17][37] ,
         \SUMB[17][36] , \SUMB[17][35] , \SUMB[17][34] , \SUMB[17][33] ,
         \SUMB[17][32] , \SUMB[17][31] , \SUMB[17][30] , \SUMB[17][29] ,
         \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] , \SUMB[17][25] ,
         \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] , \SUMB[17][21] ,
         \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] ,
         \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][46] , \SUMB[16][45] , \SUMB[16][44] , \SUMB[16][43] ,
         \SUMB[16][42] , \SUMB[16][41] , \SUMB[16][40] , \SUMB[16][39] ,
         \SUMB[16][38] , \SUMB[16][37] , \SUMB[16][36] , \SUMB[16][35] ,
         \SUMB[16][34] , \SUMB[16][33] , \SUMB[16][32] , \SUMB[16][31] ,
         \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] , \SUMB[16][27] ,
         \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] , \SUMB[16][23] ,
         \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][19] ,
         \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] , \SUMB[16][15] ,
         \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] ,
         \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] ,
         \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] ,
         \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][46] , \SUMB[15][45] ,
         \SUMB[15][44] , \SUMB[15][43] , \SUMB[15][42] , \SUMB[15][41] ,
         \SUMB[15][40] , \SUMB[15][39] , \SUMB[15][38] , \SUMB[15][37] ,
         \SUMB[15][36] , \SUMB[15][35] , \SUMB[15][34] , \SUMB[15][33] ,
         \SUMB[15][32] , \SUMB[15][31] , \SUMB[15][30] , \SUMB[15][29] ,
         \SUMB[15][28] , \SUMB[15][27] , \SUMB[15][26] , \SUMB[15][25] ,
         \SUMB[15][24] , \SUMB[15][23] , \SUMB[15][22] , \SUMB[15][21] ,
         \SUMB[15][20] , \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] ,
         \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][46] , \SUMB[14][45] , \SUMB[14][44] , \SUMB[14][43] ,
         \SUMB[14][42] , \SUMB[14][41] , \SUMB[14][40] , \SUMB[14][39] ,
         \SUMB[14][38] , \SUMB[14][37] , \SUMB[14][36] , \SUMB[14][35] ,
         \SUMB[14][34] , \SUMB[14][33] , \SUMB[14][32] , \SUMB[14][31] ,
         \SUMB[14][30] , \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] ,
         \SUMB[14][26] , \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] ,
         \SUMB[14][22] , \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] ,
         \SUMB[14][18] , \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] ,
         \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] ,
         \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] ,
         \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] ,
         \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][46] , \SUMB[13][45] ,
         \SUMB[13][44] , \SUMB[13][43] , \SUMB[13][42] , \SUMB[13][41] ,
         \SUMB[13][40] , \SUMB[13][39] , \SUMB[13][38] , \SUMB[13][37] ,
         \SUMB[13][36] , \SUMB[13][35] , \SUMB[13][34] , \SUMB[13][33] ,
         \SUMB[13][32] , \SUMB[13][31] , \SUMB[13][30] , \SUMB[13][29] ,
         \SUMB[13][28] , \SUMB[13][27] , \SUMB[13][26] , \SUMB[13][25] ,
         \SUMB[13][24] , \SUMB[13][23] , \SUMB[13][22] , \SUMB[13][21] ,
         \SUMB[13][20] , \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] ,
         \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][46] , \SUMB[12][45] , \SUMB[12][44] , \SUMB[12][43] ,
         \SUMB[12][42] , \SUMB[12][41] , \SUMB[12][40] , \SUMB[12][39] ,
         \SUMB[12][38] , \SUMB[12][37] , \SUMB[12][36] , \SUMB[12][35] ,
         \SUMB[12][34] , \SUMB[12][33] , \SUMB[12][32] , \SUMB[12][31] ,
         \SUMB[12][30] , \SUMB[12][29] , \SUMB[12][28] , \SUMB[12][27] ,
         \SUMB[12][26] , \SUMB[12][25] , \SUMB[12][24] , \SUMB[12][23] ,
         \SUMB[12][22] , \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] ,
         \SUMB[12][18] , \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] ,
         \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] ,
         \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] ,
         \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] ,
         \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][46] , \SUMB[11][45] ,
         \SUMB[11][44] , \SUMB[11][43] , \SUMB[11][42] , \SUMB[11][41] ,
         \SUMB[11][40] , \SUMB[11][39] , \SUMB[11][38] , \SUMB[11][37] ,
         \SUMB[11][36] , \SUMB[11][35] , \SUMB[11][34] , \SUMB[11][33] ,
         \SUMB[11][32] , \SUMB[11][31] , \SUMB[11][30] , \SUMB[11][29] ,
         \SUMB[11][28] , \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] ,
         \SUMB[11][24] , \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] ,
         \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] ,
         \SUMB[11][16] , \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] ,
         \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] ,
         \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] ,
         \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] ,
         \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] ,
         \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] ,
         \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] ,
         \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[67] , \A2[66] ,
         \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] ,
         \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] ,
         \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] ,
         \A2[23] , \A2[22] , \A2[21] , n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37;

  LOG_POLY_DW01_add_4 FS_1 ( .A({1'b0, \A1[66] , \A1[65] , \A1[64] , \A1[63] , 
        \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , 
        \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , 
        \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , 
        \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , 
        \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , 
        \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , 
        \A1[20] , \SUMB[21][0] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , 
        \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[67] , \A2[66] , \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , 
        \A2[60] , \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , 
        \A2[53] , \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , 
        \A2[46] , \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , 
        \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , 
        \A2[32] , \A2[31] , \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , 
        \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, PRODUCT[67:38], 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37}) );
  FA1A S3_20_46 ( .A(\ab[20][46] ), .B(\CARRYB[19][46] ), .CI(\ab[19][47] ), 
        .CO(\CARRYB[20][46] ), .S(\SUMB[20][46] ) );
  FA1A S3_19_46 ( .A(\ab[19][46] ), .B(\CARRYB[18][46] ), .CI(\ab[18][47] ), 
        .CO(\CARRYB[19][46] ), .S(\SUMB[19][46] ) );
  FA1A S3_18_46 ( .A(\ab[18][46] ), .B(\CARRYB[17][46] ), .CI(\ab[17][47] ), 
        .CO(\CARRYB[18][46] ), .S(\SUMB[18][46] ) );
  FA1A S3_17_46 ( .A(\ab[17][46] ), .B(\CARRYB[16][46] ), .CI(\ab[16][47] ), 
        .CO(\CARRYB[17][46] ), .S(\SUMB[17][46] ) );
  FA1A S3_16_46 ( .A(\ab[16][46] ), .B(\CARRYB[15][46] ), .CI(\ab[15][47] ), 
        .CO(\CARRYB[16][46] ), .S(\SUMB[16][46] ) );
  FA1A S3_15_46 ( .A(\ab[15][46] ), .B(\CARRYB[14][46] ), .CI(\ab[14][47] ), 
        .CO(\CARRYB[15][46] ), .S(\SUMB[15][46] ) );
  FA1A S3_14_46 ( .A(\ab[14][46] ), .B(\CARRYB[13][46] ), .CI(\ab[13][47] ), 
        .CO(\CARRYB[14][46] ), .S(\SUMB[14][46] ) );
  FA1A S3_13_46 ( .A(\ab[13][46] ), .B(\CARRYB[12][46] ), .CI(\ab[12][47] ), 
        .CO(\CARRYB[13][46] ), .S(\SUMB[13][46] ) );
  FA1A S3_12_46 ( .A(\ab[12][46] ), .B(\CARRYB[11][46] ), .CI(\ab[11][47] ), 
        .CO(\CARRYB[12][46] ), .S(\SUMB[12][46] ) );
  FA1A S3_11_46 ( .A(\ab[11][46] ), .B(\CARRYB[10][46] ), .CI(\ab[10][47] ), 
        .CO(\CARRYB[11][46] ), .S(\SUMB[11][46] ) );
  FA1A S3_10_46 ( .A(\ab[10][46] ), .B(\CARRYB[9][46] ), .CI(\ab[9][47] ), 
        .CO(\CARRYB[10][46] ), .S(\SUMB[10][46] ) );
  FA1A S3_9_46 ( .A(\ab[9][46] ), .B(\CARRYB[8][46] ), .CI(\ab[8][47] ), .CO(
        \CARRYB[9][46] ), .S(\SUMB[9][46] ) );
  FA1A S3_8_46 ( .A(\ab[8][46] ), .B(\CARRYB[7][46] ), .CI(\ab[7][47] ), .CO(
        \CARRYB[8][46] ), .S(\SUMB[8][46] ) );
  FA1A S3_7_46 ( .A(\ab[7][46] ), .B(\CARRYB[6][46] ), .CI(\ab[6][47] ), .CO(
        \CARRYB[7][46] ), .S(\SUMB[7][46] ) );
  FA1A S3_6_46 ( .A(\ab[6][46] ), .B(\CARRYB[5][46] ), .CI(\ab[5][47] ), .CO(
        \CARRYB[6][46] ), .S(\SUMB[6][46] ) );
  FA1A S3_5_46 ( .A(\ab[5][46] ), .B(\CARRYB[4][46] ), .CI(\ab[4][47] ), .CO(
        \CARRYB[5][46] ), .S(\SUMB[5][46] ) );
  FA1A S3_4_46 ( .A(\ab[4][46] ), .B(\CARRYB[3][46] ), .CI(\ab[3][47] ), .CO(
        \CARRYB[4][46] ), .S(\SUMB[4][46] ) );
  FA1A S3_3_46 ( .A(\ab[3][46] ), .B(\CARRYB[2][46] ), .CI(\ab[2][47] ), .CO(
        \CARRYB[3][46] ), .S(\SUMB[3][46] ) );
  FA1A S5_46 ( .A(\ab[21][46] ), .B(\CARRYB[20][46] ), .CI(\ab[20][47] ), .CO(
        \CARRYB[21][46] ), .S(\SUMB[21][46] ) );
  FA1A S2_20_45 ( .A(\ab[20][45] ), .B(\CARRYB[19][45] ), .CI(\SUMB[19][46] ), 
        .CO(\CARRYB[20][45] ), .S(\SUMB[20][45] ) );
  FA1A S2_19_45 ( .A(\ab[19][45] ), .B(\CARRYB[18][45] ), .CI(\SUMB[18][46] ), 
        .CO(\CARRYB[19][45] ), .S(\SUMB[19][45] ) );
  FA1A S2_18_45 ( .A(\ab[18][45] ), .B(\CARRYB[17][45] ), .CI(\SUMB[17][46] ), 
        .CO(\CARRYB[18][45] ), .S(\SUMB[18][45] ) );
  FA1A S2_17_45 ( .A(\ab[17][45] ), .B(\CARRYB[16][45] ), .CI(\SUMB[16][46] ), 
        .CO(\CARRYB[17][45] ), .S(\SUMB[17][45] ) );
  FA1A S2_16_45 ( .A(\ab[16][45] ), .B(\CARRYB[15][45] ), .CI(\SUMB[15][46] ), 
        .CO(\CARRYB[16][45] ), .S(\SUMB[16][45] ) );
  FA1A S2_15_45 ( .A(\ab[15][45] ), .B(\CARRYB[14][45] ), .CI(\SUMB[14][46] ), 
        .CO(\CARRYB[15][45] ), .S(\SUMB[15][45] ) );
  FA1A S2_14_45 ( .A(\ab[14][45] ), .B(\CARRYB[13][45] ), .CI(\SUMB[13][46] ), 
        .CO(\CARRYB[14][45] ), .S(\SUMB[14][45] ) );
  FA1A S2_13_45 ( .A(\ab[13][45] ), .B(\CARRYB[12][45] ), .CI(\SUMB[12][46] ), 
        .CO(\CARRYB[13][45] ), .S(\SUMB[13][45] ) );
  FA1A S2_12_45 ( .A(\ab[12][45] ), .B(\CARRYB[11][45] ), .CI(\SUMB[11][46] ), 
        .CO(\CARRYB[12][45] ), .S(\SUMB[12][45] ) );
  FA1A S2_11_45 ( .A(\ab[11][45] ), .B(\CARRYB[10][45] ), .CI(\SUMB[10][46] ), 
        .CO(\CARRYB[11][45] ), .S(\SUMB[11][45] ) );
  FA1A S2_10_45 ( .A(\ab[10][45] ), .B(\CARRYB[9][45] ), .CI(\SUMB[9][46] ), 
        .CO(\CARRYB[10][45] ), .S(\SUMB[10][45] ) );
  FA1A S2_9_45 ( .A(\ab[9][45] ), .B(\CARRYB[8][45] ), .CI(\SUMB[8][46] ), 
        .CO(\CARRYB[9][45] ), .S(\SUMB[9][45] ) );
  FA1A S2_8_45 ( .A(\ab[8][45] ), .B(\CARRYB[7][45] ), .CI(\SUMB[7][46] ), 
        .CO(\CARRYB[8][45] ), .S(\SUMB[8][45] ) );
  FA1A S2_7_45 ( .A(\ab[7][45] ), .B(\CARRYB[6][45] ), .CI(\SUMB[6][46] ), 
        .CO(\CARRYB[7][45] ), .S(\SUMB[7][45] ) );
  FA1A S2_6_45 ( .A(\ab[6][45] ), .B(\CARRYB[5][45] ), .CI(\SUMB[5][46] ), 
        .CO(\CARRYB[6][45] ), .S(\SUMB[6][45] ) );
  FA1A S2_5_45 ( .A(\ab[5][45] ), .B(\CARRYB[4][45] ), .CI(\SUMB[4][46] ), 
        .CO(\CARRYB[5][45] ), .S(\SUMB[5][45] ) );
  FA1A S2_4_45 ( .A(\ab[4][45] ), .B(\CARRYB[3][45] ), .CI(\SUMB[3][46] ), 
        .CO(\CARRYB[4][45] ), .S(\SUMB[4][45] ) );
  FA1A S2_3_45 ( .A(\ab[3][45] ), .B(\CARRYB[2][45] ), .CI(\SUMB[2][46] ), 
        .CO(\CARRYB[3][45] ), .S(\SUMB[3][45] ) );
  FA1A S3_2_46 ( .A(\ab[2][46] ), .B(\CARRYB[1][46] ), .CI(\ab[1][47] ), .CO(
        \CARRYB[2][46] ), .S(\SUMB[2][46] ) );
  FA1A S2_2_45 ( .A(\ab[2][45] ), .B(\CARRYB[1][45] ), .CI(\SUMB[1][46] ), 
        .CO(\CARRYB[2][45] ), .S(\SUMB[2][45] ) );
  FA1A S4_45 ( .A(\ab[21][45] ), .B(\CARRYB[20][45] ), .CI(\SUMB[20][46] ), 
        .CO(\CARRYB[21][45] ), .S(\SUMB[21][45] ) );
  FA1A S2_20_44 ( .A(\ab[20][44] ), .B(\CARRYB[19][44] ), .CI(\SUMB[19][45] ), 
        .CO(\CARRYB[20][44] ), .S(\SUMB[20][44] ) );
  FA1A S2_19_44 ( .A(\ab[19][44] ), .B(\CARRYB[18][44] ), .CI(\SUMB[18][45] ), 
        .CO(\CARRYB[19][44] ), .S(\SUMB[19][44] ) );
  FA1A S2_18_44 ( .A(\ab[18][44] ), .B(\CARRYB[17][44] ), .CI(\SUMB[17][45] ), 
        .CO(\CARRYB[18][44] ), .S(\SUMB[18][44] ) );
  FA1A S2_17_44 ( .A(\ab[17][44] ), .B(\CARRYB[16][44] ), .CI(\SUMB[16][45] ), 
        .CO(\CARRYB[17][44] ), .S(\SUMB[17][44] ) );
  FA1A S2_16_44 ( .A(\ab[16][44] ), .B(\CARRYB[15][44] ), .CI(\SUMB[15][45] ), 
        .CO(\CARRYB[16][44] ), .S(\SUMB[16][44] ) );
  FA1A S2_15_44 ( .A(\ab[15][44] ), .B(\CARRYB[14][44] ), .CI(\SUMB[14][45] ), 
        .CO(\CARRYB[15][44] ), .S(\SUMB[15][44] ) );
  FA1A S2_14_44 ( .A(\ab[14][44] ), .B(\CARRYB[13][44] ), .CI(\SUMB[13][45] ), 
        .CO(\CARRYB[14][44] ), .S(\SUMB[14][44] ) );
  FA1A S2_13_44 ( .A(\ab[13][44] ), .B(\CARRYB[12][44] ), .CI(\SUMB[12][45] ), 
        .CO(\CARRYB[13][44] ), .S(\SUMB[13][44] ) );
  FA1A S2_12_44 ( .A(\ab[12][44] ), .B(\CARRYB[11][44] ), .CI(\SUMB[11][45] ), 
        .CO(\CARRYB[12][44] ), .S(\SUMB[12][44] ) );
  FA1A S2_11_44 ( .A(\ab[11][44] ), .B(\CARRYB[10][44] ), .CI(\SUMB[10][45] ), 
        .CO(\CARRYB[11][44] ), .S(\SUMB[11][44] ) );
  FA1A S2_10_44 ( .A(\ab[10][44] ), .B(\CARRYB[9][44] ), .CI(\SUMB[9][45] ), 
        .CO(\CARRYB[10][44] ), .S(\SUMB[10][44] ) );
  FA1A S2_9_44 ( .A(\ab[9][44] ), .B(\CARRYB[8][44] ), .CI(\SUMB[8][45] ), 
        .CO(\CARRYB[9][44] ), .S(\SUMB[9][44] ) );
  FA1A S2_8_44 ( .A(\ab[8][44] ), .B(\CARRYB[7][44] ), .CI(\SUMB[7][45] ), 
        .CO(\CARRYB[8][44] ), .S(\SUMB[8][44] ) );
  FA1A S2_7_44 ( .A(\ab[7][44] ), .B(\CARRYB[6][44] ), .CI(\SUMB[6][45] ), 
        .CO(\CARRYB[7][44] ), .S(\SUMB[7][44] ) );
  FA1A S2_6_44 ( .A(\ab[6][44] ), .B(\CARRYB[5][44] ), .CI(\SUMB[5][45] ), 
        .CO(\CARRYB[6][44] ), .S(\SUMB[6][44] ) );
  FA1A S2_5_44 ( .A(\ab[5][44] ), .B(\CARRYB[4][44] ), .CI(\SUMB[4][45] ), 
        .CO(\CARRYB[5][44] ), .S(\SUMB[5][44] ) );
  FA1A S2_4_44 ( .A(\ab[4][44] ), .B(\CARRYB[3][44] ), .CI(\SUMB[3][45] ), 
        .CO(\CARRYB[4][44] ), .S(\SUMB[4][44] ) );
  FA1A S2_3_44 ( .A(\ab[3][44] ), .B(\CARRYB[2][44] ), .CI(\SUMB[2][45] ), 
        .CO(\CARRYB[3][44] ), .S(\SUMB[3][44] ) );
  FA1A S2_2_44 ( .A(\ab[2][44] ), .B(\CARRYB[1][44] ), .CI(\SUMB[1][45] ), 
        .CO(\CARRYB[2][44] ), .S(\SUMB[2][44] ) );
  FA1A S4_44 ( .A(\ab[21][44] ), .B(\CARRYB[20][44] ), .CI(\SUMB[20][45] ), 
        .CO(\CARRYB[21][44] ), .S(\SUMB[21][44] ) );
  FA1A S2_20_43 ( .A(\ab[20][43] ), .B(\CARRYB[19][43] ), .CI(\SUMB[19][44] ), 
        .CO(\CARRYB[20][43] ), .S(\SUMB[20][43] ) );
  FA1A S2_19_43 ( .A(\ab[19][43] ), .B(\CARRYB[18][43] ), .CI(\SUMB[18][44] ), 
        .CO(\CARRYB[19][43] ), .S(\SUMB[19][43] ) );
  FA1A S2_18_43 ( .A(\ab[18][43] ), .B(\CARRYB[17][43] ), .CI(\SUMB[17][44] ), 
        .CO(\CARRYB[18][43] ), .S(\SUMB[18][43] ) );
  FA1A S2_17_43 ( .A(\ab[17][43] ), .B(\CARRYB[16][43] ), .CI(\SUMB[16][44] ), 
        .CO(\CARRYB[17][43] ), .S(\SUMB[17][43] ) );
  FA1A S2_16_43 ( .A(\ab[16][43] ), .B(\CARRYB[15][43] ), .CI(\SUMB[15][44] ), 
        .CO(\CARRYB[16][43] ), .S(\SUMB[16][43] ) );
  FA1A S2_15_43 ( .A(\ab[15][43] ), .B(\CARRYB[14][43] ), .CI(\SUMB[14][44] ), 
        .CO(\CARRYB[15][43] ), .S(\SUMB[15][43] ) );
  FA1A S2_14_43 ( .A(\ab[14][43] ), .B(\CARRYB[13][43] ), .CI(\SUMB[13][44] ), 
        .CO(\CARRYB[14][43] ), .S(\SUMB[14][43] ) );
  FA1A S2_13_43 ( .A(\ab[13][43] ), .B(\CARRYB[12][43] ), .CI(\SUMB[12][44] ), 
        .CO(\CARRYB[13][43] ), .S(\SUMB[13][43] ) );
  FA1A S2_12_43 ( .A(\ab[12][43] ), .B(\CARRYB[11][43] ), .CI(\SUMB[11][44] ), 
        .CO(\CARRYB[12][43] ), .S(\SUMB[12][43] ) );
  FA1A S2_11_43 ( .A(\ab[11][43] ), .B(\CARRYB[10][43] ), .CI(\SUMB[10][44] ), 
        .CO(\CARRYB[11][43] ), .S(\SUMB[11][43] ) );
  FA1A S2_10_43 ( .A(\ab[10][43] ), .B(\CARRYB[9][43] ), .CI(\SUMB[9][44] ), 
        .CO(\CARRYB[10][43] ), .S(\SUMB[10][43] ) );
  FA1A S2_9_43 ( .A(\ab[9][43] ), .B(\CARRYB[8][43] ), .CI(\SUMB[8][44] ), 
        .CO(\CARRYB[9][43] ), .S(\SUMB[9][43] ) );
  FA1A S2_8_43 ( .A(\ab[8][43] ), .B(\CARRYB[7][43] ), .CI(\SUMB[7][44] ), 
        .CO(\CARRYB[8][43] ), .S(\SUMB[8][43] ) );
  FA1A S2_7_43 ( .A(\ab[7][43] ), .B(\CARRYB[6][43] ), .CI(\SUMB[6][44] ), 
        .CO(\CARRYB[7][43] ), .S(\SUMB[7][43] ) );
  FA1A S2_6_43 ( .A(\ab[6][43] ), .B(\CARRYB[5][43] ), .CI(\SUMB[5][44] ), 
        .CO(\CARRYB[6][43] ), .S(\SUMB[6][43] ) );
  FA1A S2_5_43 ( .A(\ab[5][43] ), .B(\CARRYB[4][43] ), .CI(\SUMB[4][44] ), 
        .CO(\CARRYB[5][43] ), .S(\SUMB[5][43] ) );
  FA1A S2_4_43 ( .A(\ab[4][43] ), .B(\CARRYB[3][43] ), .CI(\SUMB[3][44] ), 
        .CO(\CARRYB[4][43] ), .S(\SUMB[4][43] ) );
  FA1A S2_3_43 ( .A(\ab[3][43] ), .B(\CARRYB[2][43] ), .CI(\SUMB[2][44] ), 
        .CO(\CARRYB[3][43] ), .S(\SUMB[3][43] ) );
  FA1A S2_2_43 ( .A(\ab[2][43] ), .B(\CARRYB[1][43] ), .CI(\SUMB[1][44] ), 
        .CO(\CARRYB[2][43] ), .S(\SUMB[2][43] ) );
  FA1A S4_43 ( .A(\ab[21][43] ), .B(\CARRYB[20][43] ), .CI(\SUMB[20][44] ), 
        .CO(\CARRYB[21][43] ), .S(\SUMB[21][43] ) );
  FA1A S4_42 ( .A(\ab[21][42] ), .B(\CARRYB[20][42] ), .CI(\SUMB[20][43] ), 
        .CO(\CARRYB[21][42] ), .S(\SUMB[21][42] ) );
  FA1A S2_20_42 ( .A(\ab[20][42] ), .B(\CARRYB[19][42] ), .CI(\SUMB[19][43] ), 
        .CO(\CARRYB[20][42] ), .S(\SUMB[20][42] ) );
  FA1A S2_19_42 ( .A(\ab[19][42] ), .B(\CARRYB[18][42] ), .CI(\SUMB[18][43] ), 
        .CO(\CARRYB[19][42] ), .S(\SUMB[19][42] ) );
  FA1A S2_18_42 ( .A(\ab[18][42] ), .B(\CARRYB[17][42] ), .CI(\SUMB[17][43] ), 
        .CO(\CARRYB[18][42] ), .S(\SUMB[18][42] ) );
  FA1A S2_17_42 ( .A(\ab[17][42] ), .B(\CARRYB[16][42] ), .CI(\SUMB[16][43] ), 
        .CO(\CARRYB[17][42] ), .S(\SUMB[17][42] ) );
  FA1A S2_16_42 ( .A(\ab[16][42] ), .B(\CARRYB[15][42] ), .CI(\SUMB[15][43] ), 
        .CO(\CARRYB[16][42] ), .S(\SUMB[16][42] ) );
  FA1A S2_15_42 ( .A(\ab[15][42] ), .B(\CARRYB[14][42] ), .CI(\SUMB[14][43] ), 
        .CO(\CARRYB[15][42] ), .S(\SUMB[15][42] ) );
  FA1A S2_14_42 ( .A(\ab[14][42] ), .B(\CARRYB[13][42] ), .CI(\SUMB[13][43] ), 
        .CO(\CARRYB[14][42] ), .S(\SUMB[14][42] ) );
  FA1A S2_13_42 ( .A(\ab[13][42] ), .B(\CARRYB[12][42] ), .CI(\SUMB[12][43] ), 
        .CO(\CARRYB[13][42] ), .S(\SUMB[13][42] ) );
  FA1A S2_12_42 ( .A(\ab[12][42] ), .B(\CARRYB[11][42] ), .CI(\SUMB[11][43] ), 
        .CO(\CARRYB[12][42] ), .S(\SUMB[12][42] ) );
  FA1A S2_11_42 ( .A(\ab[11][42] ), .B(\CARRYB[10][42] ), .CI(\SUMB[10][43] ), 
        .CO(\CARRYB[11][42] ), .S(\SUMB[11][42] ) );
  FA1A S2_10_42 ( .A(\ab[10][42] ), .B(\CARRYB[9][42] ), .CI(\SUMB[9][43] ), 
        .CO(\CARRYB[10][42] ), .S(\SUMB[10][42] ) );
  FA1A S2_9_42 ( .A(\ab[9][42] ), .B(\CARRYB[8][42] ), .CI(\SUMB[8][43] ), 
        .CO(\CARRYB[9][42] ), .S(\SUMB[9][42] ) );
  FA1A S2_8_42 ( .A(\ab[8][42] ), .B(\CARRYB[7][42] ), .CI(\SUMB[7][43] ), 
        .CO(\CARRYB[8][42] ), .S(\SUMB[8][42] ) );
  FA1A S2_7_42 ( .A(\ab[7][42] ), .B(\CARRYB[6][42] ), .CI(\SUMB[6][43] ), 
        .CO(\CARRYB[7][42] ), .S(\SUMB[7][42] ) );
  FA1A S2_6_42 ( .A(\ab[6][42] ), .B(\CARRYB[5][42] ), .CI(\SUMB[5][43] ), 
        .CO(\CARRYB[6][42] ), .S(\SUMB[6][42] ) );
  FA1A S2_5_42 ( .A(\ab[5][42] ), .B(\CARRYB[4][42] ), .CI(\SUMB[4][43] ), 
        .CO(\CARRYB[5][42] ), .S(\SUMB[5][42] ) );
  FA1A S2_4_42 ( .A(\ab[4][42] ), .B(\CARRYB[3][42] ), .CI(\SUMB[3][43] ), 
        .CO(\CARRYB[4][42] ), .S(\SUMB[4][42] ) );
  FA1A S2_3_42 ( .A(\ab[3][42] ), .B(\CARRYB[2][42] ), .CI(\SUMB[2][43] ), 
        .CO(\CARRYB[3][42] ), .S(\SUMB[3][42] ) );
  FA1A S2_2_42 ( .A(\ab[2][42] ), .B(\CARRYB[1][42] ), .CI(\SUMB[1][43] ), 
        .CO(\CARRYB[2][42] ), .S(\SUMB[2][42] ) );
  FA1A S2_20_41 ( .A(\ab[20][41] ), .B(\CARRYB[19][41] ), .CI(\SUMB[19][42] ), 
        .CO(\CARRYB[20][41] ), .S(\SUMB[20][41] ) );
  FA1A S2_19_41 ( .A(\ab[19][41] ), .B(\CARRYB[18][41] ), .CI(\SUMB[18][42] ), 
        .CO(\CARRYB[19][41] ), .S(\SUMB[19][41] ) );
  FA1A S2_18_41 ( .A(\ab[18][41] ), .B(\CARRYB[17][41] ), .CI(\SUMB[17][42] ), 
        .CO(\CARRYB[18][41] ), .S(\SUMB[18][41] ) );
  FA1A S2_17_41 ( .A(\ab[17][41] ), .B(\CARRYB[16][41] ), .CI(\SUMB[16][42] ), 
        .CO(\CARRYB[17][41] ), .S(\SUMB[17][41] ) );
  FA1A S2_16_41 ( .A(\ab[16][41] ), .B(\CARRYB[15][41] ), .CI(\SUMB[15][42] ), 
        .CO(\CARRYB[16][41] ), .S(\SUMB[16][41] ) );
  FA1A S2_15_41 ( .A(\ab[15][41] ), .B(\CARRYB[14][41] ), .CI(\SUMB[14][42] ), 
        .CO(\CARRYB[15][41] ), .S(\SUMB[15][41] ) );
  FA1A S2_14_41 ( .A(\ab[14][41] ), .B(\CARRYB[13][41] ), .CI(\SUMB[13][42] ), 
        .CO(\CARRYB[14][41] ), .S(\SUMB[14][41] ) );
  FA1A S2_13_41 ( .A(\ab[13][41] ), .B(\CARRYB[12][41] ), .CI(\SUMB[12][42] ), 
        .CO(\CARRYB[13][41] ), .S(\SUMB[13][41] ) );
  FA1A S2_12_41 ( .A(\ab[12][41] ), .B(\CARRYB[11][41] ), .CI(\SUMB[11][42] ), 
        .CO(\CARRYB[12][41] ), .S(\SUMB[12][41] ) );
  FA1A S2_11_41 ( .A(\ab[11][41] ), .B(\CARRYB[10][41] ), .CI(\SUMB[10][42] ), 
        .CO(\CARRYB[11][41] ), .S(\SUMB[11][41] ) );
  FA1A S2_10_41 ( .A(\ab[10][41] ), .B(\CARRYB[9][41] ), .CI(\SUMB[9][42] ), 
        .CO(\CARRYB[10][41] ), .S(\SUMB[10][41] ) );
  FA1A S2_9_41 ( .A(\ab[9][41] ), .B(\CARRYB[8][41] ), .CI(\SUMB[8][42] ), 
        .CO(\CARRYB[9][41] ), .S(\SUMB[9][41] ) );
  FA1A S2_8_41 ( .A(\ab[8][41] ), .B(\CARRYB[7][41] ), .CI(\SUMB[7][42] ), 
        .CO(\CARRYB[8][41] ), .S(\SUMB[8][41] ) );
  FA1A S2_7_41 ( .A(\ab[7][41] ), .B(\CARRYB[6][41] ), .CI(\SUMB[6][42] ), 
        .CO(\CARRYB[7][41] ), .S(\SUMB[7][41] ) );
  FA1A S2_6_41 ( .A(\ab[6][41] ), .B(\CARRYB[5][41] ), .CI(\SUMB[5][42] ), 
        .CO(\CARRYB[6][41] ), .S(\SUMB[6][41] ) );
  FA1A S2_5_41 ( .A(\ab[5][41] ), .B(\CARRYB[4][41] ), .CI(\SUMB[4][42] ), 
        .CO(\CARRYB[5][41] ), .S(\SUMB[5][41] ) );
  FA1A S2_4_41 ( .A(\ab[4][41] ), .B(\CARRYB[3][41] ), .CI(\SUMB[3][42] ), 
        .CO(\CARRYB[4][41] ), .S(\SUMB[4][41] ) );
  FA1A S2_3_41 ( .A(\ab[3][41] ), .B(\CARRYB[2][41] ), .CI(\SUMB[2][42] ), 
        .CO(\CARRYB[3][41] ), .S(\SUMB[3][41] ) );
  FA1A S4_41 ( .A(\ab[21][41] ), .B(\CARRYB[20][41] ), .CI(\SUMB[20][42] ), 
        .CO(\CARRYB[21][41] ), .S(\SUMB[21][41] ) );
  FA1A S2_20_40 ( .A(\ab[20][40] ), .B(\CARRYB[19][40] ), .CI(\SUMB[19][41] ), 
        .CO(\CARRYB[20][40] ), .S(\SUMB[20][40] ) );
  FA1A S2_19_40 ( .A(\ab[19][40] ), .B(\CARRYB[18][40] ), .CI(\SUMB[18][41] ), 
        .CO(\CARRYB[19][40] ), .S(\SUMB[19][40] ) );
  FA1A S2_18_40 ( .A(\ab[18][40] ), .B(\CARRYB[17][40] ), .CI(\SUMB[17][41] ), 
        .CO(\CARRYB[18][40] ), .S(\SUMB[18][40] ) );
  FA1A S2_17_40 ( .A(\ab[17][40] ), .B(\CARRYB[16][40] ), .CI(\SUMB[16][41] ), 
        .CO(\CARRYB[17][40] ), .S(\SUMB[17][40] ) );
  FA1A S2_16_40 ( .A(\ab[16][40] ), .B(\CARRYB[15][40] ), .CI(\SUMB[15][41] ), 
        .CO(\CARRYB[16][40] ), .S(\SUMB[16][40] ) );
  FA1A S2_15_40 ( .A(\ab[15][40] ), .B(\CARRYB[14][40] ), .CI(\SUMB[14][41] ), 
        .CO(\CARRYB[15][40] ), .S(\SUMB[15][40] ) );
  FA1A S2_14_40 ( .A(\ab[14][40] ), .B(\CARRYB[13][40] ), .CI(\SUMB[13][41] ), 
        .CO(\CARRYB[14][40] ), .S(\SUMB[14][40] ) );
  FA1A S2_13_40 ( .A(\ab[13][40] ), .B(\CARRYB[12][40] ), .CI(\SUMB[12][41] ), 
        .CO(\CARRYB[13][40] ), .S(\SUMB[13][40] ) );
  FA1A S2_12_40 ( .A(\ab[12][40] ), .B(\CARRYB[11][40] ), .CI(\SUMB[11][41] ), 
        .CO(\CARRYB[12][40] ), .S(\SUMB[12][40] ) );
  FA1A S2_11_40 ( .A(\ab[11][40] ), .B(\CARRYB[10][40] ), .CI(\SUMB[10][41] ), 
        .CO(\CARRYB[11][40] ), .S(\SUMB[11][40] ) );
  FA1A S2_10_40 ( .A(\ab[10][40] ), .B(\CARRYB[9][40] ), .CI(\SUMB[9][41] ), 
        .CO(\CARRYB[10][40] ), .S(\SUMB[10][40] ) );
  FA1A S2_9_40 ( .A(\ab[9][40] ), .B(\CARRYB[8][40] ), .CI(\SUMB[8][41] ), 
        .CO(\CARRYB[9][40] ), .S(\SUMB[9][40] ) );
  FA1A S2_8_40 ( .A(\ab[8][40] ), .B(\CARRYB[7][40] ), .CI(\SUMB[7][41] ), 
        .CO(\CARRYB[8][40] ), .S(\SUMB[8][40] ) );
  FA1A S2_7_40 ( .A(\ab[7][40] ), .B(\CARRYB[6][40] ), .CI(\SUMB[6][41] ), 
        .CO(\CARRYB[7][40] ), .S(\SUMB[7][40] ) );
  FA1A S2_6_40 ( .A(\ab[6][40] ), .B(\CARRYB[5][40] ), .CI(\SUMB[5][41] ), 
        .CO(\CARRYB[6][40] ), .S(\SUMB[6][40] ) );
  FA1A S2_5_40 ( .A(\ab[5][40] ), .B(\CARRYB[4][40] ), .CI(\SUMB[4][41] ), 
        .CO(\CARRYB[5][40] ), .S(\SUMB[5][40] ) );
  FA1A S2_4_40 ( .A(\ab[4][40] ), .B(\CARRYB[3][40] ), .CI(\SUMB[3][41] ), 
        .CO(\CARRYB[4][40] ), .S(\SUMB[4][40] ) );
  FA1A S2_2_41 ( .A(\ab[2][41] ), .B(\CARRYB[1][41] ), .CI(\SUMB[1][42] ), 
        .CO(\CARRYB[2][41] ), .S(\SUMB[2][41] ) );
  FA1A S4_40 ( .A(\ab[21][40] ), .B(\CARRYB[20][40] ), .CI(\SUMB[20][41] ), 
        .CO(\CARRYB[21][40] ), .S(\SUMB[21][40] ) );
  FA1A S2_20_39 ( .A(\ab[20][39] ), .B(\CARRYB[19][39] ), .CI(\SUMB[19][40] ), 
        .CO(\CARRYB[20][39] ), .S(\SUMB[20][39] ) );
  FA1A S2_19_39 ( .A(\ab[19][39] ), .B(\CARRYB[18][39] ), .CI(\SUMB[18][40] ), 
        .CO(\CARRYB[19][39] ), .S(\SUMB[19][39] ) );
  FA1A S2_18_39 ( .A(\ab[18][39] ), .B(\CARRYB[17][39] ), .CI(\SUMB[17][40] ), 
        .CO(\CARRYB[18][39] ), .S(\SUMB[18][39] ) );
  FA1A S2_17_39 ( .A(\ab[17][39] ), .B(\CARRYB[16][39] ), .CI(\SUMB[16][40] ), 
        .CO(\CARRYB[17][39] ), .S(\SUMB[17][39] ) );
  FA1A S2_16_39 ( .A(\ab[16][39] ), .B(\CARRYB[15][39] ), .CI(\SUMB[15][40] ), 
        .CO(\CARRYB[16][39] ), .S(\SUMB[16][39] ) );
  FA1A S2_15_39 ( .A(\ab[15][39] ), .B(\CARRYB[14][39] ), .CI(\SUMB[14][40] ), 
        .CO(\CARRYB[15][39] ), .S(\SUMB[15][39] ) );
  FA1A S2_14_39 ( .A(\ab[14][39] ), .B(\CARRYB[13][39] ), .CI(\SUMB[13][40] ), 
        .CO(\CARRYB[14][39] ), .S(\SUMB[14][39] ) );
  FA1A S2_13_39 ( .A(\ab[13][39] ), .B(\CARRYB[12][39] ), .CI(\SUMB[12][40] ), 
        .CO(\CARRYB[13][39] ), .S(\SUMB[13][39] ) );
  FA1A S2_12_39 ( .A(\ab[12][39] ), .B(\CARRYB[11][39] ), .CI(\SUMB[11][40] ), 
        .CO(\CARRYB[12][39] ), .S(\SUMB[12][39] ) );
  FA1A S2_11_39 ( .A(\ab[11][39] ), .B(\CARRYB[10][39] ), .CI(\SUMB[10][40] ), 
        .CO(\CARRYB[11][39] ), .S(\SUMB[11][39] ) );
  FA1A S2_10_39 ( .A(\ab[10][39] ), .B(\CARRYB[9][39] ), .CI(\SUMB[9][40] ), 
        .CO(\CARRYB[10][39] ), .S(\SUMB[10][39] ) );
  FA1A S2_9_39 ( .A(\ab[9][39] ), .B(\CARRYB[8][39] ), .CI(\SUMB[8][40] ), 
        .CO(\CARRYB[9][39] ), .S(\SUMB[9][39] ) );
  FA1A S2_8_39 ( .A(\ab[8][39] ), .B(\CARRYB[7][39] ), .CI(\SUMB[7][40] ), 
        .CO(\CARRYB[8][39] ), .S(\SUMB[8][39] ) );
  FA1A S2_7_39 ( .A(\ab[7][39] ), .B(\CARRYB[6][39] ), .CI(\SUMB[6][40] ), 
        .CO(\CARRYB[7][39] ), .S(\SUMB[7][39] ) );
  FA1A S2_6_39 ( .A(\ab[6][39] ), .B(\CARRYB[5][39] ), .CI(\SUMB[5][40] ), 
        .CO(\CARRYB[6][39] ), .S(\SUMB[6][39] ) );
  FA1A S2_5_39 ( .A(\ab[5][39] ), .B(\CARRYB[4][39] ), .CI(\SUMB[4][40] ), 
        .CO(\CARRYB[5][39] ), .S(\SUMB[5][39] ) );
  FA1A S2_4_39 ( .A(\ab[4][39] ), .B(\CARRYB[3][39] ), .CI(\SUMB[3][40] ), 
        .CO(\CARRYB[4][39] ), .S(\SUMB[4][39] ) );
  FA1A S2_3_40 ( .A(\ab[3][40] ), .B(\CARRYB[2][40] ), .CI(\SUMB[2][41] ), 
        .CO(\CARRYB[3][40] ), .S(\SUMB[3][40] ) );
  FA1A S2_3_39 ( .A(\ab[3][39] ), .B(\CARRYB[2][39] ), .CI(\SUMB[2][40] ), 
        .CO(\CARRYB[3][39] ), .S(\SUMB[3][39] ) );
  FA1A S2_2_40 ( .A(\ab[2][40] ), .B(\CARRYB[1][40] ), .CI(\SUMB[1][41] ), 
        .CO(\CARRYB[2][40] ), .S(\SUMB[2][40] ) );
  FA1A S2_2_39 ( .A(\ab[2][39] ), .B(\CARRYB[1][39] ), .CI(\SUMB[1][40] ), 
        .CO(\CARRYB[2][39] ), .S(\SUMB[2][39] ) );
  FA1A S4_39 ( .A(\ab[21][39] ), .B(\CARRYB[20][39] ), .CI(\SUMB[20][40] ), 
        .CO(\CARRYB[21][39] ), .S(\SUMB[21][39] ) );
  FA1A S4_36 ( .A(\ab[21][36] ), .B(\CARRYB[20][36] ), .CI(\SUMB[20][37] ), 
        .CO(\CARRYB[21][36] ), .S(\SUMB[21][36] ) );
  FA1A S2_20_36 ( .A(\ab[20][36] ), .B(\CARRYB[19][36] ), .CI(\SUMB[19][37] ), 
        .CO(\CARRYB[20][36] ), .S(\SUMB[20][36] ) );
  FA1A S2_19_36 ( .A(\ab[19][36] ), .B(\CARRYB[18][36] ), .CI(\SUMB[18][37] ), 
        .CO(\CARRYB[19][36] ), .S(\SUMB[19][36] ) );
  FA1A S4_37 ( .A(\ab[21][37] ), .B(\CARRYB[20][37] ), .CI(\SUMB[20][38] ), 
        .CO(\CARRYB[21][37] ), .S(\SUMB[21][37] ) );
  FA1A S2_18_36 ( .A(\ab[18][36] ), .B(\CARRYB[17][36] ), .CI(\SUMB[17][37] ), 
        .CO(\CARRYB[18][36] ), .S(\SUMB[18][36] ) );
  FA1A S2_20_38 ( .A(\ab[20][38] ), .B(\CARRYB[19][38] ), .CI(\SUMB[19][39] ), 
        .CO(\CARRYB[20][38] ), .S(\SUMB[20][38] ) );
  FA1A S2_20_37 ( .A(\ab[20][37] ), .B(\CARRYB[19][37] ), .CI(\SUMB[19][38] ), 
        .CO(\CARRYB[20][37] ), .S(\SUMB[20][37] ) );
  FA1A S2_17_36 ( .A(\ab[17][36] ), .B(\CARRYB[16][36] ), .CI(\SUMB[16][37] ), 
        .CO(\CARRYB[17][36] ), .S(\SUMB[17][36] ) );
  FA1A S2_19_38 ( .A(\ab[19][38] ), .B(\CARRYB[18][38] ), .CI(\SUMB[18][39] ), 
        .CO(\CARRYB[19][38] ), .S(\SUMB[19][38] ) );
  FA1A S2_19_37 ( .A(\ab[19][37] ), .B(\CARRYB[18][37] ), .CI(\SUMB[18][38] ), 
        .CO(\CARRYB[19][37] ), .S(\SUMB[19][37] ) );
  FA1A S2_18_38 ( .A(\ab[18][38] ), .B(\CARRYB[17][38] ), .CI(\SUMB[17][39] ), 
        .CO(\CARRYB[18][38] ), .S(\SUMB[18][38] ) );
  FA1A S2_18_37 ( .A(\ab[18][37] ), .B(\CARRYB[17][37] ), .CI(\SUMB[17][38] ), 
        .CO(\CARRYB[18][37] ), .S(\SUMB[18][37] ) );
  FA1A S2_17_38 ( .A(\ab[17][38] ), .B(\CARRYB[16][38] ), .CI(\SUMB[16][39] ), 
        .CO(\CARRYB[17][38] ), .S(\SUMB[17][38] ) );
  FA1A S2_17_37 ( .A(\ab[17][37] ), .B(\CARRYB[16][37] ), .CI(\SUMB[16][38] ), 
        .CO(\CARRYB[17][37] ), .S(\SUMB[17][37] ) );
  FA1A S2_16_38 ( .A(\ab[16][38] ), .B(\CARRYB[15][38] ), .CI(\SUMB[15][39] ), 
        .CO(\CARRYB[16][38] ), .S(\SUMB[16][38] ) );
  FA1A S2_16_37 ( .A(\ab[16][37] ), .B(\CARRYB[15][37] ), .CI(\SUMB[15][38] ), 
        .CO(\CARRYB[16][37] ), .S(\SUMB[16][37] ) );
  FA1A S2_16_36 ( .A(\ab[16][36] ), .B(\CARRYB[15][36] ), .CI(\SUMB[15][37] ), 
        .CO(\CARRYB[16][36] ), .S(\SUMB[16][36] ) );
  FA1A S2_15_38 ( .A(\ab[15][38] ), .B(\CARRYB[14][38] ), .CI(\SUMB[14][39] ), 
        .CO(\CARRYB[15][38] ), .S(\SUMB[15][38] ) );
  FA1A S2_15_37 ( .A(\ab[15][37] ), .B(\CARRYB[14][37] ), .CI(\SUMB[14][38] ), 
        .CO(\CARRYB[15][37] ), .S(\SUMB[15][37] ) );
  FA1A S2_15_36 ( .A(\ab[15][36] ), .B(\CARRYB[14][36] ), .CI(\SUMB[14][37] ), 
        .CO(\CARRYB[15][36] ), .S(\SUMB[15][36] ) );
  FA1A S2_14_38 ( .A(\ab[14][38] ), .B(\CARRYB[13][38] ), .CI(\SUMB[13][39] ), 
        .CO(\CARRYB[14][38] ), .S(\SUMB[14][38] ) );
  FA1A S2_14_37 ( .A(\ab[14][37] ), .B(\CARRYB[13][37] ), .CI(\SUMB[13][38] ), 
        .CO(\CARRYB[14][37] ), .S(\SUMB[14][37] ) );
  FA1A S2_14_36 ( .A(\ab[14][36] ), .B(\CARRYB[13][36] ), .CI(\SUMB[13][37] ), 
        .CO(\CARRYB[14][36] ), .S(\SUMB[14][36] ) );
  FA1A S2_13_38 ( .A(\ab[13][38] ), .B(\CARRYB[12][38] ), .CI(\SUMB[12][39] ), 
        .CO(\CARRYB[13][38] ), .S(\SUMB[13][38] ) );
  FA1A S2_13_37 ( .A(\ab[13][37] ), .B(\CARRYB[12][37] ), .CI(\SUMB[12][38] ), 
        .CO(\CARRYB[13][37] ), .S(\SUMB[13][37] ) );
  FA1A S2_12_38 ( .A(\ab[12][38] ), .B(\CARRYB[11][38] ), .CI(\SUMB[11][39] ), 
        .CO(\CARRYB[12][38] ), .S(\SUMB[12][38] ) );
  FA1A S2_13_36 ( .A(\ab[13][36] ), .B(\CARRYB[12][36] ), .CI(\SUMB[12][37] ), 
        .CO(\CARRYB[13][36] ), .S(\SUMB[13][36] ) );
  FA1A S2_12_37 ( .A(\ab[12][37] ), .B(\CARRYB[11][37] ), .CI(\SUMB[11][38] ), 
        .CO(\CARRYB[12][37] ), .S(\SUMB[12][37] ) );
  FA1A S2_12_36 ( .A(\ab[12][36] ), .B(\CARRYB[11][36] ), .CI(\SUMB[11][37] ), 
        .CO(\CARRYB[12][36] ), .S(\SUMB[12][36] ) );
  FA1A S2_11_38 ( .A(\ab[11][38] ), .B(\CARRYB[10][38] ), .CI(\SUMB[10][39] ), 
        .CO(\CARRYB[11][38] ), .S(\SUMB[11][38] ) );
  FA1A S2_11_37 ( .A(\ab[11][37] ), .B(\CARRYB[10][37] ), .CI(\SUMB[10][38] ), 
        .CO(\CARRYB[11][37] ), .S(\SUMB[11][37] ) );
  FA1A S2_11_36 ( .A(\ab[11][36] ), .B(\CARRYB[10][36] ), .CI(\SUMB[10][37] ), 
        .CO(\CARRYB[11][36] ), .S(\SUMB[11][36] ) );
  FA1A S2_10_38 ( .A(\ab[10][38] ), .B(\CARRYB[9][38] ), .CI(\SUMB[9][39] ), 
        .CO(\CARRYB[10][38] ), .S(\SUMB[10][38] ) );
  FA1A S2_10_37 ( .A(\ab[10][37] ), .B(\CARRYB[9][37] ), .CI(\SUMB[9][38] ), 
        .CO(\CARRYB[10][37] ), .S(\SUMB[10][37] ) );
  FA1A S2_10_36 ( .A(\ab[10][36] ), .B(\CARRYB[9][36] ), .CI(\SUMB[9][37] ), 
        .CO(\CARRYB[10][36] ), .S(\SUMB[10][36] ) );
  FA1A S2_9_38 ( .A(\ab[9][38] ), .B(\CARRYB[8][38] ), .CI(\SUMB[8][39] ), 
        .CO(\CARRYB[9][38] ), .S(\SUMB[9][38] ) );
  FA1A S2_9_37 ( .A(\ab[9][37] ), .B(\CARRYB[8][37] ), .CI(\SUMB[8][38] ), 
        .CO(\CARRYB[9][37] ), .S(\SUMB[9][37] ) );
  FA1A S2_9_36 ( .A(\ab[9][36] ), .B(\CARRYB[8][36] ), .CI(\SUMB[8][37] ), 
        .CO(\CARRYB[9][36] ), .S(\SUMB[9][36] ) );
  FA1A S2_8_38 ( .A(\ab[8][38] ), .B(\CARRYB[7][38] ), .CI(\SUMB[7][39] ), 
        .CO(\CARRYB[8][38] ), .S(\SUMB[8][38] ) );
  FA1A S2_8_37 ( .A(\ab[8][37] ), .B(\CARRYB[7][37] ), .CI(\SUMB[7][38] ), 
        .CO(\CARRYB[8][37] ), .S(\SUMB[8][37] ) );
  FA1A S2_8_36 ( .A(\ab[8][36] ), .B(\CARRYB[7][36] ), .CI(\SUMB[7][37] ), 
        .CO(\CARRYB[8][36] ), .S(\SUMB[8][36] ) );
  FA1A S2_7_38 ( .A(\ab[7][38] ), .B(\CARRYB[6][38] ), .CI(\SUMB[6][39] ), 
        .CO(\CARRYB[7][38] ), .S(\SUMB[7][38] ) );
  FA1A S2_7_37 ( .A(\ab[7][37] ), .B(\CARRYB[6][37] ), .CI(\SUMB[6][38] ), 
        .CO(\CARRYB[7][37] ), .S(\SUMB[7][37] ) );
  FA1A S2_7_36 ( .A(\ab[7][36] ), .B(\CARRYB[6][36] ), .CI(\SUMB[6][37] ), 
        .CO(\CARRYB[7][36] ), .S(\SUMB[7][36] ) );
  FA1A S2_6_38 ( .A(\ab[6][38] ), .B(\CARRYB[5][38] ), .CI(\SUMB[5][39] ), 
        .CO(\CARRYB[6][38] ), .S(\SUMB[6][38] ) );
  FA1A S2_6_37 ( .A(\ab[6][37] ), .B(\CARRYB[5][37] ), .CI(\SUMB[5][38] ), 
        .CO(\CARRYB[6][37] ), .S(\SUMB[6][37] ) );
  FA1A S2_6_36 ( .A(\ab[6][36] ), .B(\CARRYB[5][36] ), .CI(\SUMB[5][37] ), 
        .CO(\CARRYB[6][36] ), .S(\SUMB[6][36] ) );
  FA1A S2_5_38 ( .A(\ab[5][38] ), .B(\CARRYB[4][38] ), .CI(\SUMB[4][39] ), 
        .CO(\CARRYB[5][38] ), .S(\SUMB[5][38] ) );
  FA1A S2_5_37 ( .A(\ab[5][37] ), .B(\CARRYB[4][37] ), .CI(\SUMB[4][38] ), 
        .CO(\CARRYB[5][37] ), .S(\SUMB[5][37] ) );
  FA1A S2_5_36 ( .A(\ab[5][36] ), .B(\CARRYB[4][36] ), .CI(\SUMB[4][37] ), 
        .CO(\CARRYB[5][36] ), .S(\SUMB[5][36] ) );
  FA1A S2_4_38 ( .A(\ab[4][38] ), .B(\CARRYB[3][38] ), .CI(\SUMB[3][39] ), 
        .CO(\CARRYB[4][38] ), .S(\SUMB[4][38] ) );
  FA1A S2_4_37 ( .A(\ab[4][37] ), .B(\CARRYB[3][37] ), .CI(\SUMB[3][38] ), 
        .CO(\CARRYB[4][37] ), .S(\SUMB[4][37] ) );
  FA1A S2_4_36 ( .A(\ab[4][36] ), .B(\CARRYB[3][36] ), .CI(\SUMB[3][37] ), 
        .CO(\CARRYB[4][36] ), .S(\SUMB[4][36] ) );
  FA1A S2_3_38 ( .A(\ab[3][38] ), .B(\CARRYB[2][38] ), .CI(\SUMB[2][39] ), 
        .CO(\CARRYB[3][38] ), .S(\SUMB[3][38] ) );
  FA1A S2_3_37 ( .A(\ab[3][37] ), .B(\CARRYB[2][37] ), .CI(\SUMB[2][38] ), 
        .CO(\CARRYB[3][37] ), .S(\SUMB[3][37] ) );
  FA1A S2_3_36 ( .A(\ab[3][36] ), .B(\CARRYB[2][36] ), .CI(\SUMB[2][37] ), 
        .CO(\CARRYB[3][36] ), .S(\SUMB[3][36] ) );
  FA1A S2_2_38 ( .A(\ab[2][38] ), .B(\CARRYB[1][38] ), .CI(\SUMB[1][39] ), 
        .CO(\CARRYB[2][38] ), .S(\SUMB[2][38] ) );
  FA1A S2_2_37 ( .A(\ab[2][37] ), .B(\CARRYB[1][37] ), .CI(\SUMB[1][38] ), 
        .CO(\CARRYB[2][37] ), .S(\SUMB[2][37] ) );
  FA1A S2_2_36 ( .A(\ab[2][36] ), .B(\CARRYB[1][36] ), .CI(\SUMB[1][37] ), 
        .CO(\CARRYB[2][36] ), .S(\SUMB[2][36] ) );
  FA1A S4_38 ( .A(\ab[21][38] ), .B(\CARRYB[20][38] ), .CI(\SUMB[20][39] ), 
        .CO(\CARRYB[21][38] ), .S(\SUMB[21][38] ) );
  FA1A S4_33 ( .A(\ab[21][33] ), .B(\CARRYB[20][33] ), .CI(\SUMB[20][34] ), 
        .CO(\CARRYB[21][33] ), .S(\SUMB[21][33] ) );
  FA1A S4_32 ( .A(\ab[21][32] ), .B(\CARRYB[20][32] ), .CI(\SUMB[20][33] ), 
        .CO(\CARRYB[21][32] ), .S(\SUMB[21][32] ) );
  FA1A S2_20_34 ( .A(\ab[20][34] ), .B(\CARRYB[19][34] ), .CI(\SUMB[19][35] ), 
        .CO(\CARRYB[20][34] ), .S(\SUMB[20][34] ) );
  FA1A S2_20_33 ( .A(\ab[20][33] ), .B(\CARRYB[19][33] ), .CI(\SUMB[19][34] ), 
        .CO(\CARRYB[20][33] ), .S(\SUMB[20][33] ) );
  FA1A S2_19_34 ( .A(\ab[19][34] ), .B(\CARRYB[18][34] ), .CI(\SUMB[18][35] ), 
        .CO(\CARRYB[19][34] ), .S(\SUMB[19][34] ) );
  FA1A S2_20_35 ( .A(\ab[20][35] ), .B(\CARRYB[19][35] ), .CI(\SUMB[19][36] ), 
        .CO(\CARRYB[20][35] ), .S(\SUMB[20][35] ) );
  FA1A S2_19_35 ( .A(\ab[19][35] ), .B(\CARRYB[18][35] ), .CI(\SUMB[18][36] ), 
        .CO(\CARRYB[19][35] ), .S(\SUMB[19][35] ) );
  FA1A S2_18_35 ( .A(\ab[18][35] ), .B(\CARRYB[17][35] ), .CI(\SUMB[17][36] ), 
        .CO(\CARRYB[18][35] ), .S(\SUMB[18][35] ) );
  FA1A S2_20_32 ( .A(\ab[20][32] ), .B(\CARRYB[19][32] ), .CI(\SUMB[19][33] ), 
        .CO(\CARRYB[20][32] ), .S(\SUMB[20][32] ) );
  FA1A S2_19_33 ( .A(\ab[19][33] ), .B(\CARRYB[18][33] ), .CI(\SUMB[18][34] ), 
        .CO(\CARRYB[19][33] ), .S(\SUMB[19][33] ) );
  FA1A S2_19_32 ( .A(\ab[19][32] ), .B(\CARRYB[18][32] ), .CI(\SUMB[18][33] ), 
        .CO(\CARRYB[19][32] ), .S(\SUMB[19][32] ) );
  FA1A S2_18_34 ( .A(\ab[18][34] ), .B(\CARRYB[17][34] ), .CI(\SUMB[17][35] ), 
        .CO(\CARRYB[18][34] ), .S(\SUMB[18][34] ) );
  FA1A S2_18_33 ( .A(\ab[18][33] ), .B(\CARRYB[17][33] ), .CI(\SUMB[17][34] ), 
        .CO(\CARRYB[18][33] ), .S(\SUMB[18][33] ) );
  FA1A S2_18_32 ( .A(\ab[18][32] ), .B(\CARRYB[17][32] ), .CI(\SUMB[17][33] ), 
        .CO(\CARRYB[18][32] ), .S(\SUMB[18][32] ) );
  FA1A S2_17_35 ( .A(\ab[17][35] ), .B(\CARRYB[16][35] ), .CI(\SUMB[16][36] ), 
        .CO(\CARRYB[17][35] ), .S(\SUMB[17][35] ) );
  FA1A S2_17_34 ( .A(\ab[17][34] ), .B(\CARRYB[16][34] ), .CI(\SUMB[16][35] ), 
        .CO(\CARRYB[17][34] ), .S(\SUMB[17][34] ) );
  FA1A S2_17_33 ( .A(\ab[17][33] ), .B(\CARRYB[16][33] ), .CI(\SUMB[16][34] ), 
        .CO(\CARRYB[17][33] ), .S(\SUMB[17][33] ) );
  FA1A S2_16_35 ( .A(\ab[16][35] ), .B(\CARRYB[15][35] ), .CI(\SUMB[15][36] ), 
        .CO(\CARRYB[16][35] ), .S(\SUMB[16][35] ) );
  FA1A S2_16_34 ( .A(\ab[16][34] ), .B(\CARRYB[15][34] ), .CI(\SUMB[15][35] ), 
        .CO(\CARRYB[16][34] ), .S(\SUMB[16][34] ) );
  FA1A S2_17_32 ( .A(\ab[17][32] ), .B(\CARRYB[16][32] ), .CI(\SUMB[16][33] ), 
        .CO(\CARRYB[17][32] ), .S(\SUMB[17][32] ) );
  FA1A S2_15_35 ( .A(\ab[15][35] ), .B(\CARRYB[14][35] ), .CI(\SUMB[14][36] ), 
        .CO(\CARRYB[15][35] ), .S(\SUMB[15][35] ) );
  FA1A S2_16_33 ( .A(\ab[16][33] ), .B(\CARRYB[15][33] ), .CI(\SUMB[15][34] ), 
        .CO(\CARRYB[16][33] ), .S(\SUMB[16][33] ) );
  FA1A S2_16_32 ( .A(\ab[16][32] ), .B(\CARRYB[15][32] ), .CI(\SUMB[15][33] ), 
        .CO(\CARRYB[16][32] ), .S(\SUMB[16][32] ) );
  FA1A S2_15_34 ( .A(\ab[15][34] ), .B(\CARRYB[14][34] ), .CI(\SUMB[14][35] ), 
        .CO(\CARRYB[15][34] ), .S(\SUMB[15][34] ) );
  FA1A S2_15_33 ( .A(\ab[15][33] ), .B(\CARRYB[14][33] ), .CI(\SUMB[14][34] ), 
        .CO(\CARRYB[15][33] ), .S(\SUMB[15][33] ) );
  FA1A S2_15_32 ( .A(\ab[15][32] ), .B(\CARRYB[14][32] ), .CI(\SUMB[14][33] ), 
        .CO(\CARRYB[15][32] ), .S(\SUMB[15][32] ) );
  FA1A S2_14_35 ( .A(\ab[14][35] ), .B(\CARRYB[13][35] ), .CI(\SUMB[13][36] ), 
        .CO(\CARRYB[14][35] ), .S(\SUMB[14][35] ) );
  FA1A S2_14_34 ( .A(\ab[14][34] ), .B(\CARRYB[13][34] ), .CI(\SUMB[13][35] ), 
        .CO(\CARRYB[14][34] ), .S(\SUMB[14][34] ) );
  FA1A S2_14_33 ( .A(\ab[14][33] ), .B(\CARRYB[13][33] ), .CI(\SUMB[13][34] ), 
        .CO(\CARRYB[14][33] ), .S(\SUMB[14][33] ) );
  FA1A S2_14_32 ( .A(\ab[14][32] ), .B(\CARRYB[13][32] ), .CI(\SUMB[13][33] ), 
        .CO(\CARRYB[14][32] ), .S(\SUMB[14][32] ) );
  FA1A S2_13_35 ( .A(\ab[13][35] ), .B(\CARRYB[12][35] ), .CI(\SUMB[12][36] ), 
        .CO(\CARRYB[13][35] ), .S(\SUMB[13][35] ) );
  FA1A S2_13_34 ( .A(\ab[13][34] ), .B(\CARRYB[12][34] ), .CI(\SUMB[12][35] ), 
        .CO(\CARRYB[13][34] ), .S(\SUMB[13][34] ) );
  FA1A S2_13_33 ( .A(\ab[13][33] ), .B(\CARRYB[12][33] ), .CI(\SUMB[12][34] ), 
        .CO(\CARRYB[13][33] ), .S(\SUMB[13][33] ) );
  FA1A S2_13_32 ( .A(\ab[13][32] ), .B(\CARRYB[12][32] ), .CI(\SUMB[12][33] ), 
        .CO(\CARRYB[13][32] ), .S(\SUMB[13][32] ) );
  FA1A S2_12_35 ( .A(\ab[12][35] ), .B(\CARRYB[11][35] ), .CI(\SUMB[11][36] ), 
        .CO(\CARRYB[12][35] ), .S(\SUMB[12][35] ) );
  FA1A S2_12_34 ( .A(\ab[12][34] ), .B(\CARRYB[11][34] ), .CI(\SUMB[11][35] ), 
        .CO(\CARRYB[12][34] ), .S(\SUMB[12][34] ) );
  FA1A S2_12_33 ( .A(\ab[12][33] ), .B(\CARRYB[11][33] ), .CI(\SUMB[11][34] ), 
        .CO(\CARRYB[12][33] ), .S(\SUMB[12][33] ) );
  FA1A S2_12_32 ( .A(\ab[12][32] ), .B(\CARRYB[11][32] ), .CI(\SUMB[11][33] ), 
        .CO(\CARRYB[12][32] ), .S(\SUMB[12][32] ) );
  FA1A S2_11_35 ( .A(\ab[11][35] ), .B(\CARRYB[10][35] ), .CI(\SUMB[10][36] ), 
        .CO(\CARRYB[11][35] ), .S(\SUMB[11][35] ) );
  FA1A S2_11_34 ( .A(\ab[11][34] ), .B(\CARRYB[10][34] ), .CI(\SUMB[10][35] ), 
        .CO(\CARRYB[11][34] ), .S(\SUMB[11][34] ) );
  FA1A S2_11_33 ( .A(\ab[11][33] ), .B(\CARRYB[10][33] ), .CI(\SUMB[10][34] ), 
        .CO(\CARRYB[11][33] ), .S(\SUMB[11][33] ) );
  FA1A S2_11_32 ( .A(\ab[11][32] ), .B(\CARRYB[10][32] ), .CI(\SUMB[10][33] ), 
        .CO(\CARRYB[11][32] ), .S(\SUMB[11][32] ) );
  FA1A S2_10_35 ( .A(\ab[10][35] ), .B(\CARRYB[9][35] ), .CI(\SUMB[9][36] ), 
        .CO(\CARRYB[10][35] ), .S(\SUMB[10][35] ) );
  FA1A S2_10_34 ( .A(\ab[10][34] ), .B(\CARRYB[9][34] ), .CI(\SUMB[9][35] ), 
        .CO(\CARRYB[10][34] ), .S(\SUMB[10][34] ) );
  FA1A S2_10_33 ( .A(\ab[10][33] ), .B(\CARRYB[9][33] ), .CI(\SUMB[9][34] ), 
        .CO(\CARRYB[10][33] ), .S(\SUMB[10][33] ) );
  FA1A S2_10_32 ( .A(\ab[10][32] ), .B(\CARRYB[9][32] ), .CI(\SUMB[9][33] ), 
        .CO(\CARRYB[10][32] ), .S(\SUMB[10][32] ) );
  FA1A S2_9_35 ( .A(\ab[9][35] ), .B(\CARRYB[8][35] ), .CI(\SUMB[8][36] ), 
        .CO(\CARRYB[9][35] ), .S(\SUMB[9][35] ) );
  FA1A S2_9_34 ( .A(\ab[9][34] ), .B(\CARRYB[8][34] ), .CI(\SUMB[8][35] ), 
        .CO(\CARRYB[9][34] ), .S(\SUMB[9][34] ) );
  FA1A S2_9_33 ( .A(\ab[9][33] ), .B(\CARRYB[8][33] ), .CI(\SUMB[8][34] ), 
        .CO(\CARRYB[9][33] ), .S(\SUMB[9][33] ) );
  FA1A S2_9_32 ( .A(\ab[9][32] ), .B(\CARRYB[8][32] ), .CI(\SUMB[8][33] ), 
        .CO(\CARRYB[9][32] ), .S(\SUMB[9][32] ) );
  FA1A S2_8_35 ( .A(\ab[8][35] ), .B(\CARRYB[7][35] ), .CI(\SUMB[7][36] ), 
        .CO(\CARRYB[8][35] ), .S(\SUMB[8][35] ) );
  FA1A S2_8_34 ( .A(\ab[8][34] ), .B(\CARRYB[7][34] ), .CI(\SUMB[7][35] ), 
        .CO(\CARRYB[8][34] ), .S(\SUMB[8][34] ) );
  FA1A S2_8_33 ( .A(\ab[8][33] ), .B(\CARRYB[7][33] ), .CI(\SUMB[7][34] ), 
        .CO(\CARRYB[8][33] ), .S(\SUMB[8][33] ) );
  FA1A S2_8_32 ( .A(\ab[8][32] ), .B(\CARRYB[7][32] ), .CI(\SUMB[7][33] ), 
        .CO(\CARRYB[8][32] ), .S(\SUMB[8][32] ) );
  FA1A S2_7_35 ( .A(\ab[7][35] ), .B(\CARRYB[6][35] ), .CI(\SUMB[6][36] ), 
        .CO(\CARRYB[7][35] ), .S(\SUMB[7][35] ) );
  FA1A S2_7_34 ( .A(\ab[7][34] ), .B(\CARRYB[6][34] ), .CI(\SUMB[6][35] ), 
        .CO(\CARRYB[7][34] ), .S(\SUMB[7][34] ) );
  FA1A S2_7_33 ( .A(\ab[7][33] ), .B(\CARRYB[6][33] ), .CI(\SUMB[6][34] ), 
        .CO(\CARRYB[7][33] ), .S(\SUMB[7][33] ) );
  FA1A S2_7_32 ( .A(\ab[7][32] ), .B(\CARRYB[6][32] ), .CI(\SUMB[6][33] ), 
        .CO(\CARRYB[7][32] ), .S(\SUMB[7][32] ) );
  FA1A S2_6_35 ( .A(\ab[6][35] ), .B(\CARRYB[5][35] ), .CI(\SUMB[5][36] ), 
        .CO(\CARRYB[6][35] ), .S(\SUMB[6][35] ) );
  FA1A S2_6_34 ( .A(\ab[6][34] ), .B(\CARRYB[5][34] ), .CI(\SUMB[5][35] ), 
        .CO(\CARRYB[6][34] ), .S(\SUMB[6][34] ) );
  FA1A S2_6_33 ( .A(\ab[6][33] ), .B(\CARRYB[5][33] ), .CI(\SUMB[5][34] ), 
        .CO(\CARRYB[6][33] ), .S(\SUMB[6][33] ) );
  FA1A S2_6_32 ( .A(\ab[6][32] ), .B(\CARRYB[5][32] ), .CI(\SUMB[5][33] ), 
        .CO(\CARRYB[6][32] ), .S(\SUMB[6][32] ) );
  FA1A S2_5_35 ( .A(\ab[5][35] ), .B(\CARRYB[4][35] ), .CI(\SUMB[4][36] ), 
        .CO(\CARRYB[5][35] ), .S(\SUMB[5][35] ) );
  FA1A S2_5_34 ( .A(\ab[5][34] ), .B(\CARRYB[4][34] ), .CI(\SUMB[4][35] ), 
        .CO(\CARRYB[5][34] ), .S(\SUMB[5][34] ) );
  FA1A S2_5_33 ( .A(\ab[5][33] ), .B(\CARRYB[4][33] ), .CI(\SUMB[4][34] ), 
        .CO(\CARRYB[5][33] ), .S(\SUMB[5][33] ) );
  FA1A S2_5_32 ( .A(\ab[5][32] ), .B(\CARRYB[4][32] ), .CI(\SUMB[4][33] ), 
        .CO(\CARRYB[5][32] ), .S(\SUMB[5][32] ) );
  FA1A S2_4_35 ( .A(\ab[4][35] ), .B(\CARRYB[3][35] ), .CI(\SUMB[3][36] ), 
        .CO(\CARRYB[4][35] ), .S(\SUMB[4][35] ) );
  FA1A S2_4_34 ( .A(\ab[4][34] ), .B(\CARRYB[3][34] ), .CI(\SUMB[3][35] ), 
        .CO(\CARRYB[4][34] ), .S(\SUMB[4][34] ) );
  FA1A S2_4_33 ( .A(\ab[4][33] ), .B(\CARRYB[3][33] ), .CI(\SUMB[3][34] ), 
        .CO(\CARRYB[4][33] ), .S(\SUMB[4][33] ) );
  FA1A S2_4_32 ( .A(\ab[4][32] ), .B(\CARRYB[3][32] ), .CI(\SUMB[3][33] ), 
        .CO(\CARRYB[4][32] ), .S(\SUMB[4][32] ) );
  FA1A S2_3_35 ( .A(\ab[3][35] ), .B(\CARRYB[2][35] ), .CI(\SUMB[2][36] ), 
        .CO(\CARRYB[3][35] ), .S(\SUMB[3][35] ) );
  FA1A S2_3_34 ( .A(\ab[3][34] ), .B(\CARRYB[2][34] ), .CI(\SUMB[2][35] ), 
        .CO(\CARRYB[3][34] ), .S(\SUMB[3][34] ) );
  FA1A S2_3_33 ( .A(\ab[3][33] ), .B(\CARRYB[2][33] ), .CI(\SUMB[2][34] ), 
        .CO(\CARRYB[3][33] ), .S(\SUMB[3][33] ) );
  FA1A S2_3_32 ( .A(\ab[3][32] ), .B(\CARRYB[2][32] ), .CI(\SUMB[2][33] ), 
        .CO(\CARRYB[3][32] ), .S(\SUMB[3][32] ) );
  FA1A S2_2_35 ( .A(\ab[2][35] ), .B(\CARRYB[1][35] ), .CI(\SUMB[1][36] ), 
        .CO(\CARRYB[2][35] ), .S(\SUMB[2][35] ) );
  FA1A S2_2_34 ( .A(\ab[2][34] ), .B(\CARRYB[1][34] ), .CI(\SUMB[1][35] ), 
        .CO(\CARRYB[2][34] ), .S(\SUMB[2][34] ) );
  FA1A S2_2_33 ( .A(\ab[2][33] ), .B(\CARRYB[1][33] ), .CI(\SUMB[1][34] ), 
        .CO(\CARRYB[2][33] ), .S(\SUMB[2][33] ) );
  FA1A S2_2_32 ( .A(\ab[2][32] ), .B(\CARRYB[1][32] ), .CI(\SUMB[1][33] ), 
        .CO(\CARRYB[2][32] ), .S(\SUMB[2][32] ) );
  FA1A S4_34 ( .A(\ab[21][34] ), .B(\CARRYB[20][34] ), .CI(\SUMB[20][35] ), 
        .CO(\CARRYB[21][34] ), .S(\SUMB[21][34] ) );
  FA1A S4_35 ( .A(\ab[21][35] ), .B(\CARRYB[20][35] ), .CI(\SUMB[20][36] ), 
        .CO(\CARRYB[21][35] ), .S(\SUMB[21][35] ) );
  FA1A S4_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA1A S2_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\SUMB[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA1A S2_20_31 ( .A(\ab[20][31] ), .B(\CARRYB[19][31] ), .CI(\SUMB[19][32] ), 
        .CO(\CARRYB[20][31] ), .S(\SUMB[20][31] ) );
  FA1A S2_19_31 ( .A(\ab[19][31] ), .B(\CARRYB[18][31] ), .CI(\SUMB[18][32] ), 
        .CO(\CARRYB[19][31] ), .S(\SUMB[19][31] ) );
  FA1A S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA1A S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA1A S2_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\SUMB[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA1A S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA1A S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA1A S2_18_31 ( .A(\ab[18][31] ), .B(\CARRYB[17][31] ), .CI(\SUMB[17][32] ), 
        .CO(\CARRYB[18][31] ), .S(\SUMB[18][31] ) );
  FA1A S2_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\SUMB[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA1A S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA1A S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA1A S2_17_31 ( .A(\ab[17][31] ), .B(\CARRYB[16][31] ), .CI(\SUMB[16][32] ), 
        .CO(\CARRYB[17][31] ), .S(\SUMB[17][31] ) );
  FA1A S2_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\SUMB[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA1A S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA1A S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA1A S2_16_31 ( .A(\ab[16][31] ), .B(\CARRYB[15][31] ), .CI(\SUMB[15][32] ), 
        .CO(\CARRYB[16][31] ), .S(\SUMB[16][31] ) );
  FA1A S2_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\SUMB[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA1A S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA1A S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA1A S2_15_31 ( .A(\ab[15][31] ), .B(\CARRYB[14][31] ), .CI(\SUMB[14][32] ), 
        .CO(\CARRYB[15][31] ), .S(\SUMB[15][31] ) );
  FA1A S2_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\SUMB[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA1A S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA1A S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA1A S2_14_31 ( .A(\ab[14][31] ), .B(\CARRYB[13][31] ), .CI(\SUMB[13][32] ), 
        .CO(\CARRYB[14][31] ), .S(\SUMB[14][31] ) );
  FA1A S2_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\SUMB[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA1A S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA1A S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA1A S2_13_31 ( .A(\ab[13][31] ), .B(\CARRYB[12][31] ), .CI(\SUMB[12][32] ), 
        .CO(\CARRYB[13][31] ), .S(\SUMB[13][31] ) );
  FA1A S2_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\SUMB[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA1A S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA1A S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA1A S2_12_31 ( .A(\ab[12][31] ), .B(\CARRYB[11][31] ), .CI(\SUMB[11][32] ), 
        .CO(\CARRYB[12][31] ), .S(\SUMB[12][31] ) );
  FA1A S2_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\SUMB[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA1A S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA1A S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA1A S2_11_31 ( .A(\ab[11][31] ), .B(\CARRYB[10][31] ), .CI(\SUMB[10][32] ), 
        .CO(\CARRYB[11][31] ), .S(\SUMB[11][31] ) );
  FA1A S2_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\SUMB[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA1A S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1A S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1A S2_10_31 ( .A(\ab[10][31] ), .B(\CARRYB[9][31] ), .CI(\SUMB[9][32] ), 
        .CO(\CARRYB[10][31] ), .S(\SUMB[10][31] ) );
  FA1A S2_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\SUMB[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA1A S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1A S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1A S2_9_31 ( .A(\ab[9][31] ), .B(\CARRYB[8][31] ), .CI(\SUMB[8][32] ), 
        .CO(\CARRYB[9][31] ), .S(\SUMB[9][31] ) );
  FA1A S2_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\SUMB[8][31] ), 
        .CO(\CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA1A S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1A S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1A S2_8_31 ( .A(\ab[8][31] ), .B(\CARRYB[7][31] ), .CI(\SUMB[7][32] ), 
        .CO(\CARRYB[8][31] ), .S(\SUMB[8][31] ) );
  FA1A S2_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\SUMB[7][31] ), 
        .CO(\CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA1A S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1A S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA1A S2_7_31 ( .A(\ab[7][31] ), .B(\CARRYB[6][31] ), .CI(\SUMB[6][32] ), 
        .CO(\CARRYB[7][31] ), .S(\SUMB[7][31] ) );
  FA1A S2_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\SUMB[6][31] ), 
        .CO(\CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA1A S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1A S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA1A S2_6_31 ( .A(\ab[6][31] ), .B(\CARRYB[5][31] ), .CI(\SUMB[5][32] ), 
        .CO(\CARRYB[6][31] ), .S(\SUMB[6][31] ) );
  FA1A S2_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\SUMB[5][31] ), 
        .CO(\CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA1A S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA1A S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1A S2_5_31 ( .A(\ab[5][31] ), .B(\CARRYB[4][31] ), .CI(\SUMB[4][32] ), 
        .CO(\CARRYB[5][31] ), .S(\SUMB[5][31] ) );
  FA1A S2_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\SUMB[4][31] ), 
        .CO(\CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA1A S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA1A S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA1A S2_4_31 ( .A(\ab[4][31] ), .B(\CARRYB[3][31] ), .CI(\SUMB[3][32] ), 
        .CO(\CARRYB[4][31] ), .S(\SUMB[4][31] ) );
  FA1A S2_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\SUMB[3][31] ), 
        .CO(\CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA1A S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\SUMB[3][30] ), 
        .CO(\CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1A S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1A S2_3_31 ( .A(\ab[3][31] ), .B(\CARRYB[2][31] ), .CI(\SUMB[2][32] ), 
        .CO(\CARRYB[3][31] ), .S(\SUMB[3][31] ) );
  FA1A S2_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .CI(\SUMB[2][31] ), 
        .CO(\CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA1A S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1A S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA1A S2_2_31 ( .A(\ab[2][31] ), .B(\CARRYB[1][31] ), .CI(\SUMB[1][32] ), 
        .CO(\CARRYB[2][31] ), .S(\SUMB[2][31] ) );
  FA1A S2_2_30 ( .A(\ab[2][30] ), .B(\CARRYB[1][30] ), .CI(\SUMB[1][31] ), 
        .CO(\CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  FA1A S2_2_29 ( .A(\ab[2][29] ), .B(\CARRYB[1][29] ), .CI(\SUMB[1][30] ), 
        .CO(\CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1A S2_2_28 ( .A(\ab[2][28] ), .B(\CARRYB[1][28] ), .CI(\SUMB[1][29] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FA1A S4_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\SUMB[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA1A S4_31 ( .A(\ab[21][31] ), .B(\CARRYB[20][31] ), .CI(\SUMB[20][32] ), 
        .CO(\CARRYB[21][31] ), .S(\SUMB[21][31] ) );
  FA1A S4_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA1A S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA1A S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA1A S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA1A S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA1A S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA1A S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA1A S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA1A S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA1A S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA1A S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA1A S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA1A S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1A S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1A S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA1A S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA1A S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1A S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1A S2_2_27 ( .A(\ab[2][27] ), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1A S4_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA1A S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA1A S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA1A S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA1A S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA1A S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA1A S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA1A S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA1A S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA1A S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA1A S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1A S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA1A S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1A S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1A S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA1A S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA1A S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1A S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1A S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1A S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1A S4_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA1A S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA1A S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA1A S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA1A S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA1A S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA1A S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA1A S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA1A S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA1A S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA1A S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1A S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1A S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1A S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1A S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA1A S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA1A S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1A S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1A S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA1A S4_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA1A S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA1A S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA1A S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA1A S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA1A S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA1A S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA1A S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA1A S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA1A S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA1A S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1A S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1A S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1A S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1A S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA1A S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1A S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1A S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1A S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA1A S2_2_25 ( .A(\ab[2][25] ), .B(\CARRYB[1][25] ), .CI(\SUMB[1][26] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1A S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), 
        .CO(\CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA1A S4_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA1A S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA1A S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA1A S4_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA1A S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA1A S4_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA1A S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA1A S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA1A S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA1A S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA1A S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA1A S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA1A S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA1A S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA1A S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA1A S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA1A S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA1A S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA1A S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA1A S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA1A S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA1A S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA1A S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA1A S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA1A S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA1A S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA1A S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA1A S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA1A S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA1A S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA1A S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA1A S2_11_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1A S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1A S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1A S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA1A S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1A S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1A S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1A S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1A S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA1A S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1A S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1A S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA1A S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1A S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA1A S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA1A S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA1A S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1A S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1A S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA1A S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1A S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1A S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1A S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1A S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA1A S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1A S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1A S4_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA1A S4_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1A S4_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA1A S4_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA1A S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA1A S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA1A S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA1A S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA1A S4_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA1A S4_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA1A S4_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA1A S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA1A S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA1A S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA1A S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA1A S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA1A S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA1A S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA1A S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA1A S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA1A S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA1A S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA1A S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA1A S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA1A S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA1A S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA1A S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA1A S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA1A S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA1A S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA1A S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA1A S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA1A S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA1A S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA1A S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA1A S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA1A S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA1A S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA1A S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA1A S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA1A S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA1A S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA1A S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA1A S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA1A S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA1A S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA1A S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1A S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA1A S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA1A S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA1A S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA1A S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1A S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA1A S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA1A S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA1A S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1A S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1A S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA1A S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA1A S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA1A S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA1A S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA1A S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1A S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1A S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1A S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA1A S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA1A S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1A S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1A S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1A S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1A S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA1A S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA1A S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA1A S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1A S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1A S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA1A S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), 
        .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA1A S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA1A S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1A S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S4_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA1A S4_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA1A S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA1A S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA1A S4_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA1A S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA1A S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA1A S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA1A S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA1A S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA1A S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA1A S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA1A S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA1A S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA1A S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA1A S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA1A S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA1A S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA1A S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA1A S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA1A S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA1A S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA1A S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA1A S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA1A S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA1A S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA1A S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA1A S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA1A S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA1A S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA1A S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA1A S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA1A S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA1A S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA1A S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1A S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1A S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1A S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1A S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1A S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1A S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1A S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1A S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S4_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA1A S4_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA1A S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA1A S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA1A S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA1A S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S4_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), .CO(
        \CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1A S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1A S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA1A S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA1A S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA1A S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA1A S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1A S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), .CO(
        \CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1A S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1A S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1A S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), .CO(
        \CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA1A S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA1A S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1A S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1A S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1A S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA1A S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1A S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1A S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1A S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1A S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S4_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), .CO(
        \CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA1A S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1A S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1A S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1A S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S4_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), .CO(
        \CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1A S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1A S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA1A S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1A S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1A S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA1A S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA1A S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1A S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1A S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1A S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1A S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1A S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA1A S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1A S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA1A S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1A S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1A S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1A S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S4_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), .CO(
        \CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA1A S4_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), .CO(
        \CARRYB[21][0] ), .S(\SUMB[21][0] ) );
  FA1A S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA1A S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA1A S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA1A S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1A S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA1A S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1A S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1A S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1A S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1A S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1A S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1A S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1A S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1A S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1A S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), .CO(
        \CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1A S4_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), .CO(
        \CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1A S4_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), .CO(
        \CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1A S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1A S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA1A S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1A S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1A S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1A S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  IVP U2 ( .A(n40), .Z(n38) );
  IVP U3 ( .A(n40), .Z(n37) );
  IVP U4 ( .A(n40), .Z(n39) );
  IVP U5 ( .A(n40), .Z(n36) );
  IVP U6 ( .A(n112), .Z(n40) );
  IVP U7 ( .A(A[0]), .Z(n112) );
  IVP U8 ( .A(n45), .Z(n41) );
  IVP U9 ( .A(n45), .Z(n42) );
  IVP U10 ( .A(n45), .Z(n43) );
  IVP U11 ( .A(n50), .Z(n47) );
  IVP U12 ( .A(n50), .Z(n48) );
  IVP U13 ( .A(n50), .Z(n49) );
  IVP U14 ( .A(n50), .Z(n46) );
  IVP U15 ( .A(n45), .Z(n44) );
  IVP U16 ( .A(n55), .Z(n52) );
  IVP U17 ( .A(n55), .Z(n53) );
  IVP U18 ( .A(n55), .Z(n51) );
  IVP U19 ( .A(n55), .Z(n54) );
  IVP U20 ( .A(n60), .Z(n57) );
  IVP U21 ( .A(n60), .Z(n56) );
  IVP U22 ( .A(n60), .Z(n58) );
  IVP U23 ( .A(n60), .Z(n59) );
  IVP U24 ( .A(n65), .Z(n62) );
  IVP U25 ( .A(n65), .Z(n61) );
  IVP U26 ( .A(n65), .Z(n64) );
  IVP U27 ( .A(n65), .Z(n63) );
  IVP U28 ( .A(n70), .Z(n67) );
  IVP U29 ( .A(n70), .Z(n66) );
  IVP U30 ( .A(n70), .Z(n69) );
  IVP U31 ( .A(n70), .Z(n68) );
  IVP U32 ( .A(n75), .Z(n72) );
  IVP U33 ( .A(n75), .Z(n71) );
  IVP U34 ( .A(n75), .Z(n73) );
  IVP U35 ( .A(n75), .Z(n74) );
  IVP U36 ( .A(n80), .Z(n76) );
  IVP U37 ( .A(n80), .Z(n77) );
  IVP U38 ( .A(n80), .Z(n78) );
  IVP U39 ( .A(n80), .Z(n79) );
  IVP U40 ( .A(n85), .Z(n82) );
  IVP U41 ( .A(n85), .Z(n83) );
  IVP U42 ( .A(n85), .Z(n81) );
  IVP U43 ( .A(n85), .Z(n84) );
  IVP U44 ( .A(n90), .Z(n87) );
  IVP U45 ( .A(n90), .Z(n88) );
  IVP U46 ( .A(n90), .Z(n86) );
  IVP U47 ( .A(n90), .Z(n89) );
  IVP U48 ( .A(n95), .Z(n92) );
  IVP U49 ( .A(n95), .Z(n93) );
  IVP U50 ( .A(n95), .Z(n91) );
  IVP U51 ( .A(n95), .Z(n94) );
  IVP U52 ( .A(n100), .Z(n97) );
  IVP U53 ( .A(n100), .Z(n98) );
  IVP U54 ( .A(n100), .Z(n96) );
  IVP U55 ( .A(n100), .Z(n99) );
  IVP U56 ( .A(n113), .Z(n45) );
  IVP U57 ( .A(A[1]), .Z(n113) );
  IVP U58 ( .A(n114), .Z(n50) );
  IVP U59 ( .A(A[2]), .Z(n114) );
  IVP U60 ( .A(n115), .Z(n55) );
  IVP U61 ( .A(A[3]), .Z(n115) );
  IVP U62 ( .A(n116), .Z(n60) );
  IVP U63 ( .A(A[4]), .Z(n116) );
  IVP U64 ( .A(n117), .Z(n65) );
  IVP U65 ( .A(A[5]), .Z(n117) );
  IVP U66 ( .A(n118), .Z(n70) );
  IVP U67 ( .A(A[6]), .Z(n118) );
  IVP U68 ( .A(n119), .Z(n75) );
  IVP U69 ( .A(A[7]), .Z(n119) );
  IVP U70 ( .A(n120), .Z(n80) );
  IVP U71 ( .A(A[8]), .Z(n120) );
  IVP U72 ( .A(n121), .Z(n85) );
  IVP U73 ( .A(A[9]), .Z(n121) );
  IVP U74 ( .A(n122), .Z(n90) );
  IVP U75 ( .A(A[10]), .Z(n122) );
  IVP U76 ( .A(n123), .Z(n95) );
  IVP U77 ( .A(A[11]), .Z(n123) );
  IVP U78 ( .A(n124), .Z(n100) );
  IVP U79 ( .A(A[12]), .Z(n124) );
  IVP U80 ( .A(n35), .Z(n32) );
  IVP U81 ( .A(n35), .Z(n33) );
  IVP U82 ( .A(n35), .Z(n31) );
  IVP U83 ( .A(n35), .Z(n34) );
  IVP U84 ( .A(n7), .Z(n4) );
  IVP U85 ( .A(n7), .Z(n3) );
  IVP U86 ( .A(n30), .Z(n27) );
  IVP U87 ( .A(n7), .Z(n5) );
  IVP U88 ( .A(n30), .Z(n26) );
  IVP U89 ( .A(n7), .Z(n6) );
  IVP U90 ( .A(n30), .Z(n28) );
  IVP U91 ( .A(n30), .Z(n29) );
  IVP U92 ( .A(A[16]), .Z(n23) );
  IVP U93 ( .A(A[16]), .Z(n24) );
  IVP U94 ( .A(A[16]), .Z(n25) );
  IVP U95 ( .A(A[17]), .Z(n22) );
  IVP U96 ( .A(A[18]), .Z(n20) );
  IVP U97 ( .A(A[18]), .Z(n21) );
  IVP U98 ( .A(A[19]), .Z(n17) );
  IVP U99 ( .A(A[19]), .Z(n16) );
  IVP U100 ( .A(A[19]), .Z(n18) );
  IVP U101 ( .A(A[19]), .Z(n19) );
  IVP U102 ( .A(A[20]), .Z(n13) );
  IVP U103 ( .A(A[20]), .Z(n12) );
  IVP U104 ( .A(A[20]), .Z(n14) );
  IVP U105 ( .A(A[20]), .Z(n15) );
  IVP U106 ( .A(A[21]), .Z(n9) );
  IVP U107 ( .A(A[21]), .Z(n10) );
  IVP U108 ( .A(A[21]), .Z(n8) );
  IVP U109 ( .A(A[21]), .Z(n11) );
  IVP U110 ( .A(n111), .Z(n35) );
  IVP U111 ( .A(A[13]), .Z(n111) );
  IVP U112 ( .A(n109), .Z(n7) );
  IVP U113 ( .A(A[14]), .Z(n109) );
  IVP U114 ( .A(n110), .Z(n30) );
  IVP U115 ( .A(A[15]), .Z(n110) );
  EO U116 ( .A(\CARRYB[21][4] ), .B(\SUMB[21][5] ), .Z(\A1[24] ) );
  EO U117 ( .A(\CARRYB[21][9] ), .B(\SUMB[21][10] ), .Z(\A1[29] ) );
  EO U118 ( .A(\CARRYB[21][1] ), .B(\SUMB[21][2] ), .Z(\A1[21] ) );
  EO U119 ( .A(\CARRYB[21][2] ), .B(\SUMB[21][3] ), .Z(\A1[22] ) );
  EO U120 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  EO U121 ( .A(\CARRYB[21][3] ), .B(\SUMB[21][4] ), .Z(\A1[23] ) );
  EO U122 ( .A(\CARRYB[21][5] ), .B(\SUMB[21][6] ), .Z(\A1[25] ) );
  EO U123 ( .A(\CARRYB[21][6] ), .B(\SUMB[21][7] ), .Z(\A1[26] ) );
  EO U124 ( .A(\CARRYB[21][7] ), .B(\SUMB[21][8] ), .Z(\A1[27] ) );
  EO U125 ( .A(\CARRYB[21][8] ), .B(\SUMB[21][9] ), .Z(\A1[28] ) );
  EO U126 ( .A(\CARRYB[21][17] ), .B(\SUMB[21][18] ), .Z(\A1[37] ) );
  EO U127 ( .A(\CARRYB[21][13] ), .B(\SUMB[21][14] ), .Z(\A1[33] ) );
  EO U128 ( .A(\CARRYB[21][12] ), .B(\SUMB[21][13] ), .Z(\A1[32] ) );
  EO U129 ( .A(\CARRYB[21][16] ), .B(\SUMB[21][17] ), .Z(\A1[36] ) );
  EO U130 ( .A(\CARRYB[21][18] ), .B(\SUMB[21][19] ), .Z(\A1[38] ) );
  EO U131 ( .A(\CARRYB[21][21] ), .B(\SUMB[21][22] ), .Z(\A1[41] ) );
  EO U132 ( .A(\CARRYB[21][19] ), .B(\SUMB[21][20] ), .Z(\A1[39] ) );
  EO U133 ( .A(\CARRYB[21][20] ), .B(\SUMB[21][21] ), .Z(\A1[40] ) );
  EO U134 ( .A(\CARRYB[21][15] ), .B(\SUMB[21][16] ), .Z(\A1[35] ) );
  EO U135 ( .A(\CARRYB[21][14] ), .B(\SUMB[21][15] ), .Z(\A1[34] ) );
  EO U136 ( .A(\CARRYB[21][22] ), .B(\SUMB[21][23] ), .Z(\A1[42] ) );
  EO U137 ( .A(\CARRYB[21][10] ), .B(\SUMB[21][11] ), .Z(\A1[30] ) );
  EO U138 ( .A(\CARRYB[21][23] ), .B(\SUMB[21][24] ), .Z(\A1[43] ) );
  EO U139 ( .A(\CARRYB[21][11] ), .B(\SUMB[21][12] ), .Z(\A1[31] ) );
  EO U140 ( .A(\CARRYB[21][24] ), .B(\SUMB[21][25] ), .Z(\A1[44] ) );
  EO U141 ( .A(\CARRYB[21][25] ), .B(\SUMB[21][26] ), .Z(\A1[45] ) );
  EO U142 ( .A(\CARRYB[21][26] ), .B(\SUMB[21][27] ), .Z(\A1[46] ) );
  EO U143 ( .A(\CARRYB[21][29] ), .B(\SUMB[21][30] ), .Z(\A1[49] ) );
  EO U144 ( .A(\CARRYB[21][27] ), .B(\SUMB[21][28] ), .Z(\A1[47] ) );
  EO U145 ( .A(\CARRYB[21][30] ), .B(\SUMB[21][31] ), .Z(\A1[50] ) );
  EO U146 ( .A(\CARRYB[21][28] ), .B(\SUMB[21][29] ), .Z(\A1[48] ) );
  EO U147 ( .A(\CARRYB[21][33] ), .B(\SUMB[21][34] ), .Z(\A1[53] ) );
  EO U148 ( .A(\CARRYB[21][34] ), .B(\SUMB[21][35] ), .Z(\A1[54] ) );
  EO U149 ( .A(\CARRYB[21][32] ), .B(\SUMB[21][33] ), .Z(\A1[52] ) );
  EO U150 ( .A(\CARRYB[21][37] ), .B(\SUMB[21][38] ), .Z(\A1[57] ) );
  EO U151 ( .A(\CARRYB[21][31] ), .B(\SUMB[21][32] ), .Z(\A1[51] ) );
  EO U152 ( .A(\CARRYB[21][35] ), .B(\SUMB[21][36] ), .Z(\A1[55] ) );
  EO U153 ( .A(\CARRYB[21][38] ), .B(\SUMB[21][39] ), .Z(\A1[58] ) );
  EO U154 ( .A(\CARRYB[21][36] ), .B(\SUMB[21][37] ), .Z(\A1[56] ) );
  EO U155 ( .A(\CARRYB[21][39] ), .B(\SUMB[21][40] ), .Z(\A1[59] ) );
  EO U156 ( .A(\CARRYB[21][40] ), .B(\SUMB[21][41] ), .Z(\A1[60] ) );
  EO U157 ( .A(\CARRYB[21][41] ), .B(\SUMB[21][42] ), .Z(\A1[61] ) );
  EO U158 ( .A(\CARRYB[21][42] ), .B(\SUMB[21][43] ), .Z(\A1[62] ) );
  EO U159 ( .A(\CARRYB[21][43] ), .B(\SUMB[21][44] ), .Z(\A1[63] ) );
  EO U160 ( .A(\CARRYB[21][44] ), .B(\SUMB[21][45] ), .Z(\A1[64] ) );
  EO U161 ( .A(\CARRYB[21][45] ), .B(\SUMB[21][46] ), .Z(\A1[65] ) );
  EO U162 ( .A(\CARRYB[21][0] ), .B(\SUMB[21][1] ), .Z(\A1[20] ) );
  EO U163 ( .A(\CARRYB[21][46] ), .B(\ab[21][47] ), .Z(\A1[66] ) );
  EO U164 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U165 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U166 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U167 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U168 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U169 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U170 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U171 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U172 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U173 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U174 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U175 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U176 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U177 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U178 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Z(\SUMB[1][18] ) );
  EO U179 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Z(\SUMB[1][19] ) );
  EO U180 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Z(\SUMB[1][16] ) );
  EO U181 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Z(\SUMB[1][17] ) );
  EO U182 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Z(\SUMB[1][20] ) );
  EO U183 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Z(\SUMB[1][22] ) );
  EO U184 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Z(\SUMB[1][23] ) );
  EO U185 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Z(\SUMB[1][21] ) );
  EO U186 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Z(\SUMB[1][24] ) );
  EO U187 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Z(\SUMB[1][25] ) );
  EO U188 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Z(\SUMB[1][26] ) );
  EO U189 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Z(\SUMB[1][27] ) );
  EO U190 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Z(\SUMB[1][28] ) );
  EO U191 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Z(\SUMB[1][29] ) );
  EO U192 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Z(\SUMB[1][30] ) );
  EO U193 ( .A(\ab[0][32] ), .B(\ab[1][31] ), .Z(\SUMB[1][31] ) );
  EO U194 ( .A(\ab[0][33] ), .B(\ab[1][32] ), .Z(\SUMB[1][32] ) );
  EO U195 ( .A(\ab[0][34] ), .B(\ab[1][33] ), .Z(\SUMB[1][33] ) );
  EO U196 ( .A(\ab[0][35] ), .B(\ab[1][34] ), .Z(\SUMB[1][34] ) );
  EO U197 ( .A(\ab[0][36] ), .B(\ab[1][35] ), .Z(\SUMB[1][35] ) );
  EO U198 ( .A(\ab[0][37] ), .B(\ab[1][36] ), .Z(\SUMB[1][36] ) );
  EO U199 ( .A(\ab[0][38] ), .B(\ab[1][37] ), .Z(\SUMB[1][37] ) );
  EO U200 ( .A(\ab[0][39] ), .B(\ab[1][38] ), .Z(\SUMB[1][38] ) );
  EO U201 ( .A(\ab[0][40] ), .B(\ab[1][39] ), .Z(\SUMB[1][39] ) );
  EO U202 ( .A(\ab[0][41] ), .B(\ab[1][40] ), .Z(\SUMB[1][40] ) );
  EO U203 ( .A(\ab[0][42] ), .B(\ab[1][41] ), .Z(\SUMB[1][41] ) );
  EO U204 ( .A(\ab[0][43] ), .B(\ab[1][42] ), .Z(\SUMB[1][42] ) );
  EO U205 ( .A(\ab[0][44] ), .B(\ab[1][43] ), .Z(\SUMB[1][43] ) );
  EO U206 ( .A(\ab[0][45] ), .B(\ab[1][44] ), .Z(\SUMB[1][44] ) );
  EO U207 ( .A(\ab[0][46] ), .B(\ab[1][45] ), .Z(\SUMB[1][45] ) );
  EO U208 ( .A(\ab[0][47] ), .B(\ab[1][46] ), .Z(\SUMB[1][46] ) );
  IVP U209 ( .A(B[2]), .Z(n162) );
  IVP U210 ( .A(B[3]), .Z(n161) );
  IVP U211 ( .A(B[4]), .Z(n160) );
  IVP U212 ( .A(B[1]), .Z(n163) );
  IVP U213 ( .A(B[5]), .Z(n159) );
  IVP U214 ( .A(B[0]), .Z(n164) );
  IVP U215 ( .A(B[6]), .Z(n158) );
  IVP U216 ( .A(B[7]), .Z(n157) );
  IVP U217 ( .A(B[8]), .Z(n156) );
  IVP U218 ( .A(B[9]), .Z(n155) );
  IVP U219 ( .A(B[10]), .Z(n154) );
  IVP U220 ( .A(B[11]), .Z(n153) );
  IVP U221 ( .A(B[12]), .Z(n152) );
  IVP U222 ( .A(B[13]), .Z(n151) );
  IVP U223 ( .A(B[14]), .Z(n150) );
  IVP U224 ( .A(B[15]), .Z(n149) );
  IVP U225 ( .A(B[16]), .Z(n148) );
  IVP U226 ( .A(B[17]), .Z(n147) );
  IVP U227 ( .A(B[18]), .Z(n146) );
  IVP U228 ( .A(B[19]), .Z(n145) );
  IVP U229 ( .A(B[20]), .Z(n144) );
  IVP U230 ( .A(B[21]), .Z(n143) );
  IVP U231 ( .A(B[22]), .Z(n142) );
  IVP U232 ( .A(B[23]), .Z(n141) );
  IVP U233 ( .A(B[24]), .Z(n140) );
  IVP U234 ( .A(B[25]), .Z(n139) );
  IVP U235 ( .A(B[26]), .Z(n138) );
  IVP U236 ( .A(B[27]), .Z(n137) );
  IVP U237 ( .A(B[28]), .Z(n136) );
  IVP U238 ( .A(B[29]), .Z(n135) );
  IVP U239 ( .A(B[30]), .Z(n134) );
  IVP U240 ( .A(B[31]), .Z(n133) );
  IVP U241 ( .A(B[32]), .Z(n132) );
  IVP U242 ( .A(B[33]), .Z(n131) );
  IVP U243 ( .A(B[34]), .Z(n130) );
  IVP U244 ( .A(B[35]), .Z(n129) );
  IVP U245 ( .A(B[36]), .Z(n128) );
  IVP U246 ( .A(B[37]), .Z(n127) );
  IVP U247 ( .A(B[38]), .Z(n126) );
  IVP U248 ( .A(B[39]), .Z(n125) );
  IVP U249 ( .A(B[40]), .Z(n101) );
  IVP U250 ( .A(B[41]), .Z(n102) );
  IVP U251 ( .A(B[42]), .Z(n103) );
  IVP U252 ( .A(B[43]), .Z(n104) );
  IVP U253 ( .A(B[44]), .Z(n105) );
  IVP U254 ( .A(B[45]), .Z(n106) );
  IVP U255 ( .A(B[47]), .Z(n108) );
  IVP U256 ( .A(B[46]), .Z(n107) );
  AN2P U257 ( .A(\CARRYB[21][0] ), .B(\SUMB[21][1] ), .Z(\A2[21] ) );
  AN2P U258 ( .A(\CARRYB[21][1] ), .B(\SUMB[21][2] ), .Z(\A2[22] ) );
  AN2P U259 ( .A(\CARRYB[21][2] ), .B(\SUMB[21][3] ), .Z(\A2[23] ) );
  AN2P U260 ( .A(\CARRYB[21][3] ), .B(\SUMB[21][4] ), .Z(\A2[24] ) );
  AN2P U261 ( .A(\CARRYB[21][4] ), .B(\SUMB[21][5] ), .Z(\A2[25] ) );
  AN2P U262 ( .A(\CARRYB[21][5] ), .B(\SUMB[21][6] ), .Z(\A2[26] ) );
  AN2P U263 ( .A(\CARRYB[21][6] ), .B(\SUMB[21][7] ), .Z(\A2[27] ) );
  AN2P U264 ( .A(\CARRYB[21][7] ), .B(\SUMB[21][8] ), .Z(\A2[28] ) );
  AN2P U265 ( .A(\CARRYB[21][8] ), .B(\SUMB[21][9] ), .Z(\A2[29] ) );
  AN2P U266 ( .A(\CARRYB[21][9] ), .B(\SUMB[21][10] ), .Z(\A2[30] ) );
  AN2P U267 ( .A(\CARRYB[21][10] ), .B(\SUMB[21][11] ), .Z(\A2[31] ) );
  AN2P U268 ( .A(\CARRYB[21][11] ), .B(\SUMB[21][12] ), .Z(\A2[32] ) );
  AN2P U269 ( .A(\CARRYB[21][12] ), .B(\SUMB[21][13] ), .Z(\A2[33] ) );
  AN2P U270 ( .A(\CARRYB[21][13] ), .B(\SUMB[21][14] ), .Z(\A2[34] ) );
  AN2P U271 ( .A(\CARRYB[21][14] ), .B(\SUMB[21][15] ), .Z(\A2[35] ) );
  AN2P U272 ( .A(\CARRYB[21][15] ), .B(\SUMB[21][16] ), .Z(\A2[36] ) );
  AN2P U273 ( .A(\CARRYB[21][16] ), .B(\SUMB[21][17] ), .Z(\A2[37] ) );
  AN2P U274 ( .A(\CARRYB[21][17] ), .B(\SUMB[21][18] ), .Z(\A2[38] ) );
  AN2P U275 ( .A(\CARRYB[21][18] ), .B(\SUMB[21][19] ), .Z(\A2[39] ) );
  AN2P U276 ( .A(\CARRYB[21][19] ), .B(\SUMB[21][20] ), .Z(\A2[40] ) );
  AN2P U277 ( .A(\CARRYB[21][20] ), .B(\SUMB[21][21] ), .Z(\A2[41] ) );
  AN2P U278 ( .A(\CARRYB[21][21] ), .B(\SUMB[21][22] ), .Z(\A2[42] ) );
  AN2P U279 ( .A(\CARRYB[21][22] ), .B(\SUMB[21][23] ), .Z(\A2[43] ) );
  AN2P U280 ( .A(\CARRYB[21][23] ), .B(\SUMB[21][24] ), .Z(\A2[44] ) );
  AN2P U281 ( .A(\CARRYB[21][24] ), .B(\SUMB[21][25] ), .Z(\A2[45] ) );
  AN2P U282 ( .A(\CARRYB[21][26] ), .B(\SUMB[21][27] ), .Z(\A2[47] ) );
  AN2P U283 ( .A(\CARRYB[21][27] ), .B(\SUMB[21][28] ), .Z(\A2[48] ) );
  AN2P U284 ( .A(\CARRYB[21][28] ), .B(\SUMB[21][29] ), .Z(\A2[49] ) );
  AN2P U285 ( .A(\CARRYB[21][29] ), .B(\SUMB[21][30] ), .Z(\A2[50] ) );
  AN2P U286 ( .A(\CARRYB[21][30] ), .B(\SUMB[21][31] ), .Z(\A2[51] ) );
  AN2P U287 ( .A(\CARRYB[21][31] ), .B(\SUMB[21][32] ), .Z(\A2[52] ) );
  AN2P U288 ( .A(\CARRYB[21][32] ), .B(\SUMB[21][33] ), .Z(\A2[53] ) );
  AN2P U289 ( .A(\CARRYB[21][33] ), .B(\SUMB[21][34] ), .Z(\A2[54] ) );
  AN2P U290 ( .A(\CARRYB[21][34] ), .B(\SUMB[21][35] ), .Z(\A2[55] ) );
  AN2P U291 ( .A(\CARRYB[21][35] ), .B(\SUMB[21][36] ), .Z(\A2[56] ) );
  AN2P U292 ( .A(\CARRYB[21][36] ), .B(\SUMB[21][37] ), .Z(\A2[57] ) );
  AN2P U293 ( .A(\CARRYB[21][37] ), .B(\SUMB[21][38] ), .Z(\A2[58] ) );
  AN2P U294 ( .A(\CARRYB[21][38] ), .B(\SUMB[21][39] ), .Z(\A2[59] ) );
  AN2P U295 ( .A(\CARRYB[21][39] ), .B(\SUMB[21][40] ), .Z(\A2[60] ) );
  AN2P U296 ( .A(\CARRYB[21][40] ), .B(\SUMB[21][41] ), .Z(\A2[61] ) );
  AN2P U297 ( .A(\CARRYB[21][41] ), .B(\SUMB[21][42] ), .Z(\A2[62] ) );
  AN2P U298 ( .A(\CARRYB[21][42] ), .B(\SUMB[21][43] ), .Z(\A2[63] ) );
  AN2P U299 ( .A(\CARRYB[21][43] ), .B(\SUMB[21][44] ), .Z(\A2[64] ) );
  AN2P U300 ( .A(\CARRYB[21][44] ), .B(\SUMB[21][45] ), .Z(\A2[65] ) );
  AN2P U301 ( .A(\CARRYB[21][45] ), .B(\SUMB[21][46] ), .Z(\A2[66] ) );
  AN2P U302 ( .A(\CARRYB[21][46] ), .B(\ab[21][47] ), .Z(\A2[67] ) );
  AN2P U303 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U304 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U305 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U306 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U307 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U308 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U309 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U310 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U311 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U312 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U313 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U314 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U315 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U316 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U317 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U318 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\CARRYB[1][16] ) );
  AN2P U319 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\CARRYB[1][17] ) );
  AN2P U320 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\CARRYB[1][18] ) );
  AN2P U321 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\CARRYB[1][19] ) );
  AN2P U322 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\CARRYB[1][20] ) );
  AN2P U323 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\CARRYB[1][21] ) );
  AN2P U324 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(\CARRYB[1][22] ) );
  AN2P U325 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(\CARRYB[1][23] ) );
  AN2P U326 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(\CARRYB[1][24] ) );
  AN2P U327 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(\CARRYB[1][25] ) );
  AN2P U328 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\CARRYB[1][26] ) );
  AN2P U329 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(\CARRYB[1][27] ) );
  AN2P U330 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(\CARRYB[1][28] ) );
  AN2P U331 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(\CARRYB[1][29] ) );
  AN2P U332 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(\CARRYB[1][30] ) );
  AN2P U333 ( .A(\ab[1][31] ), .B(\ab[0][32] ), .Z(\CARRYB[1][31] ) );
  AN2P U334 ( .A(\ab[1][32] ), .B(\ab[0][33] ), .Z(\CARRYB[1][32] ) );
  AN2P U335 ( .A(\ab[1][33] ), .B(\ab[0][34] ), .Z(\CARRYB[1][33] ) );
  AN2P U336 ( .A(\ab[1][34] ), .B(\ab[0][35] ), .Z(\CARRYB[1][34] ) );
  AN2P U337 ( .A(\ab[1][35] ), .B(\ab[0][36] ), .Z(\CARRYB[1][35] ) );
  AN2P U338 ( .A(\ab[1][36] ), .B(\ab[0][37] ), .Z(\CARRYB[1][36] ) );
  AN2P U339 ( .A(\ab[1][37] ), .B(\ab[0][38] ), .Z(\CARRYB[1][37] ) );
  AN2P U340 ( .A(\ab[1][38] ), .B(\ab[0][39] ), .Z(\CARRYB[1][38] ) );
  AN2P U341 ( .A(\ab[1][39] ), .B(\ab[0][40] ), .Z(\CARRYB[1][39] ) );
  AN2P U342 ( .A(\ab[1][40] ), .B(\ab[0][41] ), .Z(\CARRYB[1][40] ) );
  AN2P U343 ( .A(\ab[1][41] ), .B(\ab[0][42] ), .Z(\CARRYB[1][41] ) );
  AN2P U344 ( .A(\ab[1][42] ), .B(\ab[0][43] ), .Z(\CARRYB[1][42] ) );
  AN2P U345 ( .A(\ab[1][43] ), .B(\ab[0][44] ), .Z(\CARRYB[1][43] ) );
  AN2P U346 ( .A(\ab[1][44] ), .B(\ab[0][45] ), .Z(\CARRYB[1][44] ) );
  AN2P U347 ( .A(\ab[1][45] ), .B(\ab[0][46] ), .Z(\CARRYB[1][45] ) );
  AN2P U348 ( .A(\ab[1][46] ), .B(\ab[0][47] ), .Z(\CARRYB[1][46] ) );
  AN2P U349 ( .A(\CARRYB[21][25] ), .B(\SUMB[21][26] ), .Z(\A2[46] ) );
  NR2 U351 ( .A(n84), .B(n155), .Z(\ab[9][9] ) );
  NR2 U352 ( .A(n84), .B(n156), .Z(\ab[9][8] ) );
  NR2 U353 ( .A(n84), .B(n157), .Z(\ab[9][7] ) );
  NR2 U354 ( .A(n84), .B(n158), .Z(\ab[9][6] ) );
  NR2 U355 ( .A(n84), .B(n159), .Z(\ab[9][5] ) );
  NR2 U356 ( .A(n84), .B(n160), .Z(\ab[9][4] ) );
  NR2 U357 ( .A(n84), .B(n108), .Z(\ab[9][47] ) );
  NR2 U358 ( .A(n84), .B(n107), .Z(\ab[9][46] ) );
  NR2 U359 ( .A(n84), .B(n106), .Z(\ab[9][45] ) );
  NR2 U360 ( .A(n84), .B(n105), .Z(\ab[9][44] ) );
  NR2 U361 ( .A(n84), .B(n104), .Z(\ab[9][43] ) );
  NR2 U362 ( .A(n84), .B(n103), .Z(\ab[9][42] ) );
  NR2 U363 ( .A(n83), .B(n102), .Z(\ab[9][41] ) );
  NR2 U364 ( .A(n83), .B(n101), .Z(\ab[9][40] ) );
  NR2 U365 ( .A(n83), .B(n161), .Z(\ab[9][3] ) );
  NR2 U366 ( .A(n83), .B(n125), .Z(\ab[9][39] ) );
  NR2 U367 ( .A(n83), .B(n126), .Z(\ab[9][38] ) );
  NR2 U368 ( .A(n83), .B(n127), .Z(\ab[9][37] ) );
  NR2 U369 ( .A(n83), .B(n128), .Z(\ab[9][36] ) );
  NR2 U370 ( .A(n83), .B(n129), .Z(\ab[9][35] ) );
  NR2 U371 ( .A(n83), .B(n130), .Z(\ab[9][34] ) );
  NR2 U372 ( .A(n83), .B(n131), .Z(\ab[9][33] ) );
  NR2 U373 ( .A(n83), .B(n132), .Z(\ab[9][32] ) );
  NR2 U374 ( .A(n83), .B(n133), .Z(\ab[9][31] ) );
  NR2 U375 ( .A(n82), .B(n134), .Z(\ab[9][30] ) );
  NR2 U376 ( .A(n82), .B(n162), .Z(\ab[9][2] ) );
  NR2 U377 ( .A(n82), .B(n135), .Z(\ab[9][29] ) );
  NR2 U378 ( .A(n82), .B(n136), .Z(\ab[9][28] ) );
  NR2 U379 ( .A(n82), .B(n137), .Z(\ab[9][27] ) );
  NR2 U380 ( .A(n82), .B(n138), .Z(\ab[9][26] ) );
  NR2 U381 ( .A(n82), .B(n139), .Z(\ab[9][25] ) );
  NR2 U382 ( .A(n82), .B(n140), .Z(\ab[9][24] ) );
  NR2 U383 ( .A(n82), .B(n141), .Z(\ab[9][23] ) );
  NR2 U384 ( .A(n82), .B(n142), .Z(\ab[9][22] ) );
  NR2 U385 ( .A(n82), .B(n143), .Z(\ab[9][21] ) );
  NR2 U386 ( .A(n82), .B(n144), .Z(\ab[9][20] ) );
  NR2 U387 ( .A(n81), .B(n163), .Z(\ab[9][1] ) );
  NR2 U388 ( .A(n81), .B(n145), .Z(\ab[9][19] ) );
  NR2 U389 ( .A(n81), .B(n146), .Z(\ab[9][18] ) );
  NR2 U390 ( .A(n81), .B(n147), .Z(\ab[9][17] ) );
  NR2 U391 ( .A(n81), .B(n148), .Z(\ab[9][16] ) );
  NR2 U392 ( .A(n81), .B(n149), .Z(\ab[9][15] ) );
  NR2 U393 ( .A(n81), .B(n150), .Z(\ab[9][14] ) );
  NR2 U394 ( .A(n81), .B(n151), .Z(\ab[9][13] ) );
  NR2 U395 ( .A(n81), .B(n152), .Z(\ab[9][12] ) );
  NR2 U396 ( .A(n81), .B(n153), .Z(\ab[9][11] ) );
  NR2 U397 ( .A(n81), .B(n154), .Z(\ab[9][10] ) );
  NR2 U398 ( .A(n81), .B(n164), .Z(\ab[9][0] ) );
  NR2 U399 ( .A(n155), .B(n79), .Z(\ab[8][9] ) );
  NR2 U400 ( .A(n156), .B(n79), .Z(\ab[8][8] ) );
  NR2 U401 ( .A(n157), .B(n79), .Z(\ab[8][7] ) );
  NR2 U402 ( .A(n158), .B(n79), .Z(\ab[8][6] ) );
  NR2 U403 ( .A(n159), .B(n79), .Z(\ab[8][5] ) );
  NR2 U404 ( .A(n160), .B(n79), .Z(\ab[8][4] ) );
  NR2 U405 ( .A(n108), .B(n79), .Z(\ab[8][47] ) );
  NR2 U406 ( .A(n107), .B(n79), .Z(\ab[8][46] ) );
  NR2 U407 ( .A(n106), .B(n79), .Z(\ab[8][45] ) );
  NR2 U408 ( .A(n105), .B(n79), .Z(\ab[8][44] ) );
  NR2 U409 ( .A(n104), .B(n79), .Z(\ab[8][43] ) );
  NR2 U410 ( .A(n103), .B(n79), .Z(\ab[8][42] ) );
  NR2 U411 ( .A(n102), .B(n78), .Z(\ab[8][41] ) );
  NR2 U412 ( .A(n101), .B(n78), .Z(\ab[8][40] ) );
  NR2 U413 ( .A(n161), .B(n78), .Z(\ab[8][3] ) );
  NR2 U414 ( .A(n125), .B(n78), .Z(\ab[8][39] ) );
  NR2 U415 ( .A(n126), .B(n78), .Z(\ab[8][38] ) );
  NR2 U416 ( .A(n127), .B(n78), .Z(\ab[8][37] ) );
  NR2 U417 ( .A(n128), .B(n78), .Z(\ab[8][36] ) );
  NR2 U418 ( .A(n129), .B(n78), .Z(\ab[8][35] ) );
  NR2 U419 ( .A(n130), .B(n78), .Z(\ab[8][34] ) );
  NR2 U420 ( .A(n131), .B(n78), .Z(\ab[8][33] ) );
  NR2 U421 ( .A(n132), .B(n78), .Z(\ab[8][32] ) );
  NR2 U422 ( .A(n133), .B(n78), .Z(\ab[8][31] ) );
  NR2 U423 ( .A(n134), .B(n77), .Z(\ab[8][30] ) );
  NR2 U424 ( .A(n162), .B(n77), .Z(\ab[8][2] ) );
  NR2 U425 ( .A(n135), .B(n77), .Z(\ab[8][29] ) );
  NR2 U426 ( .A(n136), .B(n77), .Z(\ab[8][28] ) );
  NR2 U427 ( .A(n137), .B(n77), .Z(\ab[8][27] ) );
  NR2 U428 ( .A(n138), .B(n77), .Z(\ab[8][26] ) );
  NR2 U429 ( .A(n139), .B(n77), .Z(\ab[8][25] ) );
  NR2 U430 ( .A(n140), .B(n77), .Z(\ab[8][24] ) );
  NR2 U431 ( .A(n141), .B(n77), .Z(\ab[8][23] ) );
  NR2 U432 ( .A(n142), .B(n77), .Z(\ab[8][22] ) );
  NR2 U433 ( .A(n143), .B(n77), .Z(\ab[8][21] ) );
  NR2 U434 ( .A(n144), .B(n77), .Z(\ab[8][20] ) );
  NR2 U435 ( .A(n163), .B(n76), .Z(\ab[8][1] ) );
  NR2 U436 ( .A(n145), .B(n76), .Z(\ab[8][19] ) );
  NR2 U437 ( .A(n146), .B(n76), .Z(\ab[8][18] ) );
  NR2 U438 ( .A(n147), .B(n76), .Z(\ab[8][17] ) );
  NR2 U439 ( .A(n148), .B(n76), .Z(\ab[8][16] ) );
  NR2 U440 ( .A(n149), .B(n76), .Z(\ab[8][15] ) );
  NR2 U441 ( .A(n150), .B(n76), .Z(\ab[8][14] ) );
  NR2 U442 ( .A(n151), .B(n76), .Z(\ab[8][13] ) );
  NR2 U443 ( .A(n152), .B(n76), .Z(\ab[8][12] ) );
  NR2 U444 ( .A(n153), .B(n76), .Z(\ab[8][11] ) );
  NR2 U445 ( .A(n154), .B(n76), .Z(\ab[8][10] ) );
  NR2 U446 ( .A(n164), .B(n76), .Z(\ab[8][0] ) );
  NR2 U447 ( .A(n155), .B(n74), .Z(\ab[7][9] ) );
  NR2 U448 ( .A(n156), .B(n74), .Z(\ab[7][8] ) );
  NR2 U449 ( .A(n157), .B(n74), .Z(\ab[7][7] ) );
  NR2 U450 ( .A(n158), .B(n74), .Z(\ab[7][6] ) );
  NR2 U451 ( .A(n159), .B(n74), .Z(\ab[7][5] ) );
  NR2 U452 ( .A(n160), .B(n74), .Z(\ab[7][4] ) );
  NR2 U453 ( .A(n108), .B(n74), .Z(\ab[7][47] ) );
  NR2 U454 ( .A(n107), .B(n74), .Z(\ab[7][46] ) );
  NR2 U455 ( .A(n106), .B(n74), .Z(\ab[7][45] ) );
  NR2 U456 ( .A(n105), .B(n74), .Z(\ab[7][44] ) );
  NR2 U457 ( .A(n104), .B(n74), .Z(\ab[7][43] ) );
  NR2 U458 ( .A(n103), .B(n74), .Z(\ab[7][42] ) );
  NR2 U459 ( .A(n102), .B(n73), .Z(\ab[7][41] ) );
  NR2 U460 ( .A(n101), .B(n73), .Z(\ab[7][40] ) );
  NR2 U461 ( .A(n161), .B(n73), .Z(\ab[7][3] ) );
  NR2 U462 ( .A(n125), .B(n73), .Z(\ab[7][39] ) );
  NR2 U463 ( .A(n126), .B(n73), .Z(\ab[7][38] ) );
  NR2 U464 ( .A(n127), .B(n73), .Z(\ab[7][37] ) );
  NR2 U465 ( .A(n128), .B(n73), .Z(\ab[7][36] ) );
  NR2 U466 ( .A(n129), .B(n73), .Z(\ab[7][35] ) );
  NR2 U467 ( .A(n130), .B(n73), .Z(\ab[7][34] ) );
  NR2 U468 ( .A(n131), .B(n73), .Z(\ab[7][33] ) );
  NR2 U469 ( .A(n132), .B(n73), .Z(\ab[7][32] ) );
  NR2 U470 ( .A(n133), .B(n73), .Z(\ab[7][31] ) );
  NR2 U471 ( .A(n134), .B(n72), .Z(\ab[7][30] ) );
  NR2 U472 ( .A(n162), .B(n72), .Z(\ab[7][2] ) );
  NR2 U473 ( .A(n135), .B(n72), .Z(\ab[7][29] ) );
  NR2 U474 ( .A(n136), .B(n72), .Z(\ab[7][28] ) );
  NR2 U475 ( .A(n137), .B(n72), .Z(\ab[7][27] ) );
  NR2 U476 ( .A(n138), .B(n72), .Z(\ab[7][26] ) );
  NR2 U477 ( .A(n139), .B(n72), .Z(\ab[7][25] ) );
  NR2 U478 ( .A(n140), .B(n72), .Z(\ab[7][24] ) );
  NR2 U479 ( .A(n141), .B(n72), .Z(\ab[7][23] ) );
  NR2 U480 ( .A(n142), .B(n72), .Z(\ab[7][22] ) );
  NR2 U481 ( .A(n143), .B(n72), .Z(\ab[7][21] ) );
  NR2 U482 ( .A(n144), .B(n72), .Z(\ab[7][20] ) );
  NR2 U483 ( .A(n163), .B(n71), .Z(\ab[7][1] ) );
  NR2 U484 ( .A(n145), .B(n71), .Z(\ab[7][19] ) );
  NR2 U485 ( .A(n146), .B(n71), .Z(\ab[7][18] ) );
  NR2 U486 ( .A(n147), .B(n71), .Z(\ab[7][17] ) );
  NR2 U487 ( .A(n148), .B(n71), .Z(\ab[7][16] ) );
  NR2 U488 ( .A(n149), .B(n71), .Z(\ab[7][15] ) );
  NR2 U489 ( .A(n150), .B(n71), .Z(\ab[7][14] ) );
  NR2 U490 ( .A(n151), .B(n71), .Z(\ab[7][13] ) );
  NR2 U491 ( .A(n152), .B(n71), .Z(\ab[7][12] ) );
  NR2 U492 ( .A(n153), .B(n71), .Z(\ab[7][11] ) );
  NR2 U493 ( .A(n154), .B(n71), .Z(\ab[7][10] ) );
  NR2 U494 ( .A(n164), .B(n71), .Z(\ab[7][0] ) );
  NR2 U495 ( .A(n155), .B(n69), .Z(\ab[6][9] ) );
  NR2 U496 ( .A(n156), .B(n69), .Z(\ab[6][8] ) );
  NR2 U497 ( .A(n157), .B(n69), .Z(\ab[6][7] ) );
  NR2 U498 ( .A(n158), .B(n69), .Z(\ab[6][6] ) );
  NR2 U499 ( .A(n159), .B(n69), .Z(\ab[6][5] ) );
  NR2 U500 ( .A(n160), .B(n69), .Z(\ab[6][4] ) );
  NR2 U501 ( .A(n108), .B(n69), .Z(\ab[6][47] ) );
  NR2 U502 ( .A(n107), .B(n69), .Z(\ab[6][46] ) );
  NR2 U503 ( .A(n106), .B(n69), .Z(\ab[6][45] ) );
  NR2 U504 ( .A(n105), .B(n69), .Z(\ab[6][44] ) );
  NR2 U505 ( .A(n104), .B(n69), .Z(\ab[6][43] ) );
  NR2 U506 ( .A(n103), .B(n69), .Z(\ab[6][42] ) );
  NR2 U507 ( .A(n102), .B(n68), .Z(\ab[6][41] ) );
  NR2 U508 ( .A(n101), .B(n68), .Z(\ab[6][40] ) );
  NR2 U509 ( .A(n161), .B(n68), .Z(\ab[6][3] ) );
  NR2 U510 ( .A(n125), .B(n68), .Z(\ab[6][39] ) );
  NR2 U511 ( .A(n126), .B(n68), .Z(\ab[6][38] ) );
  NR2 U512 ( .A(n127), .B(n68), .Z(\ab[6][37] ) );
  NR2 U513 ( .A(n128), .B(n68), .Z(\ab[6][36] ) );
  NR2 U514 ( .A(n129), .B(n68), .Z(\ab[6][35] ) );
  NR2 U515 ( .A(n130), .B(n68), .Z(\ab[6][34] ) );
  NR2 U516 ( .A(n131), .B(n68), .Z(\ab[6][33] ) );
  NR2 U517 ( .A(n132), .B(n68), .Z(\ab[6][32] ) );
  NR2 U518 ( .A(n133), .B(n68), .Z(\ab[6][31] ) );
  NR2 U519 ( .A(n134), .B(n67), .Z(\ab[6][30] ) );
  NR2 U520 ( .A(n162), .B(n67), .Z(\ab[6][2] ) );
  NR2 U521 ( .A(n135), .B(n67), .Z(\ab[6][29] ) );
  NR2 U522 ( .A(n136), .B(n67), .Z(\ab[6][28] ) );
  NR2 U523 ( .A(n137), .B(n67), .Z(\ab[6][27] ) );
  NR2 U524 ( .A(n138), .B(n67), .Z(\ab[6][26] ) );
  NR2 U525 ( .A(n139), .B(n67), .Z(\ab[6][25] ) );
  NR2 U526 ( .A(n140), .B(n67), .Z(\ab[6][24] ) );
  NR2 U527 ( .A(n141), .B(n67), .Z(\ab[6][23] ) );
  NR2 U528 ( .A(n142), .B(n67), .Z(\ab[6][22] ) );
  NR2 U529 ( .A(n143), .B(n67), .Z(\ab[6][21] ) );
  NR2 U530 ( .A(n144), .B(n67), .Z(\ab[6][20] ) );
  NR2 U531 ( .A(n163), .B(n66), .Z(\ab[6][1] ) );
  NR2 U532 ( .A(n145), .B(n66), .Z(\ab[6][19] ) );
  NR2 U533 ( .A(n146), .B(n66), .Z(\ab[6][18] ) );
  NR2 U534 ( .A(n147), .B(n66), .Z(\ab[6][17] ) );
  NR2 U535 ( .A(n148), .B(n66), .Z(\ab[6][16] ) );
  NR2 U536 ( .A(n149), .B(n66), .Z(\ab[6][15] ) );
  NR2 U537 ( .A(n150), .B(n66), .Z(\ab[6][14] ) );
  NR2 U538 ( .A(n151), .B(n66), .Z(\ab[6][13] ) );
  NR2 U539 ( .A(n152), .B(n66), .Z(\ab[6][12] ) );
  NR2 U540 ( .A(n153), .B(n66), .Z(\ab[6][11] ) );
  NR2 U541 ( .A(n154), .B(n66), .Z(\ab[6][10] ) );
  NR2 U542 ( .A(n164), .B(n66), .Z(\ab[6][0] ) );
  NR2 U543 ( .A(n155), .B(n64), .Z(\ab[5][9] ) );
  NR2 U544 ( .A(n156), .B(n64), .Z(\ab[5][8] ) );
  NR2 U545 ( .A(n157), .B(n64), .Z(\ab[5][7] ) );
  NR2 U546 ( .A(n158), .B(n64), .Z(\ab[5][6] ) );
  NR2 U547 ( .A(n159), .B(n64), .Z(\ab[5][5] ) );
  NR2 U548 ( .A(n160), .B(n64), .Z(\ab[5][4] ) );
  NR2 U549 ( .A(n108), .B(n64), .Z(\ab[5][47] ) );
  NR2 U550 ( .A(n107), .B(n64), .Z(\ab[5][46] ) );
  NR2 U551 ( .A(n106), .B(n64), .Z(\ab[5][45] ) );
  NR2 U552 ( .A(n105), .B(n64), .Z(\ab[5][44] ) );
  NR2 U553 ( .A(n104), .B(n64), .Z(\ab[5][43] ) );
  NR2 U554 ( .A(n103), .B(n64), .Z(\ab[5][42] ) );
  NR2 U555 ( .A(n102), .B(n63), .Z(\ab[5][41] ) );
  NR2 U556 ( .A(n101), .B(n63), .Z(\ab[5][40] ) );
  NR2 U557 ( .A(n161), .B(n63), .Z(\ab[5][3] ) );
  NR2 U558 ( .A(n125), .B(n63), .Z(\ab[5][39] ) );
  NR2 U559 ( .A(n126), .B(n63), .Z(\ab[5][38] ) );
  NR2 U560 ( .A(n127), .B(n63), .Z(\ab[5][37] ) );
  NR2 U561 ( .A(n128), .B(n63), .Z(\ab[5][36] ) );
  NR2 U562 ( .A(n129), .B(n63), .Z(\ab[5][35] ) );
  NR2 U563 ( .A(n130), .B(n63), .Z(\ab[5][34] ) );
  NR2 U564 ( .A(n131), .B(n63), .Z(\ab[5][33] ) );
  NR2 U565 ( .A(n132), .B(n63), .Z(\ab[5][32] ) );
  NR2 U566 ( .A(n133), .B(n63), .Z(\ab[5][31] ) );
  NR2 U567 ( .A(n134), .B(n62), .Z(\ab[5][30] ) );
  NR2 U568 ( .A(n162), .B(n62), .Z(\ab[5][2] ) );
  NR2 U569 ( .A(n135), .B(n62), .Z(\ab[5][29] ) );
  NR2 U570 ( .A(n136), .B(n62), .Z(\ab[5][28] ) );
  NR2 U571 ( .A(n137), .B(n62), .Z(\ab[5][27] ) );
  NR2 U572 ( .A(n138), .B(n62), .Z(\ab[5][26] ) );
  NR2 U573 ( .A(n139), .B(n62), .Z(\ab[5][25] ) );
  NR2 U574 ( .A(n140), .B(n62), .Z(\ab[5][24] ) );
  NR2 U575 ( .A(n141), .B(n62), .Z(\ab[5][23] ) );
  NR2 U576 ( .A(n142), .B(n62), .Z(\ab[5][22] ) );
  NR2 U577 ( .A(n143), .B(n62), .Z(\ab[5][21] ) );
  NR2 U578 ( .A(n144), .B(n62), .Z(\ab[5][20] ) );
  NR2 U579 ( .A(n163), .B(n61), .Z(\ab[5][1] ) );
  NR2 U580 ( .A(n145), .B(n61), .Z(\ab[5][19] ) );
  NR2 U581 ( .A(n146), .B(n61), .Z(\ab[5][18] ) );
  NR2 U582 ( .A(n147), .B(n61), .Z(\ab[5][17] ) );
  NR2 U583 ( .A(n148), .B(n61), .Z(\ab[5][16] ) );
  NR2 U584 ( .A(n149), .B(n61), .Z(\ab[5][15] ) );
  NR2 U585 ( .A(n150), .B(n61), .Z(\ab[5][14] ) );
  NR2 U586 ( .A(n151), .B(n61), .Z(\ab[5][13] ) );
  NR2 U587 ( .A(n152), .B(n61), .Z(\ab[5][12] ) );
  NR2 U588 ( .A(n153), .B(n61), .Z(\ab[5][11] ) );
  NR2 U589 ( .A(n154), .B(n61), .Z(\ab[5][10] ) );
  NR2 U590 ( .A(n164), .B(n61), .Z(\ab[5][0] ) );
  NR2 U591 ( .A(n155), .B(n59), .Z(\ab[4][9] ) );
  NR2 U592 ( .A(n156), .B(n59), .Z(\ab[4][8] ) );
  NR2 U593 ( .A(n157), .B(n59), .Z(\ab[4][7] ) );
  NR2 U594 ( .A(n158), .B(n59), .Z(\ab[4][6] ) );
  NR2 U595 ( .A(n159), .B(n59), .Z(\ab[4][5] ) );
  NR2 U596 ( .A(n160), .B(n59), .Z(\ab[4][4] ) );
  NR2 U597 ( .A(n108), .B(n59), .Z(\ab[4][47] ) );
  NR2 U598 ( .A(n107), .B(n59), .Z(\ab[4][46] ) );
  NR2 U599 ( .A(n106), .B(n59), .Z(\ab[4][45] ) );
  NR2 U600 ( .A(n105), .B(n59), .Z(\ab[4][44] ) );
  NR2 U601 ( .A(n104), .B(n59), .Z(\ab[4][43] ) );
  NR2 U602 ( .A(n103), .B(n59), .Z(\ab[4][42] ) );
  NR2 U603 ( .A(n102), .B(n58), .Z(\ab[4][41] ) );
  NR2 U604 ( .A(n101), .B(n58), .Z(\ab[4][40] ) );
  NR2 U605 ( .A(n161), .B(n58), .Z(\ab[4][3] ) );
  NR2 U606 ( .A(n125), .B(n58), .Z(\ab[4][39] ) );
  NR2 U607 ( .A(n126), .B(n58), .Z(\ab[4][38] ) );
  NR2 U608 ( .A(n127), .B(n58), .Z(\ab[4][37] ) );
  NR2 U609 ( .A(n128), .B(n58), .Z(\ab[4][36] ) );
  NR2 U610 ( .A(n129), .B(n58), .Z(\ab[4][35] ) );
  NR2 U611 ( .A(n130), .B(n58), .Z(\ab[4][34] ) );
  NR2 U612 ( .A(n131), .B(n58), .Z(\ab[4][33] ) );
  NR2 U613 ( .A(n132), .B(n58), .Z(\ab[4][32] ) );
  NR2 U614 ( .A(n133), .B(n58), .Z(\ab[4][31] ) );
  NR2 U615 ( .A(n134), .B(n57), .Z(\ab[4][30] ) );
  NR2 U616 ( .A(n162), .B(n57), .Z(\ab[4][2] ) );
  NR2 U617 ( .A(n135), .B(n57), .Z(\ab[4][29] ) );
  NR2 U618 ( .A(n136), .B(n57), .Z(\ab[4][28] ) );
  NR2 U619 ( .A(n137), .B(n57), .Z(\ab[4][27] ) );
  NR2 U620 ( .A(n138), .B(n57), .Z(\ab[4][26] ) );
  NR2 U621 ( .A(n139), .B(n57), .Z(\ab[4][25] ) );
  NR2 U622 ( .A(n140), .B(n57), .Z(\ab[4][24] ) );
  NR2 U623 ( .A(n141), .B(n57), .Z(\ab[4][23] ) );
  NR2 U624 ( .A(n142), .B(n57), .Z(\ab[4][22] ) );
  NR2 U625 ( .A(n143), .B(n57), .Z(\ab[4][21] ) );
  NR2 U626 ( .A(n144), .B(n57), .Z(\ab[4][20] ) );
  NR2 U627 ( .A(n163), .B(n56), .Z(\ab[4][1] ) );
  NR2 U628 ( .A(n145), .B(n56), .Z(\ab[4][19] ) );
  NR2 U629 ( .A(n146), .B(n56), .Z(\ab[4][18] ) );
  NR2 U630 ( .A(n147), .B(n56), .Z(\ab[4][17] ) );
  NR2 U631 ( .A(n148), .B(n56), .Z(\ab[4][16] ) );
  NR2 U632 ( .A(n149), .B(n56), .Z(\ab[4][15] ) );
  NR2 U633 ( .A(n150), .B(n56), .Z(\ab[4][14] ) );
  NR2 U634 ( .A(n151), .B(n56), .Z(\ab[4][13] ) );
  NR2 U635 ( .A(n152), .B(n56), .Z(\ab[4][12] ) );
  NR2 U636 ( .A(n153), .B(n56), .Z(\ab[4][11] ) );
  NR2 U637 ( .A(n154), .B(n56), .Z(\ab[4][10] ) );
  NR2 U638 ( .A(n164), .B(n56), .Z(\ab[4][0] ) );
  NR2 U639 ( .A(n155), .B(n54), .Z(\ab[3][9] ) );
  NR2 U640 ( .A(n156), .B(n54), .Z(\ab[3][8] ) );
  NR2 U641 ( .A(n157), .B(n54), .Z(\ab[3][7] ) );
  NR2 U642 ( .A(n158), .B(n54), .Z(\ab[3][6] ) );
  NR2 U643 ( .A(n159), .B(n54), .Z(\ab[3][5] ) );
  NR2 U644 ( .A(n160), .B(n54), .Z(\ab[3][4] ) );
  NR2 U645 ( .A(n108), .B(n54), .Z(\ab[3][47] ) );
  NR2 U646 ( .A(n107), .B(n54), .Z(\ab[3][46] ) );
  NR2 U647 ( .A(n106), .B(n54), .Z(\ab[3][45] ) );
  NR2 U648 ( .A(n105), .B(n54), .Z(\ab[3][44] ) );
  NR2 U649 ( .A(n104), .B(n54), .Z(\ab[3][43] ) );
  NR2 U650 ( .A(n103), .B(n54), .Z(\ab[3][42] ) );
  NR2 U651 ( .A(n102), .B(n53), .Z(\ab[3][41] ) );
  NR2 U652 ( .A(n101), .B(n53), .Z(\ab[3][40] ) );
  NR2 U653 ( .A(n161), .B(n53), .Z(\ab[3][3] ) );
  NR2 U654 ( .A(n125), .B(n53), .Z(\ab[3][39] ) );
  NR2 U655 ( .A(n126), .B(n53), .Z(\ab[3][38] ) );
  NR2 U656 ( .A(n127), .B(n53), .Z(\ab[3][37] ) );
  NR2 U657 ( .A(n128), .B(n53), .Z(\ab[3][36] ) );
  NR2 U658 ( .A(n129), .B(n53), .Z(\ab[3][35] ) );
  NR2 U659 ( .A(n130), .B(n53), .Z(\ab[3][34] ) );
  NR2 U660 ( .A(n131), .B(n53), .Z(\ab[3][33] ) );
  NR2 U661 ( .A(n132), .B(n53), .Z(\ab[3][32] ) );
  NR2 U662 ( .A(n133), .B(n53), .Z(\ab[3][31] ) );
  NR2 U663 ( .A(n134), .B(n52), .Z(\ab[3][30] ) );
  NR2 U664 ( .A(n162), .B(n52), .Z(\ab[3][2] ) );
  NR2 U665 ( .A(n135), .B(n52), .Z(\ab[3][29] ) );
  NR2 U666 ( .A(n136), .B(n52), .Z(\ab[3][28] ) );
  NR2 U667 ( .A(n137), .B(n52), .Z(\ab[3][27] ) );
  NR2 U668 ( .A(n138), .B(n52), .Z(\ab[3][26] ) );
  NR2 U669 ( .A(n139), .B(n52), .Z(\ab[3][25] ) );
  NR2 U670 ( .A(n140), .B(n52), .Z(\ab[3][24] ) );
  NR2 U671 ( .A(n141), .B(n52), .Z(\ab[3][23] ) );
  NR2 U672 ( .A(n142), .B(n52), .Z(\ab[3][22] ) );
  NR2 U673 ( .A(n143), .B(n52), .Z(\ab[3][21] ) );
  NR2 U674 ( .A(n144), .B(n52), .Z(\ab[3][20] ) );
  NR2 U675 ( .A(n163), .B(n51), .Z(\ab[3][1] ) );
  NR2 U676 ( .A(n145), .B(n51), .Z(\ab[3][19] ) );
  NR2 U677 ( .A(n146), .B(n51), .Z(\ab[3][18] ) );
  NR2 U678 ( .A(n147), .B(n51), .Z(\ab[3][17] ) );
  NR2 U679 ( .A(n148), .B(n51), .Z(\ab[3][16] ) );
  NR2 U680 ( .A(n149), .B(n51), .Z(\ab[3][15] ) );
  NR2 U681 ( .A(n150), .B(n51), .Z(\ab[3][14] ) );
  NR2 U682 ( .A(n151), .B(n51), .Z(\ab[3][13] ) );
  NR2 U683 ( .A(n152), .B(n51), .Z(\ab[3][12] ) );
  NR2 U684 ( .A(n153), .B(n51), .Z(\ab[3][11] ) );
  NR2 U685 ( .A(n154), .B(n51), .Z(\ab[3][10] ) );
  NR2 U686 ( .A(n164), .B(n51), .Z(\ab[3][0] ) );
  NR2 U687 ( .A(n155), .B(n49), .Z(\ab[2][9] ) );
  NR2 U688 ( .A(n156), .B(n49), .Z(\ab[2][8] ) );
  NR2 U689 ( .A(n157), .B(n49), .Z(\ab[2][7] ) );
  NR2 U690 ( .A(n158), .B(n49), .Z(\ab[2][6] ) );
  NR2 U691 ( .A(n159), .B(n49), .Z(\ab[2][5] ) );
  NR2 U692 ( .A(n160), .B(n49), .Z(\ab[2][4] ) );
  NR2 U693 ( .A(n108), .B(n49), .Z(\ab[2][47] ) );
  NR2 U694 ( .A(n107), .B(n49), .Z(\ab[2][46] ) );
  NR2 U695 ( .A(n106), .B(n49), .Z(\ab[2][45] ) );
  NR2 U696 ( .A(n105), .B(n49), .Z(\ab[2][44] ) );
  NR2 U697 ( .A(n104), .B(n49), .Z(\ab[2][43] ) );
  NR2 U698 ( .A(n103), .B(n49), .Z(\ab[2][42] ) );
  NR2 U699 ( .A(n102), .B(n48), .Z(\ab[2][41] ) );
  NR2 U700 ( .A(n101), .B(n48), .Z(\ab[2][40] ) );
  NR2 U701 ( .A(n161), .B(n48), .Z(\ab[2][3] ) );
  NR2 U702 ( .A(n125), .B(n48), .Z(\ab[2][39] ) );
  NR2 U703 ( .A(n126), .B(n48), .Z(\ab[2][38] ) );
  NR2 U704 ( .A(n127), .B(n48), .Z(\ab[2][37] ) );
  NR2 U705 ( .A(n128), .B(n48), .Z(\ab[2][36] ) );
  NR2 U706 ( .A(n129), .B(n48), .Z(\ab[2][35] ) );
  NR2 U707 ( .A(n130), .B(n48), .Z(\ab[2][34] ) );
  NR2 U708 ( .A(n131), .B(n48), .Z(\ab[2][33] ) );
  NR2 U709 ( .A(n132), .B(n48), .Z(\ab[2][32] ) );
  NR2 U710 ( .A(n133), .B(n48), .Z(\ab[2][31] ) );
  NR2 U711 ( .A(n134), .B(n47), .Z(\ab[2][30] ) );
  NR2 U712 ( .A(n162), .B(n47), .Z(\ab[2][2] ) );
  NR2 U713 ( .A(n135), .B(n47), .Z(\ab[2][29] ) );
  NR2 U714 ( .A(n136), .B(n47), .Z(\ab[2][28] ) );
  NR2 U715 ( .A(n137), .B(n47), .Z(\ab[2][27] ) );
  NR2 U716 ( .A(n138), .B(n47), .Z(\ab[2][26] ) );
  NR2 U717 ( .A(n139), .B(n47), .Z(\ab[2][25] ) );
  NR2 U718 ( .A(n140), .B(n47), .Z(\ab[2][24] ) );
  NR2 U719 ( .A(n141), .B(n47), .Z(\ab[2][23] ) );
  NR2 U720 ( .A(n142), .B(n47), .Z(\ab[2][22] ) );
  NR2 U721 ( .A(n143), .B(n47), .Z(\ab[2][21] ) );
  NR2 U722 ( .A(n144), .B(n47), .Z(\ab[2][20] ) );
  NR2 U723 ( .A(n163), .B(n46), .Z(\ab[2][1] ) );
  NR2 U724 ( .A(n145), .B(n46), .Z(\ab[2][19] ) );
  NR2 U725 ( .A(n146), .B(n46), .Z(\ab[2][18] ) );
  NR2 U726 ( .A(n147), .B(n46), .Z(\ab[2][17] ) );
  NR2 U727 ( .A(n148), .B(n46), .Z(\ab[2][16] ) );
  NR2 U728 ( .A(n149), .B(n46), .Z(\ab[2][15] ) );
  NR2 U729 ( .A(n150), .B(n46), .Z(\ab[2][14] ) );
  NR2 U730 ( .A(n151), .B(n46), .Z(\ab[2][13] ) );
  NR2 U731 ( .A(n152), .B(n46), .Z(\ab[2][12] ) );
  NR2 U732 ( .A(n153), .B(n46), .Z(\ab[2][11] ) );
  NR2 U733 ( .A(n154), .B(n46), .Z(\ab[2][10] ) );
  NR2 U734 ( .A(n164), .B(n46), .Z(\ab[2][0] ) );
  NR2 U735 ( .A(n155), .B(n11), .Z(\ab[21][9] ) );
  NR2 U736 ( .A(n156), .B(n11), .Z(\ab[21][8] ) );
  NR2 U737 ( .A(n157), .B(n11), .Z(\ab[21][7] ) );
  NR2 U738 ( .A(n158), .B(n11), .Z(\ab[21][6] ) );
  NR2 U739 ( .A(n159), .B(n11), .Z(\ab[21][5] ) );
  NR2 U740 ( .A(n160), .B(n11), .Z(\ab[21][4] ) );
  NR2 U741 ( .A(n108), .B(n11), .Z(\ab[21][47] ) );
  NR2 U742 ( .A(n107), .B(n11), .Z(\ab[21][46] ) );
  NR2 U743 ( .A(n106), .B(n11), .Z(\ab[21][45] ) );
  NR2 U744 ( .A(n105), .B(n11), .Z(\ab[21][44] ) );
  NR2 U745 ( .A(n104), .B(n11), .Z(\ab[21][43] ) );
  NR2 U746 ( .A(n103), .B(n11), .Z(\ab[21][42] ) );
  NR2 U747 ( .A(n102), .B(n10), .Z(\ab[21][41] ) );
  NR2 U748 ( .A(n101), .B(n10), .Z(\ab[21][40] ) );
  NR2 U749 ( .A(n161), .B(n10), .Z(\ab[21][3] ) );
  NR2 U750 ( .A(n125), .B(n10), .Z(\ab[21][39] ) );
  NR2 U751 ( .A(n126), .B(n10), .Z(\ab[21][38] ) );
  NR2 U752 ( .A(n127), .B(n10), .Z(\ab[21][37] ) );
  NR2 U753 ( .A(n128), .B(n10), .Z(\ab[21][36] ) );
  NR2 U754 ( .A(n129), .B(n10), .Z(\ab[21][35] ) );
  NR2 U755 ( .A(n130), .B(n10), .Z(\ab[21][34] ) );
  NR2 U756 ( .A(n131), .B(n10), .Z(\ab[21][33] ) );
  NR2 U757 ( .A(n132), .B(n10), .Z(\ab[21][32] ) );
  NR2 U758 ( .A(n133), .B(n10), .Z(\ab[21][31] ) );
  NR2 U759 ( .A(n134), .B(n9), .Z(\ab[21][30] ) );
  NR2 U760 ( .A(n162), .B(n9), .Z(\ab[21][2] ) );
  NR2 U761 ( .A(n135), .B(n9), .Z(\ab[21][29] ) );
  NR2 U762 ( .A(n136), .B(n9), .Z(\ab[21][28] ) );
  NR2 U763 ( .A(n137), .B(n9), .Z(\ab[21][27] ) );
  NR2 U764 ( .A(n138), .B(n9), .Z(\ab[21][26] ) );
  NR2 U765 ( .A(n139), .B(n9), .Z(\ab[21][25] ) );
  NR2 U766 ( .A(n140), .B(n9), .Z(\ab[21][24] ) );
  NR2 U767 ( .A(n141), .B(n9), .Z(\ab[21][23] ) );
  NR2 U768 ( .A(n142), .B(n9), .Z(\ab[21][22] ) );
  NR2 U769 ( .A(n143), .B(n9), .Z(\ab[21][21] ) );
  NR2 U770 ( .A(n144), .B(n9), .Z(\ab[21][20] ) );
  NR2 U771 ( .A(n163), .B(n8), .Z(\ab[21][1] ) );
  NR2 U772 ( .A(n145), .B(n8), .Z(\ab[21][19] ) );
  NR2 U773 ( .A(n146), .B(n8), .Z(\ab[21][18] ) );
  NR2 U774 ( .A(n147), .B(n8), .Z(\ab[21][17] ) );
  NR2 U775 ( .A(n148), .B(n8), .Z(\ab[21][16] ) );
  NR2 U776 ( .A(n149), .B(n8), .Z(\ab[21][15] ) );
  NR2 U777 ( .A(n150), .B(n8), .Z(\ab[21][14] ) );
  NR2 U778 ( .A(n151), .B(n8), .Z(\ab[21][13] ) );
  NR2 U779 ( .A(n152), .B(n8), .Z(\ab[21][12] ) );
  NR2 U780 ( .A(n153), .B(n8), .Z(\ab[21][11] ) );
  NR2 U781 ( .A(n154), .B(n8), .Z(\ab[21][10] ) );
  NR2 U782 ( .A(n164), .B(n8), .Z(\ab[21][0] ) );
  NR2 U783 ( .A(n155), .B(n15), .Z(\ab[20][9] ) );
  NR2 U784 ( .A(n156), .B(n15), .Z(\ab[20][8] ) );
  NR2 U785 ( .A(n157), .B(n15), .Z(\ab[20][7] ) );
  NR2 U786 ( .A(n158), .B(n15), .Z(\ab[20][6] ) );
  NR2 U787 ( .A(n159), .B(n15), .Z(\ab[20][5] ) );
  NR2 U788 ( .A(n160), .B(n15), .Z(\ab[20][4] ) );
  NR2 U789 ( .A(n108), .B(n15), .Z(\ab[20][47] ) );
  NR2 U790 ( .A(n107), .B(n15), .Z(\ab[20][46] ) );
  NR2 U791 ( .A(n106), .B(n15), .Z(\ab[20][45] ) );
  NR2 U792 ( .A(n105), .B(n15), .Z(\ab[20][44] ) );
  NR2 U793 ( .A(n104), .B(n15), .Z(\ab[20][43] ) );
  NR2 U794 ( .A(n103), .B(n15), .Z(\ab[20][42] ) );
  NR2 U795 ( .A(n102), .B(n14), .Z(\ab[20][41] ) );
  NR2 U796 ( .A(n101), .B(n14), .Z(\ab[20][40] ) );
  NR2 U797 ( .A(n161), .B(n14), .Z(\ab[20][3] ) );
  NR2 U798 ( .A(n125), .B(n14), .Z(\ab[20][39] ) );
  NR2 U799 ( .A(n126), .B(n14), .Z(\ab[20][38] ) );
  NR2 U800 ( .A(n127), .B(n14), .Z(\ab[20][37] ) );
  NR2 U801 ( .A(n128), .B(n14), .Z(\ab[20][36] ) );
  NR2 U802 ( .A(n129), .B(n14), .Z(\ab[20][35] ) );
  NR2 U803 ( .A(n130), .B(n14), .Z(\ab[20][34] ) );
  NR2 U804 ( .A(n131), .B(n14), .Z(\ab[20][33] ) );
  NR2 U805 ( .A(n132), .B(n14), .Z(\ab[20][32] ) );
  NR2 U806 ( .A(n133), .B(n14), .Z(\ab[20][31] ) );
  NR2 U807 ( .A(n134), .B(n13), .Z(\ab[20][30] ) );
  NR2 U808 ( .A(n162), .B(n13), .Z(\ab[20][2] ) );
  NR2 U809 ( .A(n135), .B(n13), .Z(\ab[20][29] ) );
  NR2 U810 ( .A(n136), .B(n13), .Z(\ab[20][28] ) );
  NR2 U811 ( .A(n137), .B(n13), .Z(\ab[20][27] ) );
  NR2 U812 ( .A(n138), .B(n13), .Z(\ab[20][26] ) );
  NR2 U813 ( .A(n139), .B(n13), .Z(\ab[20][25] ) );
  NR2 U814 ( .A(n140), .B(n13), .Z(\ab[20][24] ) );
  NR2 U815 ( .A(n141), .B(n13), .Z(\ab[20][23] ) );
  NR2 U816 ( .A(n142), .B(n13), .Z(\ab[20][22] ) );
  NR2 U817 ( .A(n143), .B(n13), .Z(\ab[20][21] ) );
  NR2 U818 ( .A(n144), .B(n13), .Z(\ab[20][20] ) );
  NR2 U819 ( .A(n163), .B(n12), .Z(\ab[20][1] ) );
  NR2 U820 ( .A(n145), .B(n12), .Z(\ab[20][19] ) );
  NR2 U821 ( .A(n146), .B(n12), .Z(\ab[20][18] ) );
  NR2 U822 ( .A(n147), .B(n12), .Z(\ab[20][17] ) );
  NR2 U823 ( .A(n148), .B(n12), .Z(\ab[20][16] ) );
  NR2 U824 ( .A(n149), .B(n12), .Z(\ab[20][15] ) );
  NR2 U825 ( .A(n150), .B(n12), .Z(\ab[20][14] ) );
  NR2 U826 ( .A(n151), .B(n12), .Z(\ab[20][13] ) );
  NR2 U827 ( .A(n152), .B(n12), .Z(\ab[20][12] ) );
  NR2 U828 ( .A(n153), .B(n12), .Z(\ab[20][11] ) );
  NR2 U829 ( .A(n154), .B(n12), .Z(\ab[20][10] ) );
  NR2 U830 ( .A(n164), .B(n12), .Z(\ab[20][0] ) );
  NR2 U831 ( .A(n155), .B(n44), .Z(\ab[1][9] ) );
  NR2 U832 ( .A(n156), .B(n44), .Z(\ab[1][8] ) );
  NR2 U833 ( .A(n157), .B(n44), .Z(\ab[1][7] ) );
  NR2 U834 ( .A(n158), .B(n44), .Z(\ab[1][6] ) );
  NR2 U835 ( .A(n159), .B(n44), .Z(\ab[1][5] ) );
  NR2 U836 ( .A(n160), .B(n44), .Z(\ab[1][4] ) );
  NR2 U837 ( .A(n108), .B(n44), .Z(\ab[1][47] ) );
  NR2 U838 ( .A(n107), .B(n44), .Z(\ab[1][46] ) );
  NR2 U839 ( .A(n106), .B(n44), .Z(\ab[1][45] ) );
  NR2 U840 ( .A(n105), .B(n44), .Z(\ab[1][44] ) );
  NR2 U841 ( .A(n104), .B(n44), .Z(\ab[1][43] ) );
  NR2 U842 ( .A(n103), .B(n43), .Z(\ab[1][42] ) );
  NR2 U843 ( .A(n102), .B(n43), .Z(\ab[1][41] ) );
  NR2 U844 ( .A(n101), .B(n43), .Z(\ab[1][40] ) );
  NR2 U845 ( .A(n161), .B(n43), .Z(\ab[1][3] ) );
  NR2 U846 ( .A(n125), .B(n43), .Z(\ab[1][39] ) );
  NR2 U847 ( .A(n126), .B(n43), .Z(\ab[1][38] ) );
  NR2 U848 ( .A(n127), .B(n43), .Z(\ab[1][37] ) );
  NR2 U849 ( .A(n128), .B(n43), .Z(\ab[1][36] ) );
  NR2 U850 ( .A(n129), .B(n43), .Z(\ab[1][35] ) );
  NR2 U851 ( .A(n130), .B(n43), .Z(\ab[1][34] ) );
  NR2 U852 ( .A(n131), .B(n43), .Z(\ab[1][33] ) );
  NR2 U853 ( .A(n132), .B(n43), .Z(\ab[1][32] ) );
  NR2 U854 ( .A(n133), .B(n42), .Z(\ab[1][31] ) );
  NR2 U855 ( .A(n134), .B(n42), .Z(\ab[1][30] ) );
  NR2 U856 ( .A(n162), .B(n42), .Z(\ab[1][2] ) );
  NR2 U857 ( .A(n135), .B(n42), .Z(\ab[1][29] ) );
  NR2 U858 ( .A(n136), .B(n42), .Z(\ab[1][28] ) );
  NR2 U859 ( .A(n137), .B(n42), .Z(\ab[1][27] ) );
  NR2 U860 ( .A(n138), .B(n42), .Z(\ab[1][26] ) );
  NR2 U861 ( .A(n139), .B(n42), .Z(\ab[1][25] ) );
  NR2 U862 ( .A(n140), .B(n42), .Z(\ab[1][24] ) );
  NR2 U863 ( .A(n141), .B(n42), .Z(\ab[1][23] ) );
  NR2 U864 ( .A(n142), .B(n42), .Z(\ab[1][22] ) );
  NR2 U865 ( .A(n143), .B(n42), .Z(\ab[1][21] ) );
  NR2 U866 ( .A(n144), .B(n41), .Z(\ab[1][20] ) );
  NR2 U867 ( .A(n145), .B(n41), .Z(\ab[1][19] ) );
  NR2 U868 ( .A(n146), .B(n41), .Z(\ab[1][18] ) );
  NR2 U869 ( .A(n147), .B(n41), .Z(\ab[1][17] ) );
  NR2 U870 ( .A(n148), .B(n41), .Z(\ab[1][16] ) );
  NR2 U871 ( .A(n149), .B(n41), .Z(\ab[1][15] ) );
  NR2 U872 ( .A(n150), .B(n41), .Z(\ab[1][14] ) );
  NR2 U873 ( .A(n151), .B(n41), .Z(\ab[1][13] ) );
  NR2 U874 ( .A(n152), .B(n41), .Z(\ab[1][12] ) );
  NR2 U875 ( .A(n153), .B(n41), .Z(\ab[1][11] ) );
  NR2 U876 ( .A(n154), .B(n41), .Z(\ab[1][10] ) );
  NR2 U877 ( .A(n155), .B(n19), .Z(\ab[19][9] ) );
  NR2 U878 ( .A(n156), .B(n19), .Z(\ab[19][8] ) );
  NR2 U879 ( .A(n157), .B(n19), .Z(\ab[19][7] ) );
  NR2 U880 ( .A(n158), .B(n19), .Z(\ab[19][6] ) );
  NR2 U881 ( .A(n159), .B(n19), .Z(\ab[19][5] ) );
  NR2 U882 ( .A(n160), .B(n19), .Z(\ab[19][4] ) );
  NR2 U883 ( .A(n108), .B(n19), .Z(\ab[19][47] ) );
  NR2 U884 ( .A(n107), .B(n19), .Z(\ab[19][46] ) );
  NR2 U885 ( .A(n106), .B(n19), .Z(\ab[19][45] ) );
  NR2 U886 ( .A(n105), .B(n19), .Z(\ab[19][44] ) );
  NR2 U887 ( .A(n104), .B(n19), .Z(\ab[19][43] ) );
  NR2 U888 ( .A(n103), .B(n19), .Z(\ab[19][42] ) );
  NR2 U889 ( .A(n102), .B(n18), .Z(\ab[19][41] ) );
  NR2 U890 ( .A(n101), .B(n18), .Z(\ab[19][40] ) );
  NR2 U891 ( .A(n161), .B(n18), .Z(\ab[19][3] ) );
  NR2 U892 ( .A(n125), .B(n18), .Z(\ab[19][39] ) );
  NR2 U893 ( .A(n126), .B(n18), .Z(\ab[19][38] ) );
  NR2 U894 ( .A(n127), .B(n18), .Z(\ab[19][37] ) );
  NR2 U895 ( .A(n128), .B(n18), .Z(\ab[19][36] ) );
  NR2 U896 ( .A(n129), .B(n18), .Z(\ab[19][35] ) );
  NR2 U897 ( .A(n130), .B(n18), .Z(\ab[19][34] ) );
  NR2 U898 ( .A(n131), .B(n18), .Z(\ab[19][33] ) );
  NR2 U899 ( .A(n132), .B(n18), .Z(\ab[19][32] ) );
  NR2 U900 ( .A(n133), .B(n18), .Z(\ab[19][31] ) );
  NR2 U901 ( .A(n134), .B(n17), .Z(\ab[19][30] ) );
  NR2 U902 ( .A(n162), .B(n17), .Z(\ab[19][2] ) );
  NR2 U903 ( .A(n135), .B(n17), .Z(\ab[19][29] ) );
  NR2 U904 ( .A(n136), .B(n17), .Z(\ab[19][28] ) );
  NR2 U905 ( .A(n137), .B(n17), .Z(\ab[19][27] ) );
  NR2 U906 ( .A(n138), .B(n17), .Z(\ab[19][26] ) );
  NR2 U907 ( .A(n139), .B(n17), .Z(\ab[19][25] ) );
  NR2 U908 ( .A(n140), .B(n17), .Z(\ab[19][24] ) );
  NR2 U909 ( .A(n141), .B(n17), .Z(\ab[19][23] ) );
  NR2 U910 ( .A(n142), .B(n17), .Z(\ab[19][22] ) );
  NR2 U911 ( .A(n143), .B(n17), .Z(\ab[19][21] ) );
  NR2 U912 ( .A(n144), .B(n17), .Z(\ab[19][20] ) );
  NR2 U913 ( .A(n163), .B(n16), .Z(\ab[19][1] ) );
  NR2 U914 ( .A(n145), .B(n16), .Z(\ab[19][19] ) );
  NR2 U915 ( .A(n146), .B(n16), .Z(\ab[19][18] ) );
  NR2 U916 ( .A(n147), .B(n16), .Z(\ab[19][17] ) );
  NR2 U917 ( .A(n148), .B(n16), .Z(\ab[19][16] ) );
  NR2 U918 ( .A(n149), .B(n16), .Z(\ab[19][15] ) );
  NR2 U919 ( .A(n150), .B(n16), .Z(\ab[19][14] ) );
  NR2 U920 ( .A(n151), .B(n16), .Z(\ab[19][13] ) );
  NR2 U921 ( .A(n152), .B(n16), .Z(\ab[19][12] ) );
  NR2 U922 ( .A(n153), .B(n16), .Z(\ab[19][11] ) );
  NR2 U923 ( .A(n154), .B(n16), .Z(\ab[19][10] ) );
  NR2 U924 ( .A(n164), .B(n16), .Z(\ab[19][0] ) );
  NR2 U925 ( .A(n155), .B(n21), .Z(\ab[18][9] ) );
  NR2 U926 ( .A(n156), .B(n21), .Z(\ab[18][8] ) );
  NR2 U927 ( .A(n157), .B(n21), .Z(\ab[18][7] ) );
  NR2 U928 ( .A(n158), .B(n21), .Z(\ab[18][6] ) );
  NR2 U929 ( .A(n159), .B(n21), .Z(\ab[18][5] ) );
  NR2 U930 ( .A(n160), .B(n21), .Z(\ab[18][4] ) );
  NR2 U931 ( .A(n108), .B(n21), .Z(\ab[18][47] ) );
  NR2 U932 ( .A(n107), .B(n21), .Z(\ab[18][46] ) );
  NR2 U933 ( .A(n106), .B(n21), .Z(\ab[18][45] ) );
  NR2 U934 ( .A(n105), .B(n21), .Z(\ab[18][44] ) );
  NR2 U935 ( .A(n104), .B(n21), .Z(\ab[18][43] ) );
  NR2 U936 ( .A(n103), .B(n21), .Z(\ab[18][42] ) );
  NR2 U937 ( .A(n102), .B(n20), .Z(\ab[18][41] ) );
  NR2 U938 ( .A(n101), .B(n20), .Z(\ab[18][40] ) );
  NR2 U939 ( .A(n161), .B(n20), .Z(\ab[18][3] ) );
  NR2 U940 ( .A(n125), .B(n20), .Z(\ab[18][39] ) );
  NR2 U941 ( .A(n126), .B(n20), .Z(\ab[18][38] ) );
  NR2 U942 ( .A(n127), .B(n20), .Z(\ab[18][37] ) );
  NR2 U943 ( .A(n128), .B(n20), .Z(\ab[18][36] ) );
  NR2 U944 ( .A(n129), .B(n20), .Z(\ab[18][35] ) );
  NR2 U945 ( .A(n130), .B(n20), .Z(\ab[18][34] ) );
  NR2 U946 ( .A(n131), .B(n20), .Z(\ab[18][33] ) );
  NR2 U947 ( .A(n132), .B(n20), .Z(\ab[18][32] ) );
  NR2 U948 ( .A(n133), .B(n20), .Z(\ab[18][31] ) );
  NR2 U949 ( .A(n134), .B(n21), .Z(\ab[18][30] ) );
  NR2 U950 ( .A(n162), .B(n20), .Z(\ab[18][2] ) );
  NR2 U951 ( .A(n135), .B(n20), .Z(\ab[18][29] ) );
  NR2 U952 ( .A(n136), .B(n21), .Z(\ab[18][28] ) );
  NR2 U953 ( .A(n137), .B(n21), .Z(\ab[18][27] ) );
  NR2 U954 ( .A(n138), .B(n21), .Z(\ab[18][26] ) );
  NR2 U955 ( .A(n139), .B(n21), .Z(\ab[18][25] ) );
  NR2 U956 ( .A(n140), .B(n21), .Z(\ab[18][24] ) );
  NR2 U957 ( .A(n141), .B(n21), .Z(\ab[18][23] ) );
  NR2 U958 ( .A(n142), .B(n21), .Z(\ab[18][22] ) );
  NR2 U959 ( .A(n143), .B(n21), .Z(\ab[18][21] ) );
  NR2 U960 ( .A(n144), .B(n21), .Z(\ab[18][20] ) );
  NR2 U961 ( .A(n163), .B(n20), .Z(\ab[18][1] ) );
  NR2 U962 ( .A(n145), .B(n21), .Z(\ab[18][19] ) );
  NR2 U963 ( .A(n146), .B(n21), .Z(\ab[18][18] ) );
  NR2 U964 ( .A(n147), .B(n21), .Z(\ab[18][17] ) );
  NR2 U965 ( .A(n148), .B(n21), .Z(\ab[18][16] ) );
  NR2 U966 ( .A(n149), .B(n21), .Z(\ab[18][15] ) );
  NR2 U967 ( .A(n150), .B(n21), .Z(\ab[18][14] ) );
  NR2 U968 ( .A(n151), .B(n21), .Z(\ab[18][13] ) );
  NR2 U969 ( .A(n152), .B(n21), .Z(\ab[18][12] ) );
  NR2 U970 ( .A(n153), .B(n21), .Z(\ab[18][11] ) );
  NR2 U971 ( .A(n154), .B(n21), .Z(\ab[18][10] ) );
  NR2 U972 ( .A(n164), .B(n21), .Z(\ab[18][0] ) );
  NR2 U973 ( .A(n155), .B(n22), .Z(\ab[17][9] ) );
  NR2 U974 ( .A(n156), .B(n22), .Z(\ab[17][8] ) );
  NR2 U975 ( .A(n157), .B(n22), .Z(\ab[17][7] ) );
  NR2 U976 ( .A(n158), .B(n22), .Z(\ab[17][6] ) );
  NR2 U977 ( .A(n159), .B(n22), .Z(\ab[17][5] ) );
  NR2 U978 ( .A(n160), .B(n22), .Z(\ab[17][4] ) );
  NR2 U979 ( .A(n108), .B(n22), .Z(\ab[17][47] ) );
  NR2 U980 ( .A(n107), .B(n22), .Z(\ab[17][46] ) );
  NR2 U981 ( .A(n106), .B(n22), .Z(\ab[17][45] ) );
  NR2 U982 ( .A(n105), .B(n22), .Z(\ab[17][44] ) );
  NR2 U983 ( .A(n104), .B(n22), .Z(\ab[17][43] ) );
  NR2 U984 ( .A(n103), .B(n22), .Z(\ab[17][42] ) );
  NR2 U985 ( .A(n102), .B(n22), .Z(\ab[17][41] ) );
  NR2 U986 ( .A(n101), .B(n22), .Z(\ab[17][40] ) );
  NR2 U987 ( .A(n161), .B(n22), .Z(\ab[17][3] ) );
  NR2 U988 ( .A(n125), .B(n22), .Z(\ab[17][39] ) );
  NR2 U989 ( .A(n126), .B(n22), .Z(\ab[17][38] ) );
  NR2 U990 ( .A(n127), .B(n22), .Z(\ab[17][37] ) );
  NR2 U991 ( .A(n128), .B(n22), .Z(\ab[17][36] ) );
  NR2 U992 ( .A(n129), .B(n22), .Z(\ab[17][35] ) );
  NR2 U993 ( .A(n130), .B(n22), .Z(\ab[17][34] ) );
  NR2 U994 ( .A(n131), .B(n22), .Z(\ab[17][33] ) );
  NR2 U995 ( .A(n132), .B(n22), .Z(\ab[17][32] ) );
  NR2 U996 ( .A(n133), .B(n22), .Z(\ab[17][31] ) );
  NR2 U997 ( .A(n134), .B(n22), .Z(\ab[17][30] ) );
  NR2 U998 ( .A(n162), .B(n22), .Z(\ab[17][2] ) );
  NR2 U999 ( .A(n135), .B(n22), .Z(\ab[17][29] ) );
  NR2 U1000 ( .A(n136), .B(n22), .Z(\ab[17][28] ) );
  NR2 U1001 ( .A(n137), .B(n22), .Z(\ab[17][27] ) );
  NR2 U1002 ( .A(n138), .B(n22), .Z(\ab[17][26] ) );
  NR2 U1003 ( .A(n139), .B(n22), .Z(\ab[17][25] ) );
  NR2 U1004 ( .A(n140), .B(n22), .Z(\ab[17][24] ) );
  NR2 U1005 ( .A(n141), .B(n22), .Z(\ab[17][23] ) );
  NR2 U1006 ( .A(n142), .B(n22), .Z(\ab[17][22] ) );
  NR2 U1007 ( .A(n143), .B(n22), .Z(\ab[17][21] ) );
  NR2 U1008 ( .A(n144), .B(n22), .Z(\ab[17][20] ) );
  NR2 U1009 ( .A(n163), .B(n22), .Z(\ab[17][1] ) );
  NR2 U1010 ( .A(n145), .B(n22), .Z(\ab[17][19] ) );
  NR2 U1011 ( .A(n146), .B(n22), .Z(\ab[17][18] ) );
  NR2 U1012 ( .A(n147), .B(n22), .Z(\ab[17][17] ) );
  NR2 U1013 ( .A(n148), .B(n22), .Z(\ab[17][16] ) );
  NR2 U1014 ( .A(n149), .B(n22), .Z(\ab[17][15] ) );
  NR2 U1015 ( .A(n150), .B(n22), .Z(\ab[17][14] ) );
  NR2 U1016 ( .A(n151), .B(n22), .Z(\ab[17][13] ) );
  NR2 U1017 ( .A(n152), .B(n22), .Z(\ab[17][12] ) );
  NR2 U1018 ( .A(n153), .B(n22), .Z(\ab[17][11] ) );
  NR2 U1019 ( .A(n154), .B(n22), .Z(\ab[17][10] ) );
  NR2 U1020 ( .A(n164), .B(n22), .Z(\ab[17][0] ) );
  NR2 U1021 ( .A(n155), .B(n25), .Z(\ab[16][9] ) );
  NR2 U1022 ( .A(n156), .B(n25), .Z(\ab[16][8] ) );
  NR2 U1023 ( .A(n157), .B(n25), .Z(\ab[16][7] ) );
  NR2 U1024 ( .A(n158), .B(n25), .Z(\ab[16][6] ) );
  NR2 U1025 ( .A(n159), .B(n25), .Z(\ab[16][5] ) );
  NR2 U1026 ( .A(n160), .B(n25), .Z(\ab[16][4] ) );
  NR2 U1027 ( .A(n108), .B(n25), .Z(\ab[16][47] ) );
  NR2 U1028 ( .A(n107), .B(n25), .Z(\ab[16][46] ) );
  NR2 U1029 ( .A(n106), .B(n25), .Z(\ab[16][45] ) );
  NR2 U1030 ( .A(n105), .B(n25), .Z(\ab[16][44] ) );
  NR2 U1031 ( .A(n104), .B(n25), .Z(\ab[16][43] ) );
  NR2 U1032 ( .A(n103), .B(n25), .Z(\ab[16][42] ) );
  NR2 U1033 ( .A(n102), .B(n24), .Z(\ab[16][41] ) );
  NR2 U1034 ( .A(n101), .B(n24), .Z(\ab[16][40] ) );
  NR2 U1035 ( .A(n161), .B(n24), .Z(\ab[16][3] ) );
  NR2 U1036 ( .A(n125), .B(n24), .Z(\ab[16][39] ) );
  NR2 U1037 ( .A(n126), .B(n24), .Z(\ab[16][38] ) );
  NR2 U1038 ( .A(n127), .B(n24), .Z(\ab[16][37] ) );
  NR2 U1039 ( .A(n128), .B(n24), .Z(\ab[16][36] ) );
  NR2 U1040 ( .A(n129), .B(n24), .Z(\ab[16][35] ) );
  NR2 U1041 ( .A(n130), .B(n24), .Z(\ab[16][34] ) );
  NR2 U1042 ( .A(n131), .B(n24), .Z(\ab[16][33] ) );
  NR2 U1043 ( .A(n132), .B(n24), .Z(\ab[16][32] ) );
  NR2 U1044 ( .A(n133), .B(n24), .Z(\ab[16][31] ) );
  NR2 U1045 ( .A(n134), .B(n25), .Z(\ab[16][30] ) );
  NR2 U1046 ( .A(n162), .B(n23), .Z(\ab[16][2] ) );
  NR2 U1047 ( .A(n135), .B(n25), .Z(\ab[16][29] ) );
  NR2 U1048 ( .A(n136), .B(n25), .Z(\ab[16][28] ) );
  NR2 U1049 ( .A(n137), .B(n25), .Z(\ab[16][27] ) );
  NR2 U1050 ( .A(n138), .B(n25), .Z(\ab[16][26] ) );
  NR2 U1051 ( .A(n139), .B(n25), .Z(\ab[16][25] ) );
  NR2 U1052 ( .A(n140), .B(n25), .Z(\ab[16][24] ) );
  NR2 U1053 ( .A(n141), .B(n25), .Z(\ab[16][23] ) );
  NR2 U1054 ( .A(n142), .B(n25), .Z(\ab[16][22] ) );
  NR2 U1055 ( .A(n143), .B(n25), .Z(\ab[16][21] ) );
  NR2 U1056 ( .A(n144), .B(n25), .Z(\ab[16][20] ) );
  NR2 U1057 ( .A(n163), .B(n23), .Z(\ab[16][1] ) );
  NR2 U1058 ( .A(n145), .B(n23), .Z(\ab[16][19] ) );
  NR2 U1059 ( .A(n146), .B(n23), .Z(\ab[16][18] ) );
  NR2 U1060 ( .A(n147), .B(n23), .Z(\ab[16][17] ) );
  NR2 U1061 ( .A(n148), .B(n23), .Z(\ab[16][16] ) );
  NR2 U1062 ( .A(n149), .B(n23), .Z(\ab[16][15] ) );
  NR2 U1063 ( .A(n150), .B(n23), .Z(\ab[16][14] ) );
  NR2 U1064 ( .A(n151), .B(n23), .Z(\ab[16][13] ) );
  NR2 U1065 ( .A(n152), .B(n23), .Z(\ab[16][12] ) );
  NR2 U1066 ( .A(n153), .B(n23), .Z(\ab[16][11] ) );
  NR2 U1067 ( .A(n154), .B(n23), .Z(\ab[16][10] ) );
  NR2 U1068 ( .A(n164), .B(n23), .Z(\ab[16][0] ) );
  NR2 U1069 ( .A(n155), .B(n29), .Z(\ab[15][9] ) );
  NR2 U1070 ( .A(n156), .B(n29), .Z(\ab[15][8] ) );
  NR2 U1071 ( .A(n157), .B(n29), .Z(\ab[15][7] ) );
  NR2 U1072 ( .A(n158), .B(n29), .Z(\ab[15][6] ) );
  NR2 U1073 ( .A(n159), .B(n29), .Z(\ab[15][5] ) );
  NR2 U1074 ( .A(n160), .B(n29), .Z(\ab[15][4] ) );
  NR2 U1075 ( .A(n108), .B(n29), .Z(\ab[15][47] ) );
  NR2 U1076 ( .A(n107), .B(n29), .Z(\ab[15][46] ) );
  NR2 U1077 ( .A(n106), .B(n29), .Z(\ab[15][45] ) );
  NR2 U1078 ( .A(n105), .B(n29), .Z(\ab[15][44] ) );
  NR2 U1079 ( .A(n104), .B(n29), .Z(\ab[15][43] ) );
  NR2 U1080 ( .A(n103), .B(n29), .Z(\ab[15][42] ) );
  NR2 U1081 ( .A(n102), .B(n28), .Z(\ab[15][41] ) );
  NR2 U1082 ( .A(n101), .B(n28), .Z(\ab[15][40] ) );
  NR2 U1083 ( .A(n161), .B(n28), .Z(\ab[15][3] ) );
  NR2 U1084 ( .A(n125), .B(n28), .Z(\ab[15][39] ) );
  NR2 U1085 ( .A(n126), .B(n28), .Z(\ab[15][38] ) );
  NR2 U1086 ( .A(n127), .B(n28), .Z(\ab[15][37] ) );
  NR2 U1087 ( .A(n128), .B(n28), .Z(\ab[15][36] ) );
  NR2 U1088 ( .A(n129), .B(n28), .Z(\ab[15][35] ) );
  NR2 U1089 ( .A(n130), .B(n28), .Z(\ab[15][34] ) );
  NR2 U1090 ( .A(n131), .B(n28), .Z(\ab[15][33] ) );
  NR2 U1091 ( .A(n132), .B(n28), .Z(\ab[15][32] ) );
  NR2 U1092 ( .A(n133), .B(n28), .Z(\ab[15][31] ) );
  NR2 U1093 ( .A(n134), .B(n27), .Z(\ab[15][30] ) );
  NR2 U1094 ( .A(n162), .B(n27), .Z(\ab[15][2] ) );
  NR2 U1095 ( .A(n135), .B(n27), .Z(\ab[15][29] ) );
  NR2 U1096 ( .A(n136), .B(n27), .Z(\ab[15][28] ) );
  NR2 U1097 ( .A(n137), .B(n27), .Z(\ab[15][27] ) );
  NR2 U1098 ( .A(n138), .B(n27), .Z(\ab[15][26] ) );
  NR2 U1099 ( .A(n139), .B(n27), .Z(\ab[15][25] ) );
  NR2 U1100 ( .A(n140), .B(n27), .Z(\ab[15][24] ) );
  NR2 U1101 ( .A(n141), .B(n27), .Z(\ab[15][23] ) );
  NR2 U1102 ( .A(n142), .B(n27), .Z(\ab[15][22] ) );
  NR2 U1103 ( .A(n143), .B(n27), .Z(\ab[15][21] ) );
  NR2 U1104 ( .A(n144), .B(n27), .Z(\ab[15][20] ) );
  NR2 U1105 ( .A(n163), .B(n26), .Z(\ab[15][1] ) );
  NR2 U1106 ( .A(n145), .B(n26), .Z(\ab[15][19] ) );
  NR2 U1107 ( .A(n146), .B(n26), .Z(\ab[15][18] ) );
  NR2 U1108 ( .A(n147), .B(n26), .Z(\ab[15][17] ) );
  NR2 U1109 ( .A(n148), .B(n26), .Z(\ab[15][16] ) );
  NR2 U1110 ( .A(n149), .B(n26), .Z(\ab[15][15] ) );
  NR2 U1111 ( .A(n150), .B(n26), .Z(\ab[15][14] ) );
  NR2 U1112 ( .A(n151), .B(n26), .Z(\ab[15][13] ) );
  NR2 U1113 ( .A(n152), .B(n26), .Z(\ab[15][12] ) );
  NR2 U1114 ( .A(n153), .B(n26), .Z(\ab[15][11] ) );
  NR2 U1115 ( .A(n154), .B(n26), .Z(\ab[15][10] ) );
  NR2 U1116 ( .A(n164), .B(n26), .Z(\ab[15][0] ) );
  NR2 U1117 ( .A(n155), .B(n6), .Z(\ab[14][9] ) );
  NR2 U1118 ( .A(n156), .B(n6), .Z(\ab[14][8] ) );
  NR2 U1119 ( .A(n157), .B(n6), .Z(\ab[14][7] ) );
  NR2 U1120 ( .A(n158), .B(n6), .Z(\ab[14][6] ) );
  NR2 U1121 ( .A(n159), .B(n6), .Z(\ab[14][5] ) );
  NR2 U1122 ( .A(n160), .B(n6), .Z(\ab[14][4] ) );
  NR2 U1123 ( .A(n108), .B(n6), .Z(\ab[14][47] ) );
  NR2 U1124 ( .A(n107), .B(n6), .Z(\ab[14][46] ) );
  NR2 U1125 ( .A(n106), .B(n6), .Z(\ab[14][45] ) );
  NR2 U1126 ( .A(n105), .B(n6), .Z(\ab[14][44] ) );
  NR2 U1127 ( .A(n104), .B(n6), .Z(\ab[14][43] ) );
  NR2 U1128 ( .A(n103), .B(n6), .Z(\ab[14][42] ) );
  NR2 U1129 ( .A(n102), .B(n5), .Z(\ab[14][41] ) );
  NR2 U1130 ( .A(n101), .B(n5), .Z(\ab[14][40] ) );
  NR2 U1131 ( .A(n161), .B(n5), .Z(\ab[14][3] ) );
  NR2 U1132 ( .A(n125), .B(n5), .Z(\ab[14][39] ) );
  NR2 U1133 ( .A(n126), .B(n5), .Z(\ab[14][38] ) );
  NR2 U1134 ( .A(n127), .B(n5), .Z(\ab[14][37] ) );
  NR2 U1135 ( .A(n128), .B(n5), .Z(\ab[14][36] ) );
  NR2 U1136 ( .A(n129), .B(n5), .Z(\ab[14][35] ) );
  NR2 U1137 ( .A(n130), .B(n5), .Z(\ab[14][34] ) );
  NR2 U1138 ( .A(n131), .B(n5), .Z(\ab[14][33] ) );
  NR2 U1139 ( .A(n132), .B(n5), .Z(\ab[14][32] ) );
  NR2 U1140 ( .A(n133), .B(n5), .Z(\ab[14][31] ) );
  NR2 U1141 ( .A(n134), .B(n4), .Z(\ab[14][30] ) );
  NR2 U1142 ( .A(n162), .B(n4), .Z(\ab[14][2] ) );
  NR2 U1143 ( .A(n135), .B(n4), .Z(\ab[14][29] ) );
  NR2 U1144 ( .A(n136), .B(n4), .Z(\ab[14][28] ) );
  NR2 U1145 ( .A(n137), .B(n4), .Z(\ab[14][27] ) );
  NR2 U1146 ( .A(n138), .B(n4), .Z(\ab[14][26] ) );
  NR2 U1147 ( .A(n139), .B(n4), .Z(\ab[14][25] ) );
  NR2 U1148 ( .A(n140), .B(n4), .Z(\ab[14][24] ) );
  NR2 U1149 ( .A(n141), .B(n4), .Z(\ab[14][23] ) );
  NR2 U1150 ( .A(n142), .B(n4), .Z(\ab[14][22] ) );
  NR2 U1151 ( .A(n143), .B(n4), .Z(\ab[14][21] ) );
  NR2 U1152 ( .A(n144), .B(n4), .Z(\ab[14][20] ) );
  NR2 U1153 ( .A(n163), .B(n3), .Z(\ab[14][1] ) );
  NR2 U1154 ( .A(n145), .B(n3), .Z(\ab[14][19] ) );
  NR2 U1155 ( .A(n146), .B(n3), .Z(\ab[14][18] ) );
  NR2 U1156 ( .A(n147), .B(n3), .Z(\ab[14][17] ) );
  NR2 U1157 ( .A(n148), .B(n3), .Z(\ab[14][16] ) );
  NR2 U1158 ( .A(n149), .B(n3), .Z(\ab[14][15] ) );
  NR2 U1159 ( .A(n150), .B(n3), .Z(\ab[14][14] ) );
  NR2 U1160 ( .A(n151), .B(n3), .Z(\ab[14][13] ) );
  NR2 U1161 ( .A(n152), .B(n3), .Z(\ab[14][12] ) );
  NR2 U1162 ( .A(n153), .B(n3), .Z(\ab[14][11] ) );
  NR2 U1163 ( .A(n154), .B(n3), .Z(\ab[14][10] ) );
  NR2 U1164 ( .A(n164), .B(n3), .Z(\ab[14][0] ) );
  NR2 U1165 ( .A(n155), .B(n34), .Z(\ab[13][9] ) );
  NR2 U1166 ( .A(n156), .B(n34), .Z(\ab[13][8] ) );
  NR2 U1167 ( .A(n157), .B(n34), .Z(\ab[13][7] ) );
  NR2 U1168 ( .A(n158), .B(n34), .Z(\ab[13][6] ) );
  NR2 U1169 ( .A(n159), .B(n34), .Z(\ab[13][5] ) );
  NR2 U1170 ( .A(n160), .B(n34), .Z(\ab[13][4] ) );
  NR2 U1171 ( .A(n108), .B(n34), .Z(\ab[13][47] ) );
  NR2 U1172 ( .A(n107), .B(n34), .Z(\ab[13][46] ) );
  NR2 U1173 ( .A(n106), .B(n34), .Z(\ab[13][45] ) );
  NR2 U1174 ( .A(n105), .B(n34), .Z(\ab[13][44] ) );
  NR2 U1175 ( .A(n104), .B(n34), .Z(\ab[13][43] ) );
  NR2 U1176 ( .A(n103), .B(n34), .Z(\ab[13][42] ) );
  NR2 U1177 ( .A(n102), .B(n33), .Z(\ab[13][41] ) );
  NR2 U1178 ( .A(n101), .B(n33), .Z(\ab[13][40] ) );
  NR2 U1179 ( .A(n161), .B(n33), .Z(\ab[13][3] ) );
  NR2 U1180 ( .A(n125), .B(n33), .Z(\ab[13][39] ) );
  NR2 U1181 ( .A(n126), .B(n33), .Z(\ab[13][38] ) );
  NR2 U1182 ( .A(n127), .B(n33), .Z(\ab[13][37] ) );
  NR2 U1183 ( .A(n128), .B(n33), .Z(\ab[13][36] ) );
  NR2 U1184 ( .A(n129), .B(n33), .Z(\ab[13][35] ) );
  NR2 U1185 ( .A(n130), .B(n33), .Z(\ab[13][34] ) );
  NR2 U1186 ( .A(n131), .B(n33), .Z(\ab[13][33] ) );
  NR2 U1187 ( .A(n132), .B(n33), .Z(\ab[13][32] ) );
  NR2 U1188 ( .A(n133), .B(n33), .Z(\ab[13][31] ) );
  NR2 U1189 ( .A(n134), .B(n32), .Z(\ab[13][30] ) );
  NR2 U1190 ( .A(n162), .B(n32), .Z(\ab[13][2] ) );
  NR2 U1191 ( .A(n135), .B(n32), .Z(\ab[13][29] ) );
  NR2 U1192 ( .A(n136), .B(n32), .Z(\ab[13][28] ) );
  NR2 U1193 ( .A(n137), .B(n32), .Z(\ab[13][27] ) );
  NR2 U1194 ( .A(n138), .B(n32), .Z(\ab[13][26] ) );
  NR2 U1195 ( .A(n139), .B(n32), .Z(\ab[13][25] ) );
  NR2 U1196 ( .A(n140), .B(n32), .Z(\ab[13][24] ) );
  NR2 U1197 ( .A(n141), .B(n32), .Z(\ab[13][23] ) );
  NR2 U1198 ( .A(n142), .B(n32), .Z(\ab[13][22] ) );
  NR2 U1199 ( .A(n143), .B(n32), .Z(\ab[13][21] ) );
  NR2 U1200 ( .A(n144), .B(n32), .Z(\ab[13][20] ) );
  NR2 U1201 ( .A(n163), .B(n31), .Z(\ab[13][1] ) );
  NR2 U1202 ( .A(n145), .B(n31), .Z(\ab[13][19] ) );
  NR2 U1203 ( .A(n146), .B(n31), .Z(\ab[13][18] ) );
  NR2 U1204 ( .A(n147), .B(n31), .Z(\ab[13][17] ) );
  NR2 U1205 ( .A(n148), .B(n31), .Z(\ab[13][16] ) );
  NR2 U1206 ( .A(n149), .B(n31), .Z(\ab[13][15] ) );
  NR2 U1207 ( .A(n150), .B(n31), .Z(\ab[13][14] ) );
  NR2 U1208 ( .A(n151), .B(n31), .Z(\ab[13][13] ) );
  NR2 U1209 ( .A(n152), .B(n31), .Z(\ab[13][12] ) );
  NR2 U1210 ( .A(n153), .B(n31), .Z(\ab[13][11] ) );
  NR2 U1211 ( .A(n154), .B(n31), .Z(\ab[13][10] ) );
  NR2 U1212 ( .A(n164), .B(n31), .Z(\ab[13][0] ) );
  NR2 U1213 ( .A(n155), .B(n99), .Z(\ab[12][9] ) );
  NR2 U1214 ( .A(n156), .B(n99), .Z(\ab[12][8] ) );
  NR2 U1215 ( .A(n157), .B(n99), .Z(\ab[12][7] ) );
  NR2 U1216 ( .A(n158), .B(n99), .Z(\ab[12][6] ) );
  NR2 U1217 ( .A(n159), .B(n99), .Z(\ab[12][5] ) );
  NR2 U1218 ( .A(n160), .B(n99), .Z(\ab[12][4] ) );
  NR2 U1219 ( .A(n108), .B(n99), .Z(\ab[12][47] ) );
  NR2 U1220 ( .A(n107), .B(n99), .Z(\ab[12][46] ) );
  NR2 U1221 ( .A(n106), .B(n99), .Z(\ab[12][45] ) );
  NR2 U1222 ( .A(n105), .B(n99), .Z(\ab[12][44] ) );
  NR2 U1223 ( .A(n104), .B(n99), .Z(\ab[12][43] ) );
  NR2 U1224 ( .A(n103), .B(n99), .Z(\ab[12][42] ) );
  NR2 U1225 ( .A(n102), .B(n98), .Z(\ab[12][41] ) );
  NR2 U1226 ( .A(n101), .B(n98), .Z(\ab[12][40] ) );
  NR2 U1227 ( .A(n161), .B(n98), .Z(\ab[12][3] ) );
  NR2 U1228 ( .A(n125), .B(n98), .Z(\ab[12][39] ) );
  NR2 U1229 ( .A(n126), .B(n98), .Z(\ab[12][38] ) );
  NR2 U1230 ( .A(n127), .B(n98), .Z(\ab[12][37] ) );
  NR2 U1231 ( .A(n128), .B(n98), .Z(\ab[12][36] ) );
  NR2 U1232 ( .A(n129), .B(n98), .Z(\ab[12][35] ) );
  NR2 U1233 ( .A(n130), .B(n98), .Z(\ab[12][34] ) );
  NR2 U1234 ( .A(n131), .B(n98), .Z(\ab[12][33] ) );
  NR2 U1235 ( .A(n132), .B(n98), .Z(\ab[12][32] ) );
  NR2 U1236 ( .A(n133), .B(n98), .Z(\ab[12][31] ) );
  NR2 U1237 ( .A(n134), .B(n97), .Z(\ab[12][30] ) );
  NR2 U1238 ( .A(n162), .B(n97), .Z(\ab[12][2] ) );
  NR2 U1239 ( .A(n135), .B(n97), .Z(\ab[12][29] ) );
  NR2 U1240 ( .A(n136), .B(n97), .Z(\ab[12][28] ) );
  NR2 U1241 ( .A(n137), .B(n97), .Z(\ab[12][27] ) );
  NR2 U1242 ( .A(n138), .B(n97), .Z(\ab[12][26] ) );
  NR2 U1243 ( .A(n139), .B(n97), .Z(\ab[12][25] ) );
  NR2 U1244 ( .A(n140), .B(n97), .Z(\ab[12][24] ) );
  NR2 U1245 ( .A(n141), .B(n97), .Z(\ab[12][23] ) );
  NR2 U1246 ( .A(n142), .B(n97), .Z(\ab[12][22] ) );
  NR2 U1247 ( .A(n143), .B(n97), .Z(\ab[12][21] ) );
  NR2 U1248 ( .A(n144), .B(n97), .Z(\ab[12][20] ) );
  NR2 U1249 ( .A(n163), .B(n96), .Z(\ab[12][1] ) );
  NR2 U1250 ( .A(n145), .B(n96), .Z(\ab[12][19] ) );
  NR2 U1251 ( .A(n146), .B(n96), .Z(\ab[12][18] ) );
  NR2 U1252 ( .A(n147), .B(n96), .Z(\ab[12][17] ) );
  NR2 U1253 ( .A(n148), .B(n96), .Z(\ab[12][16] ) );
  NR2 U1254 ( .A(n149), .B(n96), .Z(\ab[12][15] ) );
  NR2 U1255 ( .A(n150), .B(n96), .Z(\ab[12][14] ) );
  NR2 U1256 ( .A(n151), .B(n96), .Z(\ab[12][13] ) );
  NR2 U1257 ( .A(n152), .B(n96), .Z(\ab[12][12] ) );
  NR2 U1258 ( .A(n153), .B(n96), .Z(\ab[12][11] ) );
  NR2 U1259 ( .A(n154), .B(n96), .Z(\ab[12][10] ) );
  NR2 U1260 ( .A(n164), .B(n96), .Z(\ab[12][0] ) );
  NR2 U1261 ( .A(n155), .B(n94), .Z(\ab[11][9] ) );
  NR2 U1262 ( .A(n156), .B(n94), .Z(\ab[11][8] ) );
  NR2 U1263 ( .A(n157), .B(n94), .Z(\ab[11][7] ) );
  NR2 U1264 ( .A(n158), .B(n94), .Z(\ab[11][6] ) );
  NR2 U1265 ( .A(n159), .B(n94), .Z(\ab[11][5] ) );
  NR2 U1266 ( .A(n160), .B(n94), .Z(\ab[11][4] ) );
  NR2 U1267 ( .A(n108), .B(n94), .Z(\ab[11][47] ) );
  NR2 U1268 ( .A(n107), .B(n94), .Z(\ab[11][46] ) );
  NR2 U1269 ( .A(n106), .B(n94), .Z(\ab[11][45] ) );
  NR2 U1270 ( .A(n105), .B(n94), .Z(\ab[11][44] ) );
  NR2 U1271 ( .A(n104), .B(n94), .Z(\ab[11][43] ) );
  NR2 U1272 ( .A(n103), .B(n94), .Z(\ab[11][42] ) );
  NR2 U1273 ( .A(n102), .B(n93), .Z(\ab[11][41] ) );
  NR2 U1274 ( .A(n101), .B(n93), .Z(\ab[11][40] ) );
  NR2 U1275 ( .A(n161), .B(n93), .Z(\ab[11][3] ) );
  NR2 U1276 ( .A(n125), .B(n93), .Z(\ab[11][39] ) );
  NR2 U1277 ( .A(n126), .B(n93), .Z(\ab[11][38] ) );
  NR2 U1278 ( .A(n127), .B(n93), .Z(\ab[11][37] ) );
  NR2 U1279 ( .A(n128), .B(n93), .Z(\ab[11][36] ) );
  NR2 U1280 ( .A(n129), .B(n93), .Z(\ab[11][35] ) );
  NR2 U1281 ( .A(n130), .B(n93), .Z(\ab[11][34] ) );
  NR2 U1282 ( .A(n131), .B(n93), .Z(\ab[11][33] ) );
  NR2 U1283 ( .A(n132), .B(n93), .Z(\ab[11][32] ) );
  NR2 U1284 ( .A(n133), .B(n93), .Z(\ab[11][31] ) );
  NR2 U1285 ( .A(n134), .B(n92), .Z(\ab[11][30] ) );
  NR2 U1286 ( .A(n162), .B(n92), .Z(\ab[11][2] ) );
  NR2 U1287 ( .A(n135), .B(n92), .Z(\ab[11][29] ) );
  NR2 U1288 ( .A(n136), .B(n92), .Z(\ab[11][28] ) );
  NR2 U1289 ( .A(n137), .B(n92), .Z(\ab[11][27] ) );
  NR2 U1290 ( .A(n138), .B(n92), .Z(\ab[11][26] ) );
  NR2 U1291 ( .A(n139), .B(n92), .Z(\ab[11][25] ) );
  NR2 U1292 ( .A(n140), .B(n92), .Z(\ab[11][24] ) );
  NR2 U1293 ( .A(n141), .B(n92), .Z(\ab[11][23] ) );
  NR2 U1294 ( .A(n142), .B(n92), .Z(\ab[11][22] ) );
  NR2 U1295 ( .A(n143), .B(n92), .Z(\ab[11][21] ) );
  NR2 U1296 ( .A(n144), .B(n92), .Z(\ab[11][20] ) );
  NR2 U1297 ( .A(n163), .B(n91), .Z(\ab[11][1] ) );
  NR2 U1298 ( .A(n145), .B(n91), .Z(\ab[11][19] ) );
  NR2 U1299 ( .A(n146), .B(n91), .Z(\ab[11][18] ) );
  NR2 U1300 ( .A(n147), .B(n91), .Z(\ab[11][17] ) );
  NR2 U1301 ( .A(n148), .B(n91), .Z(\ab[11][16] ) );
  NR2 U1302 ( .A(n149), .B(n91), .Z(\ab[11][15] ) );
  NR2 U1303 ( .A(n150), .B(n91), .Z(\ab[11][14] ) );
  NR2 U1304 ( .A(n151), .B(n91), .Z(\ab[11][13] ) );
  NR2 U1305 ( .A(n152), .B(n91), .Z(\ab[11][12] ) );
  NR2 U1306 ( .A(n153), .B(n91), .Z(\ab[11][11] ) );
  NR2 U1307 ( .A(n154), .B(n91), .Z(\ab[11][10] ) );
  NR2 U1308 ( .A(n164), .B(n91), .Z(\ab[11][0] ) );
  NR2 U1309 ( .A(n155), .B(n89), .Z(\ab[10][9] ) );
  NR2 U1310 ( .A(n156), .B(n89), .Z(\ab[10][8] ) );
  NR2 U1311 ( .A(n157), .B(n89), .Z(\ab[10][7] ) );
  NR2 U1312 ( .A(n158), .B(n89), .Z(\ab[10][6] ) );
  NR2 U1313 ( .A(n159), .B(n89), .Z(\ab[10][5] ) );
  NR2 U1314 ( .A(n160), .B(n89), .Z(\ab[10][4] ) );
  NR2 U1315 ( .A(n108), .B(n89), .Z(\ab[10][47] ) );
  NR2 U1316 ( .A(n107), .B(n89), .Z(\ab[10][46] ) );
  NR2 U1317 ( .A(n106), .B(n89), .Z(\ab[10][45] ) );
  NR2 U1318 ( .A(n105), .B(n89), .Z(\ab[10][44] ) );
  NR2 U1319 ( .A(n104), .B(n89), .Z(\ab[10][43] ) );
  NR2 U1320 ( .A(n103), .B(n89), .Z(\ab[10][42] ) );
  NR2 U1321 ( .A(n102), .B(n88), .Z(\ab[10][41] ) );
  NR2 U1322 ( .A(n101), .B(n88), .Z(\ab[10][40] ) );
  NR2 U1323 ( .A(n161), .B(n88), .Z(\ab[10][3] ) );
  NR2 U1324 ( .A(n125), .B(n88), .Z(\ab[10][39] ) );
  NR2 U1325 ( .A(n126), .B(n88), .Z(\ab[10][38] ) );
  NR2 U1326 ( .A(n127), .B(n88), .Z(\ab[10][37] ) );
  NR2 U1327 ( .A(n128), .B(n88), .Z(\ab[10][36] ) );
  NR2 U1328 ( .A(n129), .B(n88), .Z(\ab[10][35] ) );
  NR2 U1329 ( .A(n130), .B(n88), .Z(\ab[10][34] ) );
  NR2 U1330 ( .A(n131), .B(n88), .Z(\ab[10][33] ) );
  NR2 U1331 ( .A(n132), .B(n88), .Z(\ab[10][32] ) );
  NR2 U1332 ( .A(n133), .B(n88), .Z(\ab[10][31] ) );
  NR2 U1333 ( .A(n134), .B(n87), .Z(\ab[10][30] ) );
  NR2 U1334 ( .A(n162), .B(n87), .Z(\ab[10][2] ) );
  NR2 U1335 ( .A(n135), .B(n87), .Z(\ab[10][29] ) );
  NR2 U1336 ( .A(n136), .B(n87), .Z(\ab[10][28] ) );
  NR2 U1337 ( .A(n137), .B(n87), .Z(\ab[10][27] ) );
  NR2 U1338 ( .A(n138), .B(n87), .Z(\ab[10][26] ) );
  NR2 U1339 ( .A(n139), .B(n87), .Z(\ab[10][25] ) );
  NR2 U1340 ( .A(n140), .B(n87), .Z(\ab[10][24] ) );
  NR2 U1341 ( .A(n141), .B(n87), .Z(\ab[10][23] ) );
  NR2 U1342 ( .A(n142), .B(n87), .Z(\ab[10][22] ) );
  NR2 U1343 ( .A(n143), .B(n87), .Z(\ab[10][21] ) );
  NR2 U1344 ( .A(n144), .B(n87), .Z(\ab[10][20] ) );
  NR2 U1345 ( .A(n163), .B(n86), .Z(\ab[10][1] ) );
  NR2 U1346 ( .A(n145), .B(n86), .Z(\ab[10][19] ) );
  NR2 U1347 ( .A(n146), .B(n86), .Z(\ab[10][18] ) );
  NR2 U1348 ( .A(n147), .B(n86), .Z(\ab[10][17] ) );
  NR2 U1349 ( .A(n148), .B(n86), .Z(\ab[10][16] ) );
  NR2 U1350 ( .A(n149), .B(n86), .Z(\ab[10][15] ) );
  NR2 U1351 ( .A(n150), .B(n86), .Z(\ab[10][14] ) );
  NR2 U1352 ( .A(n151), .B(n86), .Z(\ab[10][13] ) );
  NR2 U1353 ( .A(n152), .B(n86), .Z(\ab[10][12] ) );
  NR2 U1354 ( .A(n153), .B(n86), .Z(\ab[10][11] ) );
  NR2 U1355 ( .A(n154), .B(n86), .Z(\ab[10][10] ) );
  NR2 U1356 ( .A(n164), .B(n86), .Z(\ab[10][0] ) );
  NR2 U1357 ( .A(n155), .B(n39), .Z(\ab[0][9] ) );
  NR2 U1358 ( .A(n156), .B(n39), .Z(\ab[0][8] ) );
  NR2 U1359 ( .A(n157), .B(n39), .Z(\ab[0][7] ) );
  NR2 U1360 ( .A(n158), .B(n39), .Z(\ab[0][6] ) );
  NR2 U1361 ( .A(n159), .B(n39), .Z(\ab[0][5] ) );
  NR2 U1362 ( .A(n160), .B(n39), .Z(\ab[0][4] ) );
  NR2 U1363 ( .A(n108), .B(n39), .Z(\ab[0][47] ) );
  NR2 U1364 ( .A(n107), .B(n39), .Z(\ab[0][46] ) );
  NR2 U1365 ( .A(n106), .B(n39), .Z(\ab[0][45] ) );
  NR2 U1366 ( .A(n105), .B(n39), .Z(\ab[0][44] ) );
  NR2 U1367 ( .A(n104), .B(n38), .Z(\ab[0][43] ) );
  NR2 U1368 ( .A(n103), .B(n38), .Z(\ab[0][42] ) );
  NR2 U1369 ( .A(n102), .B(n38), .Z(\ab[0][41] ) );
  NR2 U1370 ( .A(n101), .B(n38), .Z(\ab[0][40] ) );
  NR2 U1371 ( .A(n161), .B(n38), .Z(\ab[0][3] ) );
  NR2 U1372 ( .A(n125), .B(n38), .Z(\ab[0][39] ) );
  NR2 U1373 ( .A(n126), .B(n38), .Z(\ab[0][38] ) );
  NR2 U1374 ( .A(n127), .B(n38), .Z(\ab[0][37] ) );
  NR2 U1375 ( .A(n128), .B(n38), .Z(\ab[0][36] ) );
  NR2 U1376 ( .A(n129), .B(n38), .Z(\ab[0][35] ) );
  NR2 U1377 ( .A(n130), .B(n38), .Z(\ab[0][34] ) );
  NR2 U1378 ( .A(n131), .B(n38), .Z(\ab[0][33] ) );
  NR2 U1379 ( .A(n132), .B(n37), .Z(\ab[0][32] ) );
  NR2 U1380 ( .A(n133), .B(n37), .Z(\ab[0][31] ) );
  NR2 U1381 ( .A(n134), .B(n37), .Z(\ab[0][30] ) );
  NR2 U1382 ( .A(n162), .B(n37), .Z(\ab[0][2] ) );
  NR2 U1383 ( .A(n135), .B(n37), .Z(\ab[0][29] ) );
  NR2 U1384 ( .A(n136), .B(n37), .Z(\ab[0][28] ) );
  NR2 U1385 ( .A(n137), .B(n37), .Z(\ab[0][27] ) );
  NR2 U1386 ( .A(n138), .B(n37), .Z(\ab[0][26] ) );
  NR2 U1387 ( .A(n139), .B(n37), .Z(\ab[0][25] ) );
  NR2 U1388 ( .A(n140), .B(n37), .Z(\ab[0][24] ) );
  NR2 U1389 ( .A(n141), .B(n37), .Z(\ab[0][23] ) );
  NR2 U1390 ( .A(n142), .B(n37), .Z(\ab[0][22] ) );
  NR2 U1391 ( .A(n143), .B(n36), .Z(\ab[0][21] ) );
  NR2 U1392 ( .A(n144), .B(n36), .Z(\ab[0][20] ) );
  NR2 U1393 ( .A(n145), .B(n36), .Z(\ab[0][19] ) );
  NR2 U1394 ( .A(n146), .B(n36), .Z(\ab[0][18] ) );
  NR2 U1395 ( .A(n147), .B(n36), .Z(\ab[0][17] ) );
  NR2 U1396 ( .A(n148), .B(n36), .Z(\ab[0][16] ) );
  NR2 U1397 ( .A(n149), .B(n36), .Z(\ab[0][15] ) );
  NR2 U1398 ( .A(n150), .B(n36), .Z(\ab[0][14] ) );
  NR2 U1399 ( .A(n151), .B(n36), .Z(\ab[0][13] ) );
  NR2 U1400 ( .A(n152), .B(n36), .Z(\ab[0][12] ) );
  NR2 U1401 ( .A(n153), .B(n36), .Z(\ab[0][11] ) );
  NR2 U1402 ( .A(n154), .B(n36), .Z(\ab[0][10] ) );
  AN3 U1403 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U1404 ( .A(n41), .B(n163), .Z(\ab[1][1] ) );
endmodule


module LOG_POLY_DW01_add_6 ( A, B, CI, SUM, CO );
  input [123:0] A;
  input [123:0] B;
  output [123:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  AN4P U2 ( .A(n502), .B(n467), .C(n465), .D(n472), .Z(n1) );
  OR2P U3 ( .A(n335), .B(n336), .Z(n2) );
  AN2P U4 ( .A(B[47]), .B(A[47]), .Z(n3) );
  AN2P U5 ( .A(B[67]), .B(A[67]), .Z(n4) );
  AO7 U6 ( .A(n38), .B(n169), .C(n226), .Z(n254) );
  NR2 U7 ( .A(n2), .B(n295), .Z(n279) );
  IVP U8 ( .A(n296), .Z(n295) );
  ND2 U9 ( .A(n265), .B(n266), .Z(n43) );
  ND2 U10 ( .A(n267), .B(n87), .Z(n266) );
  ND4 U11 ( .A(n272), .B(n273), .C(n274), .D(n383), .Z(n271) );
  NR2 U12 ( .A(n368), .B(n369), .Z(n272) );
  NR3 U13 ( .A(n361), .B(n362), .C(n363), .Z(n273) );
  ND2 U14 ( .A(n275), .B(n276), .Z(n274) );
  NR2 U15 ( .A(n297), .B(n3), .Z(n277) );
  ND4 U16 ( .A(n279), .B(n280), .C(n281), .D(n282), .Z(n278) );
  AO7 U17 ( .A(n62), .B(n63), .C(n64), .Z(n60) );
  AO7 U18 ( .A(n189), .B(n158), .C(n190), .Z(n186) );
  ND2 U19 ( .A(n220), .B(n221), .Z(n217) );
  AO6 U20 ( .A(n224), .B(n167), .C(n225), .Z(n220) );
  ND2 U21 ( .A(n87), .B(n222), .Z(n221) );
  NR2 U22 ( .A(n163), .B(n169), .Z(n224) );
  IVP U23 ( .A(n375), .Z(n383) );
  AO2 U24 ( .A(n166), .B(n167), .C(n168), .D(n87), .Z(n126) );
  IVP U25 ( .A(n169), .Z(n166) );
  NR2 U26 ( .A(n169), .B(n170), .Z(n168) );
  IVP U27 ( .A(n339), .Z(n346) );
  IVP U28 ( .A(n364), .Z(n409) );
  IVP U29 ( .A(n399), .Z(n393) );
  AO7 U30 ( .A(n400), .B(n401), .C(n402), .Z(n399) );
  IVP U31 ( .A(n369), .Z(n402) );
  AO7 U32 ( .A(n409), .B(n410), .C(n411), .Z(n401) );
  IVP U33 ( .A(n367), .Z(n361) );
  IVP U34 ( .A(n370), .Z(n368) );
  NR3 U35 ( .A(n89), .B(n63), .C(n523), .Z(n532) );
  ND2 U36 ( .A(n521), .B(n522), .Z(n170) );
  NR2 U37 ( .A(n523), .B(n63), .Z(n522) );
  NR2 U38 ( .A(n89), .B(n88), .Z(n521) );
  NR2 U39 ( .A(n223), .B(n170), .Z(n222) );
  ND2 U40 ( .A(n365), .B(n366), .Z(n362) );
  NR2 U41 ( .A(n523), .B(n63), .Z(n553) );
  NR2 U42 ( .A(n88), .B(n89), .Z(n86) );
  ND2 U43 ( .A(n162), .B(n159), .Z(n134) );
  NR2 U44 ( .A(n146), .B(n158), .Z(n162) );
  ND4 U45 ( .A(n268), .B(n269), .C(n270), .D(n271), .Z(n87) );
  AO7 U46 ( .A(n443), .B(n444), .C(n445), .Z(n269) );
  ND3 U47 ( .A(A[63]), .B(B[63]), .C(n383), .Z(n268) );
  NR2 U48 ( .A(n371), .B(n372), .Z(n270) );
  NR2 U49 ( .A(n306), .B(n307), .Z(n296) );
  ND2 U50 ( .A(n301), .B(n303), .Z(n306) );
  AO7 U51 ( .A(A[44]), .B(B[44]), .C(n302), .Z(n307) );
  AO7 U52 ( .A(n246), .B(n247), .C(n234), .Z(n243) );
  AO7 U53 ( .A(n251), .B(n252), .C(n253), .Z(n248) );
  ND2 U54 ( .A(n308), .B(n309), .Z(n302) );
  IVP U55 ( .A(B[47]), .Z(n308) );
  IVP U56 ( .A(A[47]), .Z(n309) );
  EN U57 ( .A(n238), .B(n239), .Z(SUM[103]) );
  ND2 U58 ( .A(n233), .B(n228), .Z(n239) );
  ND2 U59 ( .A(n235), .B(n242), .Z(n238) );
  ND2 U60 ( .A(n232), .B(n243), .Z(n242) );
  NR2 U61 ( .A(n353), .B(n354), .Z(n282) );
  ND2 U62 ( .A(n319), .B(n323), .Z(n353) );
  AO7 U63 ( .A(A[40]), .B(B[40]), .C(n320), .Z(n354) );
  ND3 U64 ( .A(n487), .B(n1), .C(n488), .Z(n375) );
  NR2 U65 ( .A(n511), .B(n512), .Z(n487) );
  IVP U66 ( .A(n446), .Z(n488) );
  AO7 U67 ( .A(n52), .B(n53), .C(n54), .Z(n51) );
  AO7 U68 ( .A(n179), .B(n180), .C(n153), .Z(n176) );
  AO2 U69 ( .A(B[62]), .B(A[62]), .C(B[61]), .D(A[61]), .Z(n373) );
  ND2 U70 ( .A(n377), .B(n378), .Z(n376) );
  ND3 U71 ( .A(A[60]), .B(B[60]), .C(n379), .Z(n374) );
  AO7 U72 ( .A(n57), .B(n58), .C(n59), .Z(n55) );
  AO7 U73 ( .A(n184), .B(n185), .C(n147), .Z(n181) );
  ND2 U74 ( .A(n349), .B(n350), .Z(n339) );
  IVP U75 ( .A(B[37]), .Z(n349) );
  IVP U76 ( .A(A[37]), .Z(n350) );
  AO3 U77 ( .A(n324), .B(n325), .C(n293), .D(n282), .Z(n314) );
  AO3 U78 ( .A(n328), .B(n332), .C(n333), .D(n334), .Z(n324) );
  NR2 U79 ( .A(n328), .B(n329), .Z(n325) );
  ND2 U80 ( .A(A[33]), .B(B[33]), .Z(n332) );
  AO7 U81 ( .A(n304), .B(n305), .C(n296), .Z(n275) );
  ND2 U82 ( .A(n340), .B(n341), .Z(n304) );
  AO3 U83 ( .A(n2), .B(n314), .C(n315), .D(n316), .Z(n305) );
  ND3 U84 ( .A(A[39]), .B(B[39]), .C(n282), .Z(n340) );
  AO6 U85 ( .A(n380), .B(n381), .C(n382), .Z(n371) );
  AO2 U86 ( .A(B[59]), .B(A[59]), .C(n433), .D(n396), .Z(n380) );
  AO7 U87 ( .A(n392), .B(n393), .C(n370), .Z(n381) );
  ND2 U88 ( .A(n383), .B(n367), .Z(n382) );
  ND2 U89 ( .A(n343), .B(n344), .Z(n337) );
  IVP U90 ( .A(B[39]), .Z(n343) );
  IVP U91 ( .A(A[39]), .Z(n344) );
  ND2 U92 ( .A(n351), .B(n352), .Z(n338) );
  IVP U93 ( .A(B[38]), .Z(n351) );
  IVP U94 ( .A(A[38]), .Z(n352) );
  ND2 U95 ( .A(n355), .B(n356), .Z(n320) );
  IVP U96 ( .A(B[43]), .Z(n355) );
  IVP U97 ( .A(A[43]), .Z(n356) );
  ND2 U98 ( .A(n359), .B(n360), .Z(n319) );
  IVP U99 ( .A(B[42]), .Z(n359) );
  IVP U100 ( .A(A[42]), .Z(n360) );
  ND2 U101 ( .A(n330), .B(n331), .Z(n294) );
  IVP U102 ( .A(B[33]), .Z(n330) );
  IVP U103 ( .A(A[33]), .Z(n331) );
  ND2 U104 ( .A(n310), .B(n311), .Z(n303) );
  IVP U105 ( .A(B[45]), .Z(n310) );
  IVP U106 ( .A(A[45]), .Z(n311) );
  ND2 U107 ( .A(n312), .B(n313), .Z(n301) );
  IVP U108 ( .A(B[46]), .Z(n312) );
  IVP U109 ( .A(A[46]), .Z(n313) );
  ND2 U110 ( .A(n357), .B(n358), .Z(n323) );
  IVP U111 ( .A(B[41]), .Z(n357) );
  IVP U112 ( .A(A[41]), .Z(n358) );
  ND2 U113 ( .A(n84), .B(n85), .Z(n82) );
  ND2 U114 ( .A(n86), .B(n87), .Z(n85) );
  ND2 U115 ( .A(n92), .B(n93), .Z(n90) );
  ND4 U116 ( .A(n338), .B(n342), .C(n337), .D(n282), .Z(n341) );
  AO3 U117 ( .A(n345), .B(n346), .C(n347), .D(n348), .Z(n342) );
  ND2 U118 ( .A(A[36]), .B(B[36]), .Z(n345) );
  ND2 U119 ( .A(B[37]), .B(A[37]), .Z(n347) );
  ND2 U120 ( .A(n338), .B(n339), .Z(n335) );
  AO7 U121 ( .A(A[36]), .B(B[36]), .C(n337), .Z(n336) );
  ND3 U122 ( .A(B[32]), .B(A[32]), .C(n294), .Z(n329) );
  EN U123 ( .A(n51), .B(n5), .Z(SUM[94]) );
  ND2 U124 ( .A(n50), .B(n48), .Z(n5) );
  EN U125 ( .A(n44), .B(n45), .Z(SUM[95]) );
  ND2 U126 ( .A(n46), .B(n47), .Z(n45) );
  ND2 U127 ( .A(n48), .B(n49), .Z(n44) );
  ND2 U128 ( .A(n50), .B(n51), .Z(n49) );
  EN U129 ( .A(n243), .B(n6), .Z(SUM[102]) );
  ND2 U130 ( .A(n232), .B(n235), .Z(n6) );
  EN U131 ( .A(n176), .B(n7), .Z(SUM[110]) );
  ND2 U132 ( .A(n150), .B(n157), .Z(n7) );
  EN U133 ( .A(n171), .B(n172), .Z(SUM[111]) );
  ND2 U134 ( .A(n151), .B(n156), .Z(n172) );
  ND2 U135 ( .A(n157), .B(n175), .Z(n171) );
  ND2 U136 ( .A(n150), .B(n176), .Z(n175) );
  NR2 U137 ( .A(n384), .B(n385), .Z(n367) );
  ND2 U138 ( .A(n379), .B(n377), .Z(n384) );
  AO7 U139 ( .A(A[60]), .B(B[60]), .C(n378), .Z(n385) );
  NR2 U140 ( .A(n394), .B(n395), .Z(n370) );
  ND2 U141 ( .A(n397), .B(n398), .Z(n394) );
  AO7 U142 ( .A(A[56]), .B(B[56]), .C(n396), .Z(n395) );
  ND2 U143 ( .A(n419), .B(n420), .Z(n364) );
  IVP U144 ( .A(B[51]), .Z(n419) );
  IVP U145 ( .A(A[51]), .Z(n420) );
  AO7 U146 ( .A(n126), .B(n127), .C(n128), .Z(n122) );
  AO6 U147 ( .A(n129), .B(n130), .C(n131), .Z(n128) );
  AO7 U148 ( .A(n33), .B(n34), .C(n35), .Z(n32) );
  AO7 U149 ( .A(n113), .B(n114), .C(n115), .Z(n109) );
  NR3 U150 ( .A(n289), .B(n290), .C(n291), .Z(n280) );
  NR2 U151 ( .A(A[31]), .B(B[31]), .Z(n290) );
  ND2 U152 ( .A(n293), .B(n294), .Z(n289) );
  AO7 U153 ( .A(A[32]), .B(B[32]), .C(n292), .Z(n291) );
  ND2 U154 ( .A(n417), .B(n418), .Z(n365) );
  IVP U155 ( .A(B[50]), .Z(n417) );
  IVP U156 ( .A(A[50]), .Z(n418) );
  ND3 U157 ( .A(n529), .B(n530), .C(n531), .Z(n167) );
  ND2 U158 ( .A(n553), .B(n554), .Z(n530) );
  AO6 U159 ( .A(n93), .B(n532), .C(n533), .Z(n531) );
  AO2 U160 ( .A(n566), .B(n65), .C(n567), .D(n566), .Z(n529) );
  ND4 U161 ( .A(n403), .B(n404), .C(n405), .D(n406), .Z(n369) );
  ND2 U162 ( .A(n407), .B(n408), .Z(n403) );
  IVP U163 ( .A(B[52]), .Z(n407) );
  IVP U164 ( .A(A[52]), .Z(n408) );
  AO7 U165 ( .A(n80), .B(n62), .C(n81), .Z(n78) );
  AO7 U166 ( .A(n38), .B(n39), .C(n40), .Z(n36) );
  AO7 U167 ( .A(n216), .B(n189), .C(n197), .Z(n213) );
  AO7 U168 ( .A(n75), .B(n76), .C(n77), .Z(n73) );
  AO7 U169 ( .A(n199), .B(n212), .C(n198), .Z(n209) );
  AO7 U170 ( .A(n412), .B(n413), .C(n414), .Z(n400) );
  ND2 U171 ( .A(n365), .B(n366), .Z(n413) );
  ND3 U172 ( .A(B[48]), .B(A[48]), .C(n364), .Z(n412) );
  ND4 U173 ( .A(B[49]), .B(A[49]), .C(n364), .D(n365), .Z(n414) );
  AO6 U174 ( .A(n298), .B(n299), .C(n300), .Z(n297) );
  AO2 U175 ( .A(B[46]), .B(A[46]), .C(B[45]), .D(A[45]), .Z(n298) );
  ND2 U176 ( .A(n301), .B(n302), .Z(n300) );
  ND3 U177 ( .A(A[44]), .B(B[44]), .C(n303), .Z(n299) );
  AO3 U178 ( .A(n317), .B(n318), .C(n319), .D(n320), .Z(n316) );
  ND2 U179 ( .A(n321), .B(n322), .Z(n318) );
  AN3 U180 ( .A(A[40]), .B(B[40]), .C(n323), .Z(n317) );
  ND2 U181 ( .A(B[41]), .B(A[41]), .Z(n321) );
  AO3 U182 ( .A(A[64]), .B(B[64]), .C(n445), .D(n456), .Z(n512) );
  ND2 U183 ( .A(n415), .B(n416), .Z(n366) );
  IVP U184 ( .A(B[49]), .Z(n415) );
  IVP U185 ( .A(A[49]), .Z(n416) );
  ND2 U186 ( .A(n326), .B(n327), .Z(n293) );
  IVP U187 ( .A(B[35]), .Z(n326) );
  IVP U188 ( .A(A[35]), .Z(n327) );
  ND2 U189 ( .A(n425), .B(n426), .Z(n404) );
  IVP U190 ( .A(B[55]), .Z(n425) );
  IVP U191 ( .A(A[55]), .Z(n426) );
  ND2 U192 ( .A(n427), .B(n428), .Z(n405) );
  IVP U193 ( .A(B[54]), .Z(n427) );
  IVP U194 ( .A(A[54]), .Z(n428) );
  ND2 U195 ( .A(n513), .B(n514), .Z(n456) );
  IVP U196 ( .A(B[65]), .Z(n513) );
  IVP U197 ( .A(A[65]), .Z(n514) );
  ND2 U198 ( .A(n434), .B(n435), .Z(n396) );
  IVP U199 ( .A(B[59]), .Z(n434) );
  IVP U200 ( .A(A[59]), .Z(n435) );
  ND2 U201 ( .A(n390), .B(n391), .Z(n379) );
  IVP U202 ( .A(B[61]), .Z(n390) );
  IVP U203 ( .A(A[61]), .Z(n391) );
  ND2 U204 ( .A(n386), .B(n387), .Z(n378) );
  IVP U205 ( .A(B[62]), .Z(n386) );
  IVP U206 ( .A(A[62]), .Z(n387) );
  ND2 U207 ( .A(n388), .B(n389), .Z(n377) );
  IVP U208 ( .A(B[63]), .Z(n388) );
  IVP U209 ( .A(A[63]), .Z(n389) );
  ND2 U210 ( .A(n69), .B(n568), .Z(n65) );
  AO7 U211 ( .A(n569), .B(n570), .C(n68), .Z(n568) );
  ND2 U212 ( .A(n431), .B(n432), .Z(n406) );
  IVP U213 ( .A(B[53]), .Z(n431) );
  IVP U214 ( .A(A[53]), .Z(n432) );
  ND2 U215 ( .A(n120), .B(n121), .Z(n116) );
  ND2 U216 ( .A(n122), .B(n123), .Z(n121) );
  ND4 U217 ( .A(n457), .B(n458), .C(n459), .D(n460), .Z(n443) );
  NR2 U218 ( .A(n473), .B(n474), .Z(n458) );
  AO3 U219 ( .A(n479), .B(n24), .C(n480), .D(n481), .Z(n457) );
  AN3 U220 ( .A(A[52]), .B(B[52]), .C(n406), .Z(n423) );
  ND3 U221 ( .A(n284), .B(n285), .C(n283), .Z(n281) );
  ND2 U222 ( .A(B[31]), .B(A[31]), .Z(n283) );
  ND2 U223 ( .A(B[30]), .B(A[30]), .Z(n284) );
  ND3 U224 ( .A(A[29]), .B(B[29]), .C(n286), .Z(n285) );
  ND3 U225 ( .A(A[64]), .B(B[64]), .C(n456), .Z(n451) );
  ND2 U226 ( .A(n287), .B(n288), .Z(n286) );
  IVP U227 ( .A(B[30]), .Z(n287) );
  IVP U228 ( .A(A[30]), .Z(n288) );
  ND2 U229 ( .A(n454), .B(n455), .Z(n511) );
  ND2 U230 ( .A(n421), .B(n422), .Z(n392) );
  ND2 U231 ( .A(B[55]), .B(A[55]), .Z(n421) );
  AO3 U232 ( .A(n423), .B(n424), .C(n405), .D(n404), .Z(n422) );
  ND2 U233 ( .A(n429), .B(n430), .Z(n424) );
  EO U234 ( .A(n66), .B(n67), .Z(SUM[91]) );
  AO7 U235 ( .A(n70), .B(n71), .C(n72), .Z(n66) );
  EN U236 ( .A(n25), .B(n26), .Z(SUM[99]) );
  ND2 U237 ( .A(n27), .B(n28), .Z(n26) );
  ND2 U238 ( .A(n29), .B(n30), .Z(n25) );
  ND2 U239 ( .A(n31), .B(n32), .Z(n30) );
  EO U240 ( .A(n204), .B(n205), .Z(SUM[107]) );
  AO7 U241 ( .A(n200), .B(n208), .C(n196), .Z(n204) );
  EN U242 ( .A(n109), .B(n8), .Z(SUM[115]) );
  ND2 U243 ( .A(n110), .B(n107), .Z(n8) );
  ND2 U244 ( .A(n109), .B(n110), .Z(n108) );
  ND4 U245 ( .A(n68), .B(n74), .C(n79), .D(n83), .Z(n63) );
  ND4 U246 ( .A(n61), .B(n56), .C(n50), .D(n46), .Z(n523) );
  ND3 U247 ( .A(n96), .B(n103), .C(n102), .Z(n89) );
  AO7 U248 ( .A(n555), .B(n101), .C(n96), .Z(n91) );
  AO7 U249 ( .A(n436), .B(n437), .C(n438), .Z(n433) );
  ND2 U250 ( .A(B[58]), .B(A[58]), .Z(n438) );
  AO2 U251 ( .A(B[57]), .B(A[57]), .C(B[56]), .D(A[56]), .Z(n436) );
  ND2 U252 ( .A(n397), .B(n398), .Z(n437) );
  AO7 U253 ( .A(A[48]), .B(B[48]), .C(n364), .Z(n363) );
  NR2 U254 ( .A(A[34]), .B(B[34]), .Z(n328) );
  ND2 U255 ( .A(n439), .B(n440), .Z(n398) );
  IVP U256 ( .A(B[57]), .Z(n439) );
  IVP U257 ( .A(A[57]), .Z(n440) );
  ND2 U258 ( .A(n441), .B(n442), .Z(n397) );
  IVP U259 ( .A(B[58]), .Z(n441) );
  IVP U260 ( .A(A[58]), .Z(n442) );
  IVP U261 ( .A(n104), .Z(n88) );
  ND2 U262 ( .A(B[35]), .B(A[35]), .Z(n334) );
  ND2 U263 ( .A(B[34]), .B(A[34]), .Z(n333) );
  ND2 U264 ( .A(B[42]), .B(A[42]), .Z(n322) );
  ND2 U265 ( .A(B[38]), .B(A[38]), .Z(n348) );
  ND2 U266 ( .A(B[51]), .B(A[51]), .Z(n411) );
  ND2 U267 ( .A(A[50]), .B(B[50]), .Z(n410) );
  ND2 U268 ( .A(B[53]), .B(A[53]), .Z(n430) );
  ND2 U269 ( .A(B[54]), .B(A[54]), .Z(n429) );
  EN U270 ( .A(n73), .B(n9), .Z(SUM[90]) );
  ND2 U271 ( .A(n74), .B(n72), .Z(n9) );
  EN U272 ( .A(n55), .B(n10), .Z(SUM[93]) );
  ND2 U273 ( .A(n56), .B(n54), .Z(n10) );
  EN U274 ( .A(n32), .B(n11), .Z(SUM[98]) );
  ND2 U275 ( .A(n31), .B(n29), .Z(n11) );
  EN U276 ( .A(n248), .B(n12), .Z(SUM[101]) );
  ND2 U277 ( .A(n236), .B(n234), .Z(n12) );
  EN U278 ( .A(n209), .B(n13), .Z(SUM[106]) );
  ND2 U279 ( .A(n201), .B(n196), .Z(n13) );
  EN U280 ( .A(n181), .B(n14), .Z(SUM[109]) );
  ND2 U281 ( .A(n165), .B(n153), .Z(n14) );
  EN U282 ( .A(n116), .B(n15), .Z(SUM[114]) );
  ND2 U283 ( .A(n117), .B(n115), .Z(n15) );
  IVP U284 ( .A(n472), .Z(n469) );
  ND4 U285 ( .A(n27), .B(n41), .C(n37), .D(n31), .Z(n169) );
  ND4 U286 ( .A(n233), .B(n232), .C(n236), .D(n237), .Z(n163) );
  AO7 U287 ( .A(n140), .B(n141), .C(n142), .Z(n129) );
  AO6 U288 ( .A(n159), .B(n160), .C(n161), .Z(n140) );
  AO6 U289 ( .A(n143), .B(n144), .C(n145), .Z(n142) );
  AO3 U290 ( .A(n54), .B(n534), .C(n535), .D(n47), .Z(n533) );
  ND2 U291 ( .A(n50), .B(n46), .Z(n534) );
  ND2 U292 ( .A(n536), .B(n46), .Z(n535) );
  AO7 U293 ( .A(n226), .B(n163), .C(n227), .Z(n225) );
  AO6 U294 ( .A(n104), .B(n87), .C(n93), .Z(n98) );
  ND2 U295 ( .A(n191), .B(n192), .Z(n144) );
  AO7 U296 ( .A(n193), .B(n194), .C(n195), .Z(n192) );
  ND2 U297 ( .A(B[43]), .B(A[43]), .Z(n315) );
  EN U298 ( .A(n94), .B(n95), .Z(SUM[87]) );
  ND2 U299 ( .A(n96), .B(n97), .Z(n95) );
  AO7 U300 ( .A(n98), .B(n99), .C(n100), .Z(n94) );
  ND2 U301 ( .A(n102), .B(n103), .Z(n99) );
  EN U302 ( .A(n78), .B(n16), .Z(SUM[89]) );
  ND2 U303 ( .A(n79), .B(n77), .Z(n16) );
  EN U304 ( .A(n60), .B(n17), .Z(SUM[92]) );
  ND2 U305 ( .A(n61), .B(n59), .Z(n17) );
  EN U306 ( .A(n36), .B(n18), .Z(SUM[97]) );
  ND2 U307 ( .A(n37), .B(n35), .Z(n18) );
  EN U308 ( .A(n255), .B(n254), .Z(SUM[100]) );
  ND2 U309 ( .A(n253), .B(n237), .Z(n255) );
  EN U310 ( .A(n213), .B(n19), .Z(SUM[105]) );
  ND2 U311 ( .A(n202), .B(n198), .Z(n19) );
  EN U312 ( .A(n186), .B(n20), .Z(SUM[108]) );
  ND2 U313 ( .A(n164), .B(n147), .Z(n20) );
  EO U314 ( .A(n135), .B(n136), .Z(SUM[112]) );
  AO7 U315 ( .A(n126), .B(n134), .C(n139), .Z(n135) );
  EN U316 ( .A(n122), .B(n21), .Z(SUM[113]) );
  ND2 U317 ( .A(n123), .B(n120), .Z(n21) );
  ND4 U318 ( .A(n164), .B(n165), .C(n150), .D(n151), .Z(n146) );
  AO3 U319 ( .A(n146), .B(n147), .C(n148), .D(n149), .Z(n145) );
  ND3 U320 ( .A(n150), .B(n151), .C(n152), .Z(n149) );
  AO6 U321 ( .A(n154), .B(n151), .C(n155), .Z(n148) );
  EN U322 ( .A(n82), .B(n22), .Z(SUM[88]) );
  ND2 U323 ( .A(n81), .B(n83), .Z(n22) );
  EN U324 ( .A(n42), .B(n43), .Z(SUM[96]) );
  ND2 U325 ( .A(n40), .B(n41), .Z(n42) );
  EN U326 ( .A(n217), .B(n23), .Z(SUM[104]) );
  ND2 U327 ( .A(n197), .B(n203), .Z(n23) );
  ND4 U328 ( .A(n195), .B(n201), .C(n202), .D(n203), .Z(n158) );
  IVP U329 ( .A(n101), .Z(n100) );
  ND2 U330 ( .A(n489), .B(n481), .Z(n446) );
  NR2 U331 ( .A(n494), .B(n495), .Z(n489) );
  ND2 U332 ( .A(n485), .B(n486), .Z(n495) );
  AO7 U333 ( .A(A[72]), .B(B[72]), .C(n480), .Z(n494) );
  AO3 U334 ( .A(A[76]), .B(B[76]), .C(n463), .D(n464), .Z(n477) );
  ND2 U335 ( .A(n492), .B(n493), .Z(n463) );
  IVP U336 ( .A(B[78]), .Z(n492) );
  IVP U337 ( .A(A[78]), .Z(n493) );
  ND2 U338 ( .A(n498), .B(n499), .Z(n485) );
  IVP U339 ( .A(B[73]), .Z(n498) );
  IVP U340 ( .A(A[73]), .Z(n499) );
  ND2 U341 ( .A(n496), .B(n497), .Z(n486) );
  IVP U342 ( .A(B[74]), .Z(n496) );
  IVP U343 ( .A(A[74]), .Z(n497) );
  ND2 U344 ( .A(n490), .B(n491), .Z(n464) );
  IVP U345 ( .A(B[77]), .Z(n490) );
  IVP U346 ( .A(A[77]), .Z(n491) );
  ND2 U347 ( .A(n500), .B(n501), .Z(n480) );
  IVP U348 ( .A(B[75]), .Z(n500) );
  IVP U349 ( .A(A[75]), .Z(n501) );
  ND2 U350 ( .A(n509), .B(n510), .Z(n502) );
  IVP U351 ( .A(B[68]), .Z(n509) );
  IVP U352 ( .A(A[68]), .Z(n510) );
  NR3 U353 ( .A(n482), .B(n483), .C(n484), .Z(n479) );
  AO2 U354 ( .A(B[73]), .B(A[73]), .C(B[72]), .D(A[72]), .Z(n483) );
  IVP U355 ( .A(n486), .Z(n482) );
  IVP U356 ( .A(n485), .Z(n484) );
  AO2 U357 ( .A(B[66]), .B(A[66]), .C(B[65]), .D(A[65]), .Z(n450) );
  IVP U358 ( .A(n455), .Z(n452) );
  IVP U359 ( .A(n454), .Z(n453) );
  ND2 U360 ( .A(n519), .B(n520), .Z(n454) );
  IVP U361 ( .A(B[66]), .Z(n519) );
  IVP U362 ( .A(A[66]), .Z(n520) );
  ND2 U363 ( .A(n517), .B(n518), .Z(n455) );
  IVP U364 ( .A(B[67]), .Z(n517) );
  IVP U365 ( .A(A[67]), .Z(n518) );
  ND2 U366 ( .A(n503), .B(n504), .Z(n472) );
  IVP U367 ( .A(B[69]), .Z(n503) );
  IVP U368 ( .A(A[69]), .Z(n504) );
  ND2 U369 ( .A(n573), .B(n574), .Z(n74) );
  IVP U370 ( .A(B[90]), .Z(n573) );
  IVP U371 ( .A(A[90]), .Z(n574) );
  ND2 U372 ( .A(n575), .B(n576), .Z(n79) );
  IVP U373 ( .A(B[89]), .Z(n575) );
  IVP U374 ( .A(A[89]), .Z(n576) );
  AO7 U375 ( .A(n446), .B(n447), .C(n448), .Z(n444) );
  AO7 U376 ( .A(n449), .B(n4), .C(n1), .Z(n447) );
  ND3 U377 ( .A(A[71]), .B(B[71]), .C(n488), .Z(n448) );
  ND2 U378 ( .A(n505), .B(n506), .Z(n465) );
  IVP U379 ( .A(B[70]), .Z(n505) );
  IVP U380 ( .A(A[70]), .Z(n506) );
  ND2 U381 ( .A(n507), .B(n508), .Z(n467) );
  IVP U382 ( .A(B[71]), .Z(n507) );
  IVP U383 ( .A(A[71]), .Z(n508) );
  ND2 U384 ( .A(n515), .B(n516), .Z(n445) );
  IVP U385 ( .A(B[79]), .Z(n515) );
  IVP U386 ( .A(A[79]), .Z(n516) );
  ND4 U387 ( .A(n465), .B(n466), .C(n467), .D(n488), .Z(n459) );
  AO3 U388 ( .A(n468), .B(n469), .C(n470), .D(n471), .Z(n466) );
  ND2 U389 ( .A(A[68]), .B(B[68]), .Z(n468) );
  AO7 U390 ( .A(n537), .B(n558), .C(n559), .Z(n101) );
  ND2 U391 ( .A(A[84]), .B(B[84]), .Z(n558) );
  AO2 U392 ( .A(B[86]), .B(A[86]), .C(n560), .D(n561), .Z(n559) );
  NR2 U393 ( .A(n524), .B(n525), .Z(n104) );
  ND2 U394 ( .A(n527), .B(n528), .Z(n524) );
  AO7 U395 ( .A(A[80]), .B(B[80]), .C(n526), .Z(n525) );
  ND2 U396 ( .A(n577), .B(n578), .Z(n46) );
  IVP U397 ( .A(B[95]), .Z(n577) );
  IVP U398 ( .A(A[95]), .Z(n578) );
  AO7 U399 ( .A(A[85]), .B(B[85]), .C(n561), .Z(n537) );
  NR3 U400 ( .A(n546), .B(n547), .C(n548), .Z(n542) );
  AO2 U401 ( .A(B[80]), .B(A[80]), .C(B[81]), .D(A[81]), .Z(n546) );
  ND2 U402 ( .A(n556), .B(n557), .Z(n96) );
  IVP U403 ( .A(B[87]), .Z(n556) );
  IVP U404 ( .A(A[87]), .Z(n557) );
  ND2 U405 ( .A(n540), .B(n541), .Z(n93) );
  ND2 U406 ( .A(B[83]), .B(A[83]), .Z(n540) );
  AO7 U407 ( .A(n542), .B(n543), .C(n526), .Z(n541) );
  ND2 U408 ( .A(B[89]), .B(A[89]), .Z(n77) );
  ND2 U409 ( .A(B[88]), .B(A[88]), .Z(n81) );
  ND2 U410 ( .A(n571), .B(n572), .Z(n68) );
  IVP U411 ( .A(B[91]), .Z(n571) );
  IVP U412 ( .A(A[91]), .Z(n572) );
  ND2 U413 ( .A(n581), .B(n582), .Z(n56) );
  IVP U414 ( .A(B[93]), .Z(n581) );
  IVP U415 ( .A(A[93]), .Z(n582) );
  ND2 U416 ( .A(n583), .B(n584), .Z(n61) );
  IVP U417 ( .A(B[92]), .Z(n583) );
  IVP U418 ( .A(A[92]), .Z(n584) );
  ND2 U419 ( .A(n564), .B(n565), .Z(n83) );
  IVP U420 ( .A(B[88]), .Z(n564) );
  IVP U421 ( .A(A[88]), .Z(n565) );
  NR2 U422 ( .A(n477), .B(n478), .Z(n473) );
  ND2 U423 ( .A(A[75]), .B(B[75]), .Z(n478) );
  ND2 U424 ( .A(n562), .B(n563), .Z(n561) );
  IVP U425 ( .A(B[86]), .Z(n562) );
  IVP U426 ( .A(A[86]), .Z(n563) );
  ND2 U427 ( .A(n544), .B(n545), .Z(n526) );
  IVP U428 ( .A(B[83]), .Z(n544) );
  IVP U429 ( .A(A[83]), .Z(n545) );
  ND2 U430 ( .A(n551), .B(n552), .Z(n528) );
  IVP U431 ( .A(B[81]), .Z(n551) );
  IVP U432 ( .A(A[81]), .Z(n552) );
  ND2 U433 ( .A(n549), .B(n550), .Z(n527) );
  IVP U434 ( .A(B[82]), .Z(n549) );
  IVP U435 ( .A(A[82]), .Z(n550) );
  ND4 U436 ( .A(B[76]), .B(A[76]), .C(n463), .D(n464), .Z(n462) );
  ND2 U437 ( .A(n579), .B(n580), .Z(n50) );
  IVP U438 ( .A(B[94]), .Z(n579) );
  IVP U439 ( .A(A[94]), .Z(n580) );
  ND3 U440 ( .A(A[77]), .B(B[77]), .C(n463), .Z(n461) );
  ND2 U441 ( .A(n259), .B(n260), .Z(n31) );
  IVP U442 ( .A(B[98]), .Z(n259) );
  IVP U443 ( .A(A[98]), .Z(n260) );
  ND2 U444 ( .A(n244), .B(n245), .Z(n232) );
  IVP U445 ( .A(B[102]), .Z(n244) );
  IVP U446 ( .A(A[102]), .Z(n245) );
  ND2 U447 ( .A(n263), .B(n264), .Z(n27) );
  IVP U448 ( .A(B[99]), .Z(n263) );
  IVP U449 ( .A(A[99]), .Z(n264) );
  ND2 U450 ( .A(n240), .B(n241), .Z(n233) );
  IVP U451 ( .A(B[103]), .Z(n240) );
  IVP U452 ( .A(A[103]), .Z(n241) );
  ND2 U453 ( .A(n261), .B(n262), .Z(n37) );
  IVP U454 ( .A(B[97]), .Z(n261) );
  IVP U455 ( .A(A[97]), .Z(n262) );
  ND2 U456 ( .A(n249), .B(n250), .Z(n236) );
  IVP U457 ( .A(B[101]), .Z(n249) );
  IVP U458 ( .A(A[101]), .Z(n250) );
  ND2 U459 ( .A(n214), .B(n215), .Z(n202) );
  IVP U460 ( .A(B[105]), .Z(n214) );
  IVP U461 ( .A(A[105]), .Z(n215) );
  ND2 U462 ( .A(n210), .B(n211), .Z(n201) );
  IVP U463 ( .A(B[106]), .Z(n210) );
  IVP U464 ( .A(A[106]), .Z(n211) );
  ND2 U465 ( .A(n538), .B(n539), .Z(n103) );
  IVP U466 ( .A(B[84]), .Z(n538) );
  IVP U467 ( .A(A[84]), .Z(n539) );
  ND2 U468 ( .A(n28), .B(n256), .Z(n160) );
  AO3 U469 ( .A(n257), .B(n258), .C(n31), .D(n27), .Z(n256) );
  ND2 U470 ( .A(n35), .B(n29), .Z(n258) );
  AN3 U471 ( .A(A[96]), .B(B[96]), .C(n37), .Z(n257) );
  ND2 U472 ( .A(n228), .B(n229), .Z(n161) );
  AO3 U473 ( .A(n230), .B(n231), .C(n232), .D(n233), .Z(n229) );
  ND2 U474 ( .A(n234), .B(n235), .Z(n231) );
  AN3 U475 ( .A(A[100]), .B(B[100]), .C(n236), .Z(n230) );
  ND2 U476 ( .A(B[69]), .B(A[69]), .Z(n471) );
  ND2 U477 ( .A(B[70]), .B(A[70]), .Z(n470) );
  ND2 U478 ( .A(n475), .B(n476), .Z(n474) );
  ND2 U479 ( .A(B[78]), .B(A[78]), .Z(n475) );
  ND2 U480 ( .A(B[79]), .B(A[79]), .Z(n476) );
  AN2P U481 ( .A(B[74]), .B(A[74]), .Z(n24) );
  ND2 U482 ( .A(n173), .B(n174), .Z(n151) );
  IVP U483 ( .A(B[111]), .Z(n173) );
  IVP U484 ( .A(A[111]), .Z(n174) );
  ND2 U485 ( .A(B[93]), .B(A[93]), .Z(n54) );
  ND2 U486 ( .A(B[98]), .B(A[98]), .Z(n29) );
  ND2 U487 ( .A(B[97]), .B(A[97]), .Z(n35) );
  ND2 U488 ( .A(B[104]), .B(A[104]), .Z(n197) );
  ND2 U489 ( .A(B[101]), .B(A[101]), .Z(n234) );
  ND2 U490 ( .A(B[105]), .B(A[105]), .Z(n198) );
  ND2 U491 ( .A(B[102]), .B(A[102]), .Z(n235) );
  ND2 U492 ( .A(B[90]), .B(A[90]), .Z(n72) );
  ND2 U493 ( .A(B[94]), .B(A[94]), .Z(n48) );
  ND2 U494 ( .A(B[110]), .B(A[110]), .Z(n157) );
  ND2 U495 ( .A(B[95]), .B(A[95]), .Z(n47) );
  ND2 U496 ( .A(B[87]), .B(A[87]), .Z(n97) );
  ND2 U497 ( .A(B[111]), .B(A[111]), .Z(n156) );
  ND2 U498 ( .A(B[91]), .B(A[91]), .Z(n69) );
  ND2 U499 ( .A(n177), .B(n178), .Z(n150) );
  IVP U500 ( .A(B[110]), .Z(n177) );
  IVP U501 ( .A(A[110]), .Z(n178) );
  ND2 U502 ( .A(n206), .B(n207), .Z(n195) );
  IVP U503 ( .A(B[107]), .Z(n206) );
  IVP U504 ( .A(A[107]), .Z(n207) );
  ND2 U505 ( .A(B[92]), .B(A[92]), .Z(n59) );
  ND2 U506 ( .A(n218), .B(n219), .Z(n203) );
  IVP U507 ( .A(B[104]), .Z(n218) );
  IVP U508 ( .A(A[104]), .Z(n219) );
  ND2 U509 ( .A(n182), .B(n183), .Z(n165) );
  IVP U510 ( .A(B[109]), .Z(n182) );
  IVP U511 ( .A(A[109]), .Z(n183) );
  ND2 U512 ( .A(n187), .B(n188), .Z(n164) );
  IVP U513 ( .A(B[108]), .Z(n187) );
  IVP U514 ( .A(A[108]), .Z(n188) );
  ND2 U515 ( .A(B[109]), .B(A[109]), .Z(n153) );
  ND2 U516 ( .A(B[106]), .B(A[106]), .Z(n196) );
  ND2 U517 ( .A(B[99]), .B(A[99]), .Z(n28) );
  ND2 U518 ( .A(B[103]), .B(A[103]), .Z(n228) );
  ND2 U519 ( .A(B[108]), .B(A[108]), .Z(n147) );
  ND2 U520 ( .A(B[107]), .B(A[107]), .Z(n191) );
  ND2 U521 ( .A(n137), .B(n138), .Z(n130) );
  IVP U522 ( .A(B[112]), .Z(n137) );
  IVP U523 ( .A(A[112]), .Z(n138) );
  ND2 U524 ( .A(B[112]), .B(A[112]), .Z(n132) );
  ND2 U525 ( .A(B[96]), .B(A[96]), .Z(n40) );
  ND2 U526 ( .A(B[100]), .B(A[100]), .Z(n253) );
  ND2 U527 ( .A(n124), .B(n125), .Z(n123) );
  IVP U528 ( .A(B[113]), .Z(n124) );
  IVP U529 ( .A(A[113]), .Z(n125) );
  ND2 U530 ( .A(B[113]), .B(A[113]), .Z(n120) );
  ND2 U531 ( .A(n118), .B(n119), .Z(n117) );
  IVP U532 ( .A(B[114]), .Z(n118) );
  IVP U533 ( .A(A[114]), .Z(n119) );
  ND2 U534 ( .A(B[114]), .B(A[114]), .Z(n115) );
  ND2 U535 ( .A(n111), .B(n112), .Z(n110) );
  IVP U536 ( .A(B[115]), .Z(n111) );
  IVP U537 ( .A(A[115]), .Z(n112) );
  ND2 U538 ( .A(B[115]), .B(A[115]), .Z(n107) );
  EO U539 ( .A(n105), .B(n106), .Z(SUM[116]) );
  EO U540 ( .A(B[116]), .B(A[116]), .Z(n106) );
  IVA U541 ( .A(n36), .Z(n34) );
  IVA U542 ( .A(n37), .Z(n33) );
  IVA U543 ( .A(n41), .Z(n39) );
  IVA U544 ( .A(n55), .Z(n53) );
  IVA U545 ( .A(n56), .Z(n52) );
  IVA U546 ( .A(n60), .Z(n58) );
  IVA U547 ( .A(n61), .Z(n57) );
  IVA U548 ( .A(n65), .Z(n64) );
  AN2P U549 ( .A(n68), .B(n69), .Z(n67) );
  IVA U550 ( .A(n73), .Z(n71) );
  IVA U551 ( .A(n78), .Z(n76) );
  IVA U552 ( .A(n82), .Z(n62) );
  IVA U553 ( .A(n83), .Z(n80) );
  AN2P U554 ( .A(n90), .B(n91), .Z(n84) );
  IVA U555 ( .A(n89), .Z(n92) );
  ND2 U556 ( .A(n107), .B(n108), .Z(n105) );
  IVA U557 ( .A(n116), .Z(n114) );
  IVA U558 ( .A(n117), .Z(n113) );
  IVA U559 ( .A(n132), .Z(n131) );
  ND2 U560 ( .A(n133), .B(n130), .Z(n127) );
  IVA U561 ( .A(n134), .Z(n133) );
  AN2P U562 ( .A(n130), .B(n132), .Z(n136) );
  IVA U563 ( .A(n129), .Z(n139) );
  IVA U564 ( .A(n153), .Z(n152) );
  IVA U565 ( .A(n156), .Z(n155) );
  IVA U566 ( .A(n157), .Z(n154) );
  IVA U567 ( .A(n146), .Z(n143) );
  OR2 U568 ( .A(n158), .B(n146), .Z(n141) );
  IVA U569 ( .A(n163), .Z(n159) );
  IVA U570 ( .A(n181), .Z(n180) );
  IVA U571 ( .A(n165), .Z(n179) );
  IVA U572 ( .A(n186), .Z(n185) );
  IVA U573 ( .A(n164), .Z(n184) );
  IVA U574 ( .A(n144), .Z(n190) );
  IVA U575 ( .A(n196), .Z(n194) );
  AO1P U576 ( .A(n197), .B(n198), .C(n199), .D(n200), .Z(n193) );
  AN2P U577 ( .A(n195), .B(n191), .Z(n205) );
  IVA U578 ( .A(n209), .Z(n208) );
  IVA U579 ( .A(n201), .Z(n200) );
  IVA U580 ( .A(n213), .Z(n212) );
  IVA U581 ( .A(n202), .Z(n199) );
  IVA U582 ( .A(n217), .Z(n189) );
  IVA U583 ( .A(n203), .Z(n216) );
  OR2 U584 ( .A(n169), .B(n163), .Z(n223) );
  IVA U585 ( .A(n161), .Z(n227) );
  IVA U586 ( .A(n248), .Z(n247) );
  IVA U587 ( .A(n236), .Z(n246) );
  IVA U588 ( .A(n254), .Z(n252) );
  IVA U589 ( .A(n237), .Z(n251) );
  IVA U590 ( .A(n160), .Z(n226) );
  OR2 U591 ( .A(A[96]), .B(B[96]), .Z(n41) );
  IVA U592 ( .A(n43), .Z(n38) );
  AN2P U593 ( .A(n277), .B(n278), .Z(n276) );
  OR2 U594 ( .A(A[34]), .B(B[34]), .Z(n292) );
  AO1P U595 ( .A(n373), .B(n374), .C(n375), .D(n376), .Z(n372) );
  AO1P U596 ( .A(n450), .B(n451), .C(n452), .D(n453), .Z(n449) );
  AN2P U597 ( .A(n461), .B(n462), .Z(n460) );
  IVA U598 ( .A(n477), .Z(n481) );
  IVA U599 ( .A(n170), .Z(n267) );
  IVA U600 ( .A(n167), .Z(n265) );
  IVA U601 ( .A(n48), .Z(n536) );
  IVA U602 ( .A(n537), .Z(n102) );
  AN2P U603 ( .A(B[82]), .B(A[82]), .Z(n543) );
  IVA U604 ( .A(n527), .Z(n548) );
  IVA U605 ( .A(n528), .Z(n547) );
  IVA U606 ( .A(n91), .Z(n554) );
  AN2P U607 ( .A(A[85]), .B(B[85]), .Z(n560) );
  IVA U608 ( .A(n97), .Z(n555) );
  IVA U609 ( .A(n59), .Z(n567) );
  IVA U610 ( .A(n72), .Z(n570) );
  AO1P U611 ( .A(n81), .B(n77), .C(n75), .D(n70), .Z(n569) );
  IVA U612 ( .A(n74), .Z(n70) );
  IVA U613 ( .A(n79), .Z(n75) );
  IVA U614 ( .A(n523), .Z(n566) );
  OR2 U615 ( .A(A[100]), .B(B[100]), .Z(n237) );
endmodule


module LOG_POLY_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [29:0] A;
  input [95:0] B;
  output [125:0] PRODUCT;
  input TC;
  wire   \ab[29][95] , \ab[29][94] , \ab[29][93] , \ab[29][92] , \ab[29][91] ,
         \ab[29][90] , \ab[29][89] , \ab[29][88] , \ab[29][87] , \ab[29][86] ,
         \ab[29][85] , \ab[29][84] , \ab[29][83] , \ab[29][82] , \ab[29][81] ,
         \ab[29][80] , \ab[29][79] , \ab[29][78] , \ab[29][77] , \ab[29][76] ,
         \ab[29][75] , \ab[29][74] , \ab[29][73] , \ab[29][72] , \ab[29][71] ,
         \ab[29][70] , \ab[29][69] , \ab[29][68] , \ab[29][67] , \ab[29][66] ,
         \ab[29][65] , \ab[29][64] , \ab[29][63] , \ab[29][62] , \ab[29][61] ,
         \ab[29][60] , \ab[29][59] , \ab[29][58] , \ab[29][57] , \ab[29][56] ,
         \ab[29][55] , \ab[29][54] , \ab[29][53] , \ab[29][52] , \ab[29][51] ,
         \ab[29][50] , \ab[29][49] , \ab[29][48] , \ab[29][47] , \ab[29][46] ,
         \ab[29][45] , \ab[29][44] , \ab[29][43] , \ab[29][42] , \ab[29][41] ,
         \ab[29][40] , \ab[29][39] , \ab[29][38] , \ab[29][37] , \ab[29][36] ,
         \ab[29][35] , \ab[29][34] , \ab[29][33] , \ab[29][32] , \ab[29][31] ,
         \ab[29][30] , \ab[29][29] , \ab[29][28] , \ab[29][27] , \ab[29][26] ,
         \ab[29][25] , \ab[29][24] , \ab[29][23] , \ab[29][22] , \ab[29][21] ,
         \ab[29][20] , \ab[29][19] , \ab[29][18] , \ab[29][17] , \ab[29][16] ,
         \ab[29][15] , \ab[29][14] , \ab[29][13] , \ab[29][12] , \ab[29][11] ,
         \ab[29][10] , \ab[29][9] , \ab[29][8] , \ab[29][7] , \ab[29][6] ,
         \ab[29][5] , \ab[29][4] , \ab[29][3] , \ab[29][2] , \ab[29][1] ,
         \ab[29][0] , \ab[28][95] , \ab[28][94] , \ab[28][93] , \ab[28][92] ,
         \ab[28][91] , \ab[28][90] , \ab[28][89] , \ab[28][88] , \ab[28][87] ,
         \ab[28][86] , \ab[28][85] , \ab[28][84] , \ab[28][83] , \ab[28][82] ,
         \ab[28][81] , \ab[28][80] , \ab[28][79] , \ab[28][78] , \ab[28][77] ,
         \ab[28][76] , \ab[28][75] , \ab[28][74] , \ab[28][73] , \ab[28][72] ,
         \ab[28][71] , \ab[28][70] , \ab[28][69] , \ab[28][68] , \ab[28][67] ,
         \ab[28][66] , \ab[28][65] , \ab[28][64] , \ab[28][63] , \ab[28][62] ,
         \ab[28][61] , \ab[28][60] , \ab[28][59] , \ab[28][58] , \ab[28][57] ,
         \ab[28][56] , \ab[28][55] , \ab[28][54] , \ab[28][53] , \ab[28][52] ,
         \ab[28][51] , \ab[28][50] , \ab[28][49] , \ab[28][48] , \ab[28][47] ,
         \ab[28][46] , \ab[28][45] , \ab[28][44] , \ab[28][43] , \ab[28][42] ,
         \ab[28][41] , \ab[28][40] , \ab[28][39] , \ab[28][38] , \ab[28][37] ,
         \ab[28][36] , \ab[28][35] , \ab[28][34] , \ab[28][33] , \ab[28][32] ,
         \ab[28][31] , \ab[28][30] , \ab[28][29] , \ab[28][28] , \ab[28][27] ,
         \ab[28][26] , \ab[28][25] , \ab[28][24] , \ab[28][23] , \ab[28][22] ,
         \ab[28][21] , \ab[28][20] , \ab[28][19] , \ab[28][18] , \ab[28][17] ,
         \ab[28][16] , \ab[28][15] , \ab[28][14] , \ab[28][13] , \ab[28][12] ,
         \ab[28][11] , \ab[28][10] , \ab[28][9] , \ab[28][8] , \ab[28][7] ,
         \ab[28][6] , \ab[28][5] , \ab[28][4] , \ab[28][3] , \ab[28][2] ,
         \ab[28][1] , \ab[28][0] , \ab[27][95] , \ab[27][94] , \ab[27][93] ,
         \ab[27][92] , \ab[27][91] , \ab[27][90] , \ab[27][89] , \ab[27][88] ,
         \ab[27][87] , \ab[27][86] , \ab[27][85] , \ab[27][84] , \ab[27][83] ,
         \ab[27][82] , \ab[27][81] , \ab[27][80] , \ab[27][79] , \ab[27][78] ,
         \ab[27][77] , \ab[27][76] , \ab[27][75] , \ab[27][74] , \ab[27][73] ,
         \ab[27][72] , \ab[27][71] , \ab[27][70] , \ab[27][69] , \ab[27][68] ,
         \ab[27][67] , \ab[27][66] , \ab[27][65] , \ab[27][64] , \ab[27][63] ,
         \ab[27][62] , \ab[27][61] , \ab[27][60] , \ab[27][59] , \ab[27][58] ,
         \ab[27][57] , \ab[27][56] , \ab[27][55] , \ab[27][54] , \ab[27][53] ,
         \ab[27][52] , \ab[27][51] , \ab[27][50] , \ab[27][49] , \ab[27][48] ,
         \ab[27][47] , \ab[27][46] , \ab[27][45] , \ab[27][44] , \ab[27][43] ,
         \ab[27][42] , \ab[27][41] , \ab[27][40] , \ab[27][39] , \ab[27][38] ,
         \ab[27][37] , \ab[27][36] , \ab[27][35] , \ab[27][34] , \ab[27][33] ,
         \ab[27][32] , \ab[27][31] , \ab[27][30] , \ab[27][29] , \ab[27][28] ,
         \ab[27][27] , \ab[27][26] , \ab[27][25] , \ab[27][24] , \ab[27][23] ,
         \ab[27][22] , \ab[27][21] , \ab[27][20] , \ab[27][19] , \ab[27][18] ,
         \ab[27][17] , \ab[27][16] , \ab[27][15] , \ab[27][14] , \ab[27][13] ,
         \ab[27][12] , \ab[27][11] , \ab[27][10] , \ab[27][9] , \ab[27][8] ,
         \ab[27][7] , \ab[27][6] , \ab[27][5] , \ab[27][4] , \ab[27][3] ,
         \ab[27][2] , \ab[27][1] , \ab[27][0] , \ab[26][95] , \ab[26][94] ,
         \ab[26][93] , \ab[26][92] , \ab[26][91] , \ab[26][90] , \ab[26][89] ,
         \ab[26][88] , \ab[26][87] , \ab[26][86] , \ab[26][85] , \ab[26][84] ,
         \ab[26][83] , \ab[26][82] , \ab[26][81] , \ab[26][80] , \ab[26][79] ,
         \ab[26][78] , \ab[26][77] , \ab[26][76] , \ab[26][75] , \ab[26][74] ,
         \ab[26][73] , \ab[26][72] , \ab[26][71] , \ab[26][70] , \ab[26][69] ,
         \ab[26][68] , \ab[26][67] , \ab[26][66] , \ab[26][65] , \ab[26][64] ,
         \ab[26][63] , \ab[26][62] , \ab[26][61] , \ab[26][60] , \ab[26][59] ,
         \ab[26][58] , \ab[26][57] , \ab[26][56] , \ab[26][55] , \ab[26][54] ,
         \ab[26][53] , \ab[26][52] , \ab[26][51] , \ab[26][50] , \ab[26][49] ,
         \ab[26][48] , \ab[26][47] , \ab[26][46] , \ab[26][45] , \ab[26][44] ,
         \ab[26][43] , \ab[26][42] , \ab[26][41] , \ab[26][40] , \ab[26][39] ,
         \ab[26][38] , \ab[26][37] , \ab[26][36] , \ab[26][35] , \ab[26][34] ,
         \ab[26][33] , \ab[26][32] , \ab[26][31] , \ab[26][30] , \ab[26][29] ,
         \ab[26][28] , \ab[26][27] , \ab[26][26] , \ab[26][25] , \ab[26][24] ,
         \ab[26][23] , \ab[26][22] , \ab[26][21] , \ab[26][20] , \ab[26][19] ,
         \ab[26][18] , \ab[26][17] , \ab[26][16] , \ab[26][15] , \ab[26][14] ,
         \ab[26][13] , \ab[26][12] , \ab[26][11] , \ab[26][10] , \ab[26][9] ,
         \ab[26][8] , \ab[26][7] , \ab[26][6] , \ab[26][5] , \ab[26][4] ,
         \ab[26][3] , \ab[26][2] , \ab[26][1] , \ab[26][0] , \ab[25][95] ,
         \ab[25][94] , \ab[25][93] , \ab[25][92] , \ab[25][91] , \ab[25][90] ,
         \ab[25][89] , \ab[25][88] , \ab[25][87] , \ab[25][86] , \ab[25][85] ,
         \ab[25][84] , \ab[25][83] , \ab[25][82] , \ab[25][81] , \ab[25][80] ,
         \ab[25][79] , \ab[25][78] , \ab[25][77] , \ab[25][76] , \ab[25][75] ,
         \ab[25][74] , \ab[25][73] , \ab[25][72] , \ab[25][71] , \ab[25][70] ,
         \ab[25][69] , \ab[25][68] , \ab[25][67] , \ab[25][66] , \ab[25][65] ,
         \ab[25][64] , \ab[25][63] , \ab[25][62] , \ab[25][61] , \ab[25][60] ,
         \ab[25][59] , \ab[25][58] , \ab[25][57] , \ab[25][56] , \ab[25][55] ,
         \ab[25][54] , \ab[25][53] , \ab[25][52] , \ab[25][51] , \ab[25][50] ,
         \ab[25][49] , \ab[25][48] , \ab[25][47] , \ab[25][46] , \ab[25][45] ,
         \ab[25][44] , \ab[25][43] , \ab[25][42] , \ab[25][41] , \ab[25][40] ,
         \ab[25][39] , \ab[25][38] , \ab[25][37] , \ab[25][36] , \ab[25][35] ,
         \ab[25][34] , \ab[25][33] , \ab[25][32] , \ab[25][31] , \ab[25][30] ,
         \ab[25][29] , \ab[25][28] , \ab[25][27] , \ab[25][26] , \ab[25][25] ,
         \ab[25][24] , \ab[25][23] , \ab[25][22] , \ab[25][21] , \ab[25][20] ,
         \ab[25][19] , \ab[25][18] , \ab[25][17] , \ab[25][16] , \ab[25][15] ,
         \ab[25][14] , \ab[25][13] , \ab[25][12] , \ab[25][11] , \ab[25][10] ,
         \ab[25][9] , \ab[25][8] , \ab[25][7] , \ab[25][6] , \ab[25][5] ,
         \ab[25][4] , \ab[25][3] , \ab[25][2] , \ab[25][1] , \ab[25][0] ,
         \ab[24][95] , \ab[24][94] , \ab[24][93] , \ab[24][92] , \ab[24][91] ,
         \ab[24][90] , \ab[24][89] , \ab[24][88] , \ab[24][87] , \ab[24][86] ,
         \ab[24][85] , \ab[24][84] , \ab[24][83] , \ab[24][82] , \ab[24][81] ,
         \ab[24][80] , \ab[24][79] , \ab[24][78] , \ab[24][77] , \ab[24][76] ,
         \ab[24][75] , \ab[24][74] , \ab[24][73] , \ab[24][72] , \ab[24][71] ,
         \ab[24][70] , \ab[24][69] , \ab[24][68] , \ab[24][67] , \ab[24][66] ,
         \ab[24][65] , \ab[24][64] , \ab[24][63] , \ab[24][62] , \ab[24][61] ,
         \ab[24][60] , \ab[24][59] , \ab[24][58] , \ab[24][57] , \ab[24][56] ,
         \ab[24][55] , \ab[24][54] , \ab[24][53] , \ab[24][52] , \ab[24][51] ,
         \ab[24][50] , \ab[24][49] , \ab[24][48] , \ab[24][47] , \ab[24][46] ,
         \ab[24][45] , \ab[24][44] , \ab[24][43] , \ab[24][42] , \ab[24][41] ,
         \ab[24][40] , \ab[24][39] , \ab[24][38] , \ab[24][37] , \ab[24][36] ,
         \ab[24][35] , \ab[24][34] , \ab[24][33] , \ab[24][32] , \ab[24][31] ,
         \ab[24][30] , \ab[24][29] , \ab[24][28] , \ab[24][27] , \ab[24][26] ,
         \ab[24][25] , \ab[24][24] , \ab[24][23] , \ab[24][22] , \ab[24][21] ,
         \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] , \ab[24][16] ,
         \ab[24][15] , \ab[24][14] , \ab[24][13] , \ab[24][12] , \ab[24][11] ,
         \ab[24][10] , \ab[24][9] , \ab[24][8] , \ab[24][7] , \ab[24][6] ,
         \ab[24][5] , \ab[24][4] , \ab[24][3] , \ab[24][2] , \ab[24][1] ,
         \ab[24][0] , \ab[23][95] , \ab[23][94] , \ab[23][93] , \ab[23][92] ,
         \ab[23][91] , \ab[23][90] , \ab[23][89] , \ab[23][88] , \ab[23][87] ,
         \ab[23][86] , \ab[23][85] , \ab[23][84] , \ab[23][83] , \ab[23][82] ,
         \ab[23][81] , \ab[23][80] , \ab[23][79] , \ab[23][78] , \ab[23][77] ,
         \ab[23][76] , \ab[23][75] , \ab[23][74] , \ab[23][73] , \ab[23][72] ,
         \ab[23][71] , \ab[23][70] , \ab[23][69] , \ab[23][68] , \ab[23][67] ,
         \ab[23][66] , \ab[23][65] , \ab[23][64] , \ab[23][63] , \ab[23][62] ,
         \ab[23][61] , \ab[23][60] , \ab[23][59] , \ab[23][58] , \ab[23][57] ,
         \ab[23][56] , \ab[23][55] , \ab[23][54] , \ab[23][53] , \ab[23][52] ,
         \ab[23][51] , \ab[23][50] , \ab[23][49] , \ab[23][48] , \ab[23][47] ,
         \ab[23][46] , \ab[23][45] , \ab[23][44] , \ab[23][43] , \ab[23][42] ,
         \ab[23][41] , \ab[23][40] , \ab[23][39] , \ab[23][38] , \ab[23][37] ,
         \ab[23][36] , \ab[23][35] , \ab[23][34] , \ab[23][33] , \ab[23][32] ,
         \ab[23][31] , \ab[23][30] , \ab[23][29] , \ab[23][28] , \ab[23][27] ,
         \ab[23][26] , \ab[23][25] , \ab[23][24] , \ab[23][23] , \ab[23][22] ,
         \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] , \ab[23][17] ,
         \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] , \ab[23][12] ,
         \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] , \ab[23][7] ,
         \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] , \ab[23][2] ,
         \ab[23][1] , \ab[23][0] , \ab[22][95] , \ab[22][94] , \ab[22][93] ,
         \ab[22][92] , \ab[22][91] , \ab[22][90] , \ab[22][89] , \ab[22][88] ,
         \ab[22][87] , \ab[22][86] , \ab[22][85] , \ab[22][84] , \ab[22][83] ,
         \ab[22][82] , \ab[22][81] , \ab[22][80] , \ab[22][79] , \ab[22][78] ,
         \ab[22][77] , \ab[22][76] , \ab[22][75] , \ab[22][74] , \ab[22][73] ,
         \ab[22][72] , \ab[22][71] , \ab[22][70] , \ab[22][69] , \ab[22][68] ,
         \ab[22][67] , \ab[22][66] , \ab[22][65] , \ab[22][64] , \ab[22][63] ,
         \ab[22][62] , \ab[22][61] , \ab[22][60] , \ab[22][59] , \ab[22][58] ,
         \ab[22][57] , \ab[22][56] , \ab[22][55] , \ab[22][54] , \ab[22][53] ,
         \ab[22][52] , \ab[22][51] , \ab[22][50] , \ab[22][49] , \ab[22][48] ,
         \ab[22][47] , \ab[22][46] , \ab[22][45] , \ab[22][44] , \ab[22][43] ,
         \ab[22][42] , \ab[22][41] , \ab[22][40] , \ab[22][39] , \ab[22][38] ,
         \ab[22][37] , \ab[22][36] , \ab[22][35] , \ab[22][34] , \ab[22][33] ,
         \ab[22][32] , \ab[22][31] , \ab[22][30] , \ab[22][29] , \ab[22][28] ,
         \ab[22][27] , \ab[22][26] , \ab[22][25] , \ab[22][24] , \ab[22][23] ,
         \ab[22][22] , \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] ,
         \ab[22][17] , \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] ,
         \ab[22][12] , \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] ,
         \ab[22][7] , \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] ,
         \ab[22][2] , \ab[22][1] , \ab[22][0] , \ab[21][95] , \ab[21][94] ,
         \ab[21][93] , \ab[21][92] , \ab[21][91] , \ab[21][90] , \ab[21][89] ,
         \ab[21][88] , \ab[21][87] , \ab[21][86] , \ab[21][85] , \ab[21][84] ,
         \ab[21][83] , \ab[21][82] , \ab[21][81] , \ab[21][80] , \ab[21][79] ,
         \ab[21][78] , \ab[21][77] , \ab[21][76] , \ab[21][75] , \ab[21][74] ,
         \ab[21][73] , \ab[21][72] , \ab[21][71] , \ab[21][70] , \ab[21][69] ,
         \ab[21][68] , \ab[21][67] , \ab[21][66] , \ab[21][65] , \ab[21][64] ,
         \ab[21][63] , \ab[21][62] , \ab[21][61] , \ab[21][60] , \ab[21][59] ,
         \ab[21][58] , \ab[21][57] , \ab[21][56] , \ab[21][55] , \ab[21][54] ,
         \ab[21][53] , \ab[21][52] , \ab[21][51] , \ab[21][50] , \ab[21][49] ,
         \ab[21][48] , \ab[21][47] , \ab[21][46] , \ab[21][45] , \ab[21][44] ,
         \ab[21][43] , \ab[21][42] , \ab[21][41] , \ab[21][40] , \ab[21][39] ,
         \ab[21][38] , \ab[21][37] , \ab[21][36] , \ab[21][35] , \ab[21][34] ,
         \ab[21][33] , \ab[21][32] , \ab[21][31] , \ab[21][30] , \ab[21][29] ,
         \ab[21][28] , \ab[21][27] , \ab[21][26] , \ab[21][25] , \ab[21][24] ,
         \ab[21][23] , \ab[21][22] , \ab[21][21] , \ab[21][20] , \ab[21][19] ,
         \ab[21][18] , \ab[21][17] , \ab[21][16] , \ab[21][15] , \ab[21][14] ,
         \ab[21][13] , \ab[21][12] , \ab[21][11] , \ab[21][10] , \ab[21][9] ,
         \ab[21][8] , \ab[21][7] , \ab[21][6] , \ab[21][5] , \ab[21][4] ,
         \ab[21][3] , \ab[21][2] , \ab[21][1] , \ab[21][0] , \ab[20][95] ,
         \ab[20][94] , \ab[20][93] , \ab[20][92] , \ab[20][91] , \ab[20][90] ,
         \ab[20][89] , \ab[20][88] , \ab[20][87] , \ab[20][86] , \ab[20][85] ,
         \ab[20][84] , \ab[20][83] , \ab[20][82] , \ab[20][81] , \ab[20][80] ,
         \ab[20][79] , \ab[20][78] , \ab[20][77] , \ab[20][76] , \ab[20][75] ,
         \ab[20][74] , \ab[20][73] , \ab[20][72] , \ab[20][71] , \ab[20][70] ,
         \ab[20][69] , \ab[20][68] , \ab[20][67] , \ab[20][66] , \ab[20][65] ,
         \ab[20][64] , \ab[20][63] , \ab[20][62] , \ab[20][61] , \ab[20][60] ,
         \ab[20][59] , \ab[20][58] , \ab[20][57] , \ab[20][56] , \ab[20][55] ,
         \ab[20][54] , \ab[20][53] , \ab[20][52] , \ab[20][51] , \ab[20][50] ,
         \ab[20][49] , \ab[20][48] , \ab[20][47] , \ab[20][46] , \ab[20][45] ,
         \ab[20][44] , \ab[20][43] , \ab[20][42] , \ab[20][41] , \ab[20][40] ,
         \ab[20][39] , \ab[20][38] , \ab[20][37] , \ab[20][36] , \ab[20][35] ,
         \ab[20][34] , \ab[20][33] , \ab[20][32] , \ab[20][31] , \ab[20][30] ,
         \ab[20][29] , \ab[20][28] , \ab[20][27] , \ab[20][26] , \ab[20][25] ,
         \ab[20][24] , \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] ,
         \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] ,
         \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] ,
         \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] ,
         \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] ,
         \ab[19][95] , \ab[19][94] , \ab[19][93] , \ab[19][92] , \ab[19][91] ,
         \ab[19][90] , \ab[19][89] , \ab[19][88] , \ab[19][87] , \ab[19][86] ,
         \ab[19][85] , \ab[19][84] , \ab[19][83] , \ab[19][82] , \ab[19][81] ,
         \ab[19][80] , \ab[19][79] , \ab[19][78] , \ab[19][77] , \ab[19][76] ,
         \ab[19][75] , \ab[19][74] , \ab[19][73] , \ab[19][72] , \ab[19][71] ,
         \ab[19][70] , \ab[19][69] , \ab[19][68] , \ab[19][67] , \ab[19][66] ,
         \ab[19][65] , \ab[19][64] , \ab[19][63] , \ab[19][62] , \ab[19][61] ,
         \ab[19][60] , \ab[19][59] , \ab[19][58] , \ab[19][57] , \ab[19][56] ,
         \ab[19][55] , \ab[19][54] , \ab[19][53] , \ab[19][52] , \ab[19][51] ,
         \ab[19][50] , \ab[19][49] , \ab[19][48] , \ab[19][47] , \ab[19][46] ,
         \ab[19][45] , \ab[19][44] , \ab[19][43] , \ab[19][42] , \ab[19][41] ,
         \ab[19][40] , \ab[19][39] , \ab[19][38] , \ab[19][37] , \ab[19][36] ,
         \ab[19][35] , \ab[19][34] , \ab[19][33] , \ab[19][32] , \ab[19][31] ,
         \ab[19][30] , \ab[19][29] , \ab[19][28] , \ab[19][27] , \ab[19][26] ,
         \ab[19][25] , \ab[19][24] , \ab[19][23] , \ab[19][22] , \ab[19][21] ,
         \ab[19][20] , \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] ,
         \ab[19][15] , \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] ,
         \ab[19][10] , \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] ,
         \ab[19][5] , \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] ,
         \ab[19][0] , \ab[18][95] , \ab[18][94] , \ab[18][93] , \ab[18][92] ,
         \ab[18][91] , \ab[18][90] , \ab[18][89] , \ab[18][88] , \ab[18][87] ,
         \ab[18][86] , \ab[18][85] , \ab[18][84] , \ab[18][83] , \ab[18][82] ,
         \ab[18][81] , \ab[18][80] , \ab[18][79] , \ab[18][78] , \ab[18][77] ,
         \ab[18][76] , \ab[18][75] , \ab[18][74] , \ab[18][73] , \ab[18][72] ,
         \ab[18][71] , \ab[18][70] , \ab[18][69] , \ab[18][68] , \ab[18][67] ,
         \ab[18][66] , \ab[18][65] , \ab[18][64] , \ab[18][63] , \ab[18][62] ,
         \ab[18][61] , \ab[18][60] , \ab[18][59] , \ab[18][58] , \ab[18][57] ,
         \ab[18][56] , \ab[18][55] , \ab[18][54] , \ab[18][53] , \ab[18][52] ,
         \ab[18][51] , \ab[18][50] , \ab[18][49] , \ab[18][48] , \ab[18][47] ,
         \ab[18][46] , \ab[18][45] , \ab[18][44] , \ab[18][43] , \ab[18][42] ,
         \ab[18][41] , \ab[18][40] , \ab[18][39] , \ab[18][38] , \ab[18][37] ,
         \ab[18][36] , \ab[18][35] , \ab[18][34] , \ab[18][33] , \ab[18][32] ,
         \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] , \ab[18][27] ,
         \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] , \ab[18][22] ,
         \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] , \ab[18][17] ,
         \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] , \ab[18][12] ,
         \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] , \ab[18][7] ,
         \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] , \ab[18][2] ,
         \ab[18][1] , \ab[18][0] , \ab[17][95] , \ab[17][94] , \ab[17][93] ,
         \ab[17][92] , \ab[17][91] , \ab[17][90] , \ab[17][89] , \ab[17][88] ,
         \ab[17][87] , \ab[17][86] , \ab[17][85] , \ab[17][84] , \ab[17][83] ,
         \ab[17][82] , \ab[17][81] , \ab[17][80] , \ab[17][79] , \ab[17][78] ,
         \ab[17][77] , \ab[17][76] , \ab[17][75] , \ab[17][74] , \ab[17][73] ,
         \ab[17][72] , \ab[17][71] , \ab[17][70] , \ab[17][69] , \ab[17][68] ,
         \ab[17][67] , \ab[17][66] , \ab[17][65] , \ab[17][64] , \ab[17][63] ,
         \ab[17][62] , \ab[17][61] , \ab[17][60] , \ab[17][59] , \ab[17][58] ,
         \ab[17][57] , \ab[17][56] , \ab[17][55] , \ab[17][54] , \ab[17][53] ,
         \ab[17][52] , \ab[17][51] , \ab[17][50] , \ab[17][49] , \ab[17][48] ,
         \ab[17][47] , \ab[17][46] , \ab[17][45] , \ab[17][44] , \ab[17][43] ,
         \ab[17][42] , \ab[17][41] , \ab[17][40] , \ab[17][39] , \ab[17][38] ,
         \ab[17][37] , \ab[17][36] , \ab[17][35] , \ab[17][34] , \ab[17][33] ,
         \ab[17][32] , \ab[17][31] , \ab[17][30] , \ab[17][29] , \ab[17][28] ,
         \ab[17][27] , \ab[17][26] , \ab[17][25] , \ab[17][24] , \ab[17][23] ,
         \ab[17][22] , \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] ,
         \ab[17][17] , \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] ,
         \ab[17][12] , \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] ,
         \ab[17][7] , \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] ,
         \ab[17][2] , \ab[17][1] , \ab[17][0] , \ab[16][95] , \ab[16][94] ,
         \ab[16][93] , \ab[16][92] , \ab[16][91] , \ab[16][90] , \ab[16][89] ,
         \ab[16][88] , \ab[16][87] , \ab[16][86] , \ab[16][85] , \ab[16][84] ,
         \ab[16][83] , \ab[16][82] , \ab[16][81] , \ab[16][80] , \ab[16][79] ,
         \ab[16][78] , \ab[16][77] , \ab[16][76] , \ab[16][75] , \ab[16][74] ,
         \ab[16][73] , \ab[16][72] , \ab[16][71] , \ab[16][70] , \ab[16][69] ,
         \ab[16][68] , \ab[16][67] , \ab[16][66] , \ab[16][65] , \ab[16][64] ,
         \ab[16][63] , \ab[16][62] , \ab[16][61] , \ab[16][60] , \ab[16][59] ,
         \ab[16][58] , \ab[16][57] , \ab[16][56] , \ab[16][55] , \ab[16][54] ,
         \ab[16][53] , \ab[16][52] , \ab[16][51] , \ab[16][50] , \ab[16][49] ,
         \ab[16][48] , \ab[16][47] , \ab[16][46] , \ab[16][45] , \ab[16][44] ,
         \ab[16][43] , \ab[16][42] , \ab[16][41] , \ab[16][40] , \ab[16][39] ,
         \ab[16][38] , \ab[16][37] , \ab[16][36] , \ab[16][35] , \ab[16][34] ,
         \ab[16][33] , \ab[16][32] , \ab[16][31] , \ab[16][30] , \ab[16][29] ,
         \ab[16][28] , \ab[16][27] , \ab[16][26] , \ab[16][25] , \ab[16][24] ,
         \ab[16][23] , \ab[16][22] , \ab[16][21] , \ab[16][20] , \ab[16][19] ,
         \ab[16][18] , \ab[16][17] , \ab[16][16] , \ab[16][15] , \ab[16][14] ,
         \ab[16][13] , \ab[16][12] , \ab[16][11] , \ab[16][10] , \ab[16][9] ,
         \ab[16][8] , \ab[16][7] , \ab[16][6] , \ab[16][5] , \ab[16][4] ,
         \ab[16][3] , \ab[16][2] , \ab[16][1] , \ab[16][0] , \ab[15][95] ,
         \ab[15][94] , \ab[15][93] , \ab[15][92] , \ab[15][91] , \ab[15][90] ,
         \ab[15][89] , \ab[15][88] , \ab[15][87] , \ab[15][86] , \ab[15][85] ,
         \ab[15][84] , \ab[15][83] , \ab[15][82] , \ab[15][81] , \ab[15][80] ,
         \ab[15][79] , \ab[15][78] , \ab[15][77] , \ab[15][76] , \ab[15][75] ,
         \ab[15][74] , \ab[15][73] , \ab[15][72] , \ab[15][71] , \ab[15][70] ,
         \ab[15][69] , \ab[15][68] , \ab[15][67] , \ab[15][66] , \ab[15][65] ,
         \ab[15][64] , \ab[15][63] , \ab[15][62] , \ab[15][61] , \ab[15][60] ,
         \ab[15][59] , \ab[15][58] , \ab[15][57] , \ab[15][56] , \ab[15][55] ,
         \ab[15][54] , \ab[15][53] , \ab[15][52] , \ab[15][51] , \ab[15][50] ,
         \ab[15][49] , \ab[15][48] , \ab[15][47] , \ab[15][46] , \ab[15][45] ,
         \ab[15][44] , \ab[15][43] , \ab[15][42] , \ab[15][41] , \ab[15][40] ,
         \ab[15][39] , \ab[15][38] , \ab[15][37] , \ab[15][36] , \ab[15][35] ,
         \ab[15][34] , \ab[15][33] , \ab[15][32] , \ab[15][31] , \ab[15][30] ,
         \ab[15][29] , \ab[15][28] , \ab[15][27] , \ab[15][26] , \ab[15][25] ,
         \ab[15][24] , \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] ,
         \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] ,
         \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] ,
         \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] ,
         \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] ,
         \ab[14][95] , \ab[14][94] , \ab[14][93] , \ab[14][92] , \ab[14][91] ,
         \ab[14][90] , \ab[14][89] , \ab[14][88] , \ab[14][87] , \ab[14][86] ,
         \ab[14][85] , \ab[14][84] , \ab[14][83] , \ab[14][82] , \ab[14][81] ,
         \ab[14][80] , \ab[14][79] , \ab[14][78] , \ab[14][77] , \ab[14][76] ,
         \ab[14][75] , \ab[14][74] , \ab[14][73] , \ab[14][72] , \ab[14][71] ,
         \ab[14][70] , \ab[14][69] , \ab[14][68] , \ab[14][67] , \ab[14][66] ,
         \ab[14][65] , \ab[14][64] , \ab[14][63] , \ab[14][62] , \ab[14][61] ,
         \ab[14][60] , \ab[14][59] , \ab[14][58] , \ab[14][57] , \ab[14][56] ,
         \ab[14][55] , \ab[14][54] , \ab[14][53] , \ab[14][52] , \ab[14][51] ,
         \ab[14][50] , \ab[14][49] , \ab[14][48] , \ab[14][47] , \ab[14][46] ,
         \ab[14][45] , \ab[14][44] , \ab[14][43] , \ab[14][42] , \ab[14][41] ,
         \ab[14][40] , \ab[14][39] , \ab[14][38] , \ab[14][37] , \ab[14][36] ,
         \ab[14][35] , \ab[14][34] , \ab[14][33] , \ab[14][32] , \ab[14][31] ,
         \ab[14][30] , \ab[14][29] , \ab[14][28] , \ab[14][27] , \ab[14][26] ,
         \ab[14][25] , \ab[14][24] , \ab[14][23] , \ab[14][22] , \ab[14][21] ,
         \ab[14][20] , \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] ,
         \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] ,
         \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] ,
         \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] ,
         \ab[14][0] , \ab[13][95] , \ab[13][94] , \ab[13][93] , \ab[13][92] ,
         \ab[13][91] , \ab[13][90] , \ab[13][89] , \ab[13][88] , \ab[13][87] ,
         \ab[13][86] , \ab[13][85] , \ab[13][84] , \ab[13][83] , \ab[13][82] ,
         \ab[13][81] , \ab[13][80] , \ab[13][79] , \ab[13][78] , \ab[13][77] ,
         \ab[13][76] , \ab[13][75] , \ab[13][74] , \ab[13][73] , \ab[13][72] ,
         \ab[13][71] , \ab[13][70] , \ab[13][69] , \ab[13][68] , \ab[13][67] ,
         \ab[13][66] , \ab[13][65] , \ab[13][64] , \ab[13][63] , \ab[13][62] ,
         \ab[13][61] , \ab[13][60] , \ab[13][59] , \ab[13][58] , \ab[13][57] ,
         \ab[13][56] , \ab[13][55] , \ab[13][54] , \ab[13][53] , \ab[13][52] ,
         \ab[13][51] , \ab[13][50] , \ab[13][49] , \ab[13][48] , \ab[13][47] ,
         \ab[13][46] , \ab[13][45] , \ab[13][44] , \ab[13][43] , \ab[13][42] ,
         \ab[13][41] , \ab[13][40] , \ab[13][39] , \ab[13][38] , \ab[13][37] ,
         \ab[13][36] , \ab[13][35] , \ab[13][34] , \ab[13][33] , \ab[13][32] ,
         \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] , \ab[13][27] ,
         \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] , \ab[13][22] ,
         \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] , \ab[13][17] ,
         \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] , \ab[13][12] ,
         \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] , \ab[13][7] ,
         \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] , \ab[13][2] ,
         \ab[13][1] , \ab[13][0] , \ab[12][95] , \ab[12][94] , \ab[12][93] ,
         \ab[12][92] , \ab[12][91] , \ab[12][90] , \ab[12][89] , \ab[12][88] ,
         \ab[12][87] , \ab[12][86] , \ab[12][85] , \ab[12][84] , \ab[12][83] ,
         \ab[12][82] , \ab[12][81] , \ab[12][80] , \ab[12][79] , \ab[12][78] ,
         \ab[12][77] , \ab[12][76] , \ab[12][75] , \ab[12][74] , \ab[12][73] ,
         \ab[12][72] , \ab[12][71] , \ab[12][70] , \ab[12][69] , \ab[12][68] ,
         \ab[12][67] , \ab[12][66] , \ab[12][65] , \ab[12][64] , \ab[12][63] ,
         \ab[12][62] , \ab[12][61] , \ab[12][60] , \ab[12][59] , \ab[12][58] ,
         \ab[12][57] , \ab[12][56] , \ab[12][55] , \ab[12][54] , \ab[12][53] ,
         \ab[12][52] , \ab[12][51] , \ab[12][50] , \ab[12][49] , \ab[12][48] ,
         \ab[12][47] , \ab[12][46] , \ab[12][45] , \ab[12][44] , \ab[12][43] ,
         \ab[12][42] , \ab[12][41] , \ab[12][40] , \ab[12][39] , \ab[12][38] ,
         \ab[12][37] , \ab[12][36] , \ab[12][35] , \ab[12][34] , \ab[12][33] ,
         \ab[12][32] , \ab[12][31] , \ab[12][30] , \ab[12][29] , \ab[12][28] ,
         \ab[12][27] , \ab[12][26] , \ab[12][25] , \ab[12][24] , \ab[12][23] ,
         \ab[12][22] , \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] ,
         \ab[12][17] , \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] ,
         \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] ,
         \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] ,
         \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][95] , \ab[11][94] ,
         \ab[11][93] , \ab[11][92] , \ab[11][91] , \ab[11][90] , \ab[11][89] ,
         \ab[11][88] , \ab[11][87] , \ab[11][86] , \ab[11][85] , \ab[11][84] ,
         \ab[11][83] , \ab[11][82] , \ab[11][81] , \ab[11][80] , \ab[11][79] ,
         \ab[11][78] , \ab[11][77] , \ab[11][76] , \ab[11][75] , \ab[11][74] ,
         \ab[11][73] , \ab[11][72] , \ab[11][71] , \ab[11][70] , \ab[11][69] ,
         \ab[11][68] , \ab[11][67] , \ab[11][66] , \ab[11][65] , \ab[11][64] ,
         \ab[11][63] , \ab[11][62] , \ab[11][61] , \ab[11][60] , \ab[11][59] ,
         \ab[11][58] , \ab[11][57] , \ab[11][56] , \ab[11][55] , \ab[11][54] ,
         \ab[11][53] , \ab[11][52] , \ab[11][51] , \ab[11][50] , \ab[11][49] ,
         \ab[11][48] , \ab[11][47] , \ab[11][46] , \ab[11][45] , \ab[11][44] ,
         \ab[11][43] , \ab[11][42] , \ab[11][41] , \ab[11][40] , \ab[11][39] ,
         \ab[11][38] , \ab[11][37] , \ab[11][36] , \ab[11][35] , \ab[11][34] ,
         \ab[11][33] , \ab[11][32] , \ab[11][31] , \ab[11][30] , \ab[11][29] ,
         \ab[11][28] , \ab[11][27] , \ab[11][26] , \ab[11][25] , \ab[11][24] ,
         \ab[11][23] , \ab[11][22] , \ab[11][21] , \ab[11][20] , \ab[11][19] ,
         \ab[11][18] , \ab[11][17] , \ab[11][16] , \ab[11][15] , \ab[11][14] ,
         \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][95] ,
         \ab[10][94] , \ab[10][93] , \ab[10][92] , \ab[10][91] , \ab[10][90] ,
         \ab[10][89] , \ab[10][88] , \ab[10][87] , \ab[10][86] , \ab[10][85] ,
         \ab[10][84] , \ab[10][83] , \ab[10][82] , \ab[10][81] , \ab[10][80] ,
         \ab[10][79] , \ab[10][78] , \ab[10][77] , \ab[10][76] , \ab[10][75] ,
         \ab[10][74] , \ab[10][73] , \ab[10][72] , \ab[10][71] , \ab[10][70] ,
         \ab[10][69] , \ab[10][68] , \ab[10][67] , \ab[10][66] , \ab[10][65] ,
         \ab[10][64] , \ab[10][63] , \ab[10][62] , \ab[10][61] , \ab[10][60] ,
         \ab[10][59] , \ab[10][58] , \ab[10][57] , \ab[10][56] , \ab[10][55] ,
         \ab[10][54] , \ab[10][53] , \ab[10][52] , \ab[10][51] , \ab[10][50] ,
         \ab[10][49] , \ab[10][48] , \ab[10][47] , \ab[10][46] , \ab[10][45] ,
         \ab[10][44] , \ab[10][43] , \ab[10][42] , \ab[10][41] , \ab[10][40] ,
         \ab[10][39] , \ab[10][38] , \ab[10][37] , \ab[10][36] , \ab[10][35] ,
         \ab[10][34] , \ab[10][33] , \ab[10][32] , \ab[10][31] , \ab[10][30] ,
         \ab[10][29] , \ab[10][28] , \ab[10][27] , \ab[10][26] , \ab[10][25] ,
         \ab[10][24] , \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] ,
         \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][95] , \ab[9][94] , \ab[9][93] , \ab[9][92] , \ab[9][91] ,
         \ab[9][90] , \ab[9][89] , \ab[9][88] , \ab[9][87] , \ab[9][86] ,
         \ab[9][85] , \ab[9][84] , \ab[9][83] , \ab[9][82] , \ab[9][81] ,
         \ab[9][80] , \ab[9][79] , \ab[9][78] , \ab[9][77] , \ab[9][76] ,
         \ab[9][75] , \ab[9][74] , \ab[9][73] , \ab[9][72] , \ab[9][71] ,
         \ab[9][70] , \ab[9][69] , \ab[9][68] , \ab[9][67] , \ab[9][66] ,
         \ab[9][65] , \ab[9][64] , \ab[9][63] , \ab[9][62] , \ab[9][61] ,
         \ab[9][60] , \ab[9][59] , \ab[9][58] , \ab[9][57] , \ab[9][56] ,
         \ab[9][55] , \ab[9][54] , \ab[9][53] , \ab[9][52] , \ab[9][51] ,
         \ab[9][50] , \ab[9][49] , \ab[9][48] , \ab[9][47] , \ab[9][46] ,
         \ab[9][45] , \ab[9][44] , \ab[9][43] , \ab[9][42] , \ab[9][41] ,
         \ab[9][40] , \ab[9][39] , \ab[9][38] , \ab[9][37] , \ab[9][36] ,
         \ab[9][35] , \ab[9][34] , \ab[9][33] , \ab[9][32] , \ab[9][31] ,
         \ab[9][30] , \ab[9][29] , \ab[9][28] , \ab[9][27] , \ab[9][26] ,
         \ab[9][25] , \ab[9][24] , \ab[9][23] , \ab[9][22] , \ab[9][21] ,
         \ab[9][20] , \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] ,
         \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] ,
         \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] ,
         \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] ,
         \ab[9][0] , \ab[8][95] , \ab[8][94] , \ab[8][93] , \ab[8][92] ,
         \ab[8][91] , \ab[8][90] , \ab[8][89] , \ab[8][88] , \ab[8][87] ,
         \ab[8][86] , \ab[8][85] , \ab[8][84] , \ab[8][83] , \ab[8][82] ,
         \ab[8][81] , \ab[8][80] , \ab[8][79] , \ab[8][78] , \ab[8][77] ,
         \ab[8][76] , \ab[8][75] , \ab[8][74] , \ab[8][73] , \ab[8][72] ,
         \ab[8][71] , \ab[8][70] , \ab[8][69] , \ab[8][68] , \ab[8][67] ,
         \ab[8][66] , \ab[8][65] , \ab[8][64] , \ab[8][63] , \ab[8][62] ,
         \ab[8][61] , \ab[8][60] , \ab[8][59] , \ab[8][58] , \ab[8][57] ,
         \ab[8][56] , \ab[8][55] , \ab[8][54] , \ab[8][53] , \ab[8][52] ,
         \ab[8][51] , \ab[8][50] , \ab[8][49] , \ab[8][48] , \ab[8][47] ,
         \ab[8][46] , \ab[8][45] , \ab[8][44] , \ab[8][43] , \ab[8][42] ,
         \ab[8][41] , \ab[8][40] , \ab[8][39] , \ab[8][38] , \ab[8][37] ,
         \ab[8][36] , \ab[8][35] , \ab[8][34] , \ab[8][33] , \ab[8][32] ,
         \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] , \ab[8][27] ,
         \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] , \ab[8][22] ,
         \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] , \ab[8][17] ,
         \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] , \ab[8][12] ,
         \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] ,
         \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] ,
         \ab[8][1] , \ab[8][0] , \ab[7][95] , \ab[7][94] , \ab[7][93] ,
         \ab[7][92] , \ab[7][91] , \ab[7][90] , \ab[7][89] , \ab[7][88] ,
         \ab[7][87] , \ab[7][86] , \ab[7][85] , \ab[7][84] , \ab[7][83] ,
         \ab[7][82] , \ab[7][81] , \ab[7][80] , \ab[7][79] , \ab[7][78] ,
         \ab[7][77] , \ab[7][76] , \ab[7][75] , \ab[7][74] , \ab[7][73] ,
         \ab[7][72] , \ab[7][71] , \ab[7][70] , \ab[7][69] , \ab[7][68] ,
         \ab[7][67] , \ab[7][66] , \ab[7][65] , \ab[7][64] , \ab[7][63] ,
         \ab[7][62] , \ab[7][61] , \ab[7][60] , \ab[7][59] , \ab[7][58] ,
         \ab[7][57] , \ab[7][56] , \ab[7][55] , \ab[7][54] , \ab[7][53] ,
         \ab[7][52] , \ab[7][51] , \ab[7][50] , \ab[7][49] , \ab[7][48] ,
         \ab[7][47] , \ab[7][46] , \ab[7][45] , \ab[7][44] , \ab[7][43] ,
         \ab[7][42] , \ab[7][41] , \ab[7][40] , \ab[7][39] , \ab[7][38] ,
         \ab[7][37] , \ab[7][36] , \ab[7][35] , \ab[7][34] , \ab[7][33] ,
         \ab[7][32] , \ab[7][31] , \ab[7][30] , \ab[7][29] , \ab[7][28] ,
         \ab[7][27] , \ab[7][26] , \ab[7][25] , \ab[7][24] , \ab[7][23] ,
         \ab[7][22] , \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] ,
         \ab[7][17] , \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] ,
         \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] ,
         \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][95] , \ab[6][94] ,
         \ab[6][93] , \ab[6][92] , \ab[6][91] , \ab[6][90] , \ab[6][89] ,
         \ab[6][88] , \ab[6][87] , \ab[6][86] , \ab[6][85] , \ab[6][84] ,
         \ab[6][83] , \ab[6][82] , \ab[6][81] , \ab[6][80] , \ab[6][79] ,
         \ab[6][78] , \ab[6][77] , \ab[6][76] , \ab[6][75] , \ab[6][74] ,
         \ab[6][73] , \ab[6][72] , \ab[6][71] , \ab[6][70] , \ab[6][69] ,
         \ab[6][68] , \ab[6][67] , \ab[6][66] , \ab[6][65] , \ab[6][64] ,
         \ab[6][63] , \ab[6][62] , \ab[6][61] , \ab[6][60] , \ab[6][59] ,
         \ab[6][58] , \ab[6][57] , \ab[6][56] , \ab[6][55] , \ab[6][54] ,
         \ab[6][53] , \ab[6][52] , \ab[6][51] , \ab[6][50] , \ab[6][49] ,
         \ab[6][48] , \ab[6][47] , \ab[6][46] , \ab[6][45] , \ab[6][44] ,
         \ab[6][43] , \ab[6][42] , \ab[6][41] , \ab[6][40] , \ab[6][39] ,
         \ab[6][38] , \ab[6][37] , \ab[6][36] , \ab[6][35] , \ab[6][34] ,
         \ab[6][33] , \ab[6][32] , \ab[6][31] , \ab[6][30] , \ab[6][29] ,
         \ab[6][28] , \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] ,
         \ab[6][23] , \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] ,
         \ab[6][18] , \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][95] ,
         \ab[5][94] , \ab[5][93] , \ab[5][92] , \ab[5][91] , \ab[5][90] ,
         \ab[5][89] , \ab[5][88] , \ab[5][87] , \ab[5][86] , \ab[5][85] ,
         \ab[5][84] , \ab[5][83] , \ab[5][82] , \ab[5][81] , \ab[5][80] ,
         \ab[5][79] , \ab[5][78] , \ab[5][77] , \ab[5][76] , \ab[5][75] ,
         \ab[5][74] , \ab[5][73] , \ab[5][72] , \ab[5][71] , \ab[5][70] ,
         \ab[5][69] , \ab[5][68] , \ab[5][67] , \ab[5][66] , \ab[5][65] ,
         \ab[5][64] , \ab[5][63] , \ab[5][62] , \ab[5][61] , \ab[5][60] ,
         \ab[5][59] , \ab[5][58] , \ab[5][57] , \ab[5][56] , \ab[5][55] ,
         \ab[5][54] , \ab[5][53] , \ab[5][52] , \ab[5][51] , \ab[5][50] ,
         \ab[5][49] , \ab[5][48] , \ab[5][47] , \ab[5][46] , \ab[5][45] ,
         \ab[5][44] , \ab[5][43] , \ab[5][42] , \ab[5][41] , \ab[5][40] ,
         \ab[5][39] , \ab[5][38] , \ab[5][37] , \ab[5][36] , \ab[5][35] ,
         \ab[5][34] , \ab[5][33] , \ab[5][32] , \ab[5][31] , \ab[5][30] ,
         \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] , \ab[5][25] ,
         \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] ,
         \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][95] , \ab[4][94] , \ab[4][93] , \ab[4][92] , \ab[4][91] ,
         \ab[4][90] , \ab[4][89] , \ab[4][88] , \ab[4][87] , \ab[4][86] ,
         \ab[4][85] , \ab[4][84] , \ab[4][83] , \ab[4][82] , \ab[4][81] ,
         \ab[4][80] , \ab[4][79] , \ab[4][78] , \ab[4][77] , \ab[4][76] ,
         \ab[4][75] , \ab[4][74] , \ab[4][73] , \ab[4][72] , \ab[4][71] ,
         \ab[4][70] , \ab[4][69] , \ab[4][68] , \ab[4][67] , \ab[4][66] ,
         \ab[4][65] , \ab[4][64] , \ab[4][63] , \ab[4][62] , \ab[4][61] ,
         \ab[4][60] , \ab[4][59] , \ab[4][58] , \ab[4][57] , \ab[4][56] ,
         \ab[4][55] , \ab[4][54] , \ab[4][53] , \ab[4][52] , \ab[4][51] ,
         \ab[4][50] , \ab[4][49] , \ab[4][48] , \ab[4][47] , \ab[4][46] ,
         \ab[4][45] , \ab[4][44] , \ab[4][43] , \ab[4][42] , \ab[4][41] ,
         \ab[4][40] , \ab[4][39] , \ab[4][38] , \ab[4][37] , \ab[4][36] ,
         \ab[4][35] , \ab[4][34] , \ab[4][33] , \ab[4][32] , \ab[4][31] ,
         \ab[4][30] , \ab[4][29] , \ab[4][28] , \ab[4][27] , \ab[4][26] ,
         \ab[4][25] , \ab[4][24] , \ab[4][23] , \ab[4][22] , \ab[4][21] ,
         \ab[4][20] , \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] ,
         \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] ,
         \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] ,
         \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] ,
         \ab[4][0] , \ab[3][95] , \ab[3][94] , \ab[3][93] , \ab[3][92] ,
         \ab[3][91] , \ab[3][90] , \ab[3][89] , \ab[3][88] , \ab[3][87] ,
         \ab[3][86] , \ab[3][85] , \ab[3][84] , \ab[3][83] , \ab[3][82] ,
         \ab[3][81] , \ab[3][80] , \ab[3][79] , \ab[3][78] , \ab[3][77] ,
         \ab[3][76] , \ab[3][75] , \ab[3][74] , \ab[3][73] , \ab[3][72] ,
         \ab[3][71] , \ab[3][70] , \ab[3][69] , \ab[3][68] , \ab[3][67] ,
         \ab[3][66] , \ab[3][65] , \ab[3][64] , \ab[3][63] , \ab[3][62] ,
         \ab[3][61] , \ab[3][60] , \ab[3][59] , \ab[3][58] , \ab[3][57] ,
         \ab[3][56] , \ab[3][55] , \ab[3][54] , \ab[3][53] , \ab[3][52] ,
         \ab[3][51] , \ab[3][50] , \ab[3][49] , \ab[3][48] , \ab[3][47] ,
         \ab[3][46] , \ab[3][45] , \ab[3][44] , \ab[3][43] , \ab[3][42] ,
         \ab[3][41] , \ab[3][40] , \ab[3][39] , \ab[3][38] , \ab[3][37] ,
         \ab[3][36] , \ab[3][35] , \ab[3][34] , \ab[3][33] , \ab[3][32] ,
         \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] , \ab[3][27] ,
         \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] , \ab[3][22] ,
         \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] , \ab[3][17] ,
         \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] , \ab[3][12] ,
         \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] ,
         \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] ,
         \ab[3][1] , \ab[3][0] , \ab[2][95] , \ab[2][94] , \ab[2][93] ,
         \ab[2][92] , \ab[2][91] , \ab[2][90] , \ab[2][89] , \ab[2][88] ,
         \ab[2][87] , \ab[2][86] , \ab[2][85] , \ab[2][84] , \ab[2][83] ,
         \ab[2][82] , \ab[2][81] , \ab[2][80] , \ab[2][79] , \ab[2][78] ,
         \ab[2][77] , \ab[2][76] , \ab[2][75] , \ab[2][74] , \ab[2][73] ,
         \ab[2][72] , \ab[2][71] , \ab[2][70] , \ab[2][69] , \ab[2][68] ,
         \ab[2][67] , \ab[2][66] , \ab[2][65] , \ab[2][64] , \ab[2][63] ,
         \ab[2][62] , \ab[2][61] , \ab[2][60] , \ab[2][59] , \ab[2][58] ,
         \ab[2][57] , \ab[2][56] , \ab[2][55] , \ab[2][54] , \ab[2][53] ,
         \ab[2][52] , \ab[2][51] , \ab[2][50] , \ab[2][49] , \ab[2][48] ,
         \ab[2][47] , \ab[2][46] , \ab[2][45] , \ab[2][44] , \ab[2][43] ,
         \ab[2][42] , \ab[2][41] , \ab[2][40] , \ab[2][39] , \ab[2][38] ,
         \ab[2][37] , \ab[2][36] , \ab[2][35] , \ab[2][34] , \ab[2][33] ,
         \ab[2][32] , \ab[2][31] , \ab[2][30] , \ab[2][29] , \ab[2][28] ,
         \ab[2][27] , \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] ,
         \ab[2][22] , \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] ,
         \ab[2][17] , \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] ,
         \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][95] , \ab[1][94] ,
         \ab[1][93] , \ab[1][92] , \ab[1][91] , \ab[1][90] , \ab[1][89] ,
         \ab[1][88] , \ab[1][87] , \ab[1][86] , \ab[1][85] , \ab[1][84] ,
         \ab[1][83] , \ab[1][82] , \ab[1][81] , \ab[1][80] , \ab[1][79] ,
         \ab[1][78] , \ab[1][77] , \ab[1][76] , \ab[1][75] , \ab[1][74] ,
         \ab[1][73] , \ab[1][72] , \ab[1][71] , \ab[1][70] , \ab[1][69] ,
         \ab[1][68] , \ab[1][67] , \ab[1][66] , \ab[1][65] , \ab[1][64] ,
         \ab[1][63] , \ab[1][62] , \ab[1][61] , \ab[1][60] , \ab[1][59] ,
         \ab[1][58] , \ab[1][57] , \ab[1][56] , \ab[1][55] , \ab[1][54] ,
         \ab[1][53] , \ab[1][52] , \ab[1][51] , \ab[1][50] , \ab[1][49] ,
         \ab[1][48] , \ab[1][47] , \ab[1][46] , \ab[1][45] , \ab[1][44] ,
         \ab[1][43] , \ab[1][42] , \ab[1][41] , \ab[1][40] , \ab[1][39] ,
         \ab[1][38] , \ab[1][37] , \ab[1][36] , \ab[1][35] , \ab[1][34] ,
         \ab[1][33] , \ab[1][32] , \ab[1][31] , \ab[1][30] , \ab[1][29] ,
         \ab[1][28] , \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] ,
         \ab[1][23] , \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] ,
         \ab[1][18] , \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[0][95] , \ab[0][94] , \ab[0][93] ,
         \ab[0][92] , \ab[0][91] , \ab[0][90] , \ab[0][89] , \ab[0][88] ,
         \ab[0][87] , \ab[0][86] , \ab[0][85] , \ab[0][84] , \ab[0][83] ,
         \ab[0][82] , \ab[0][81] , \ab[0][80] , \ab[0][79] , \ab[0][78] ,
         \ab[0][77] , \ab[0][76] , \ab[0][75] , \ab[0][74] , \ab[0][73] ,
         \ab[0][72] , \ab[0][71] , \ab[0][70] , \ab[0][69] , \ab[0][68] ,
         \ab[0][67] , \ab[0][66] , \ab[0][65] , \ab[0][64] , \ab[0][63] ,
         \ab[0][62] , \ab[0][61] , \ab[0][60] , \ab[0][59] , \ab[0][58] ,
         \ab[0][57] , \ab[0][56] , \ab[0][55] , \ab[0][54] , \ab[0][53] ,
         \ab[0][52] , \ab[0][51] , \ab[0][50] , \ab[0][49] , \ab[0][48] ,
         \ab[0][47] , \ab[0][46] , \ab[0][45] , \ab[0][44] , \ab[0][43] ,
         \ab[0][42] , \ab[0][41] , \ab[0][40] , \ab[0][39] , \ab[0][38] ,
         \ab[0][37] , \ab[0][36] , \ab[0][35] , \ab[0][34] , \ab[0][33] ,
         \ab[0][32] , \ab[0][31] , \ab[0][30] , \ab[0][29] , \ab[0][28] ,
         \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] , \ab[0][23] ,
         \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] , \ab[0][18] ,
         \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] , \ab[0][13] ,
         \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] , \ab[0][8] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \CARRYB[3][31] , \CARRYB[3][30] , \CARRYB[3][29] ,
         \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] ,
         \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] ,
         \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] ,
         \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][94] , \CARRYB[2][93] , \CARRYB[2][92] ,
         \CARRYB[2][91] , \CARRYB[2][90] , \CARRYB[2][89] , \CARRYB[2][88] ,
         \CARRYB[2][87] , \CARRYB[2][86] , \CARRYB[2][85] , \CARRYB[2][84] ,
         \CARRYB[2][83] , \CARRYB[2][82] , \CARRYB[2][81] , \CARRYB[2][80] ,
         \CARRYB[2][79] , \CARRYB[2][78] , \CARRYB[2][77] , \CARRYB[2][76] ,
         \CARRYB[2][75] , \CARRYB[2][74] , \CARRYB[2][73] , \CARRYB[2][72] ,
         \CARRYB[2][71] , \CARRYB[2][70] , \CARRYB[2][69] , \CARRYB[2][68] ,
         \CARRYB[2][67] , \CARRYB[2][66] , \CARRYB[2][65] , \CARRYB[2][64] ,
         \CARRYB[2][63] , \CARRYB[2][62] , \CARRYB[2][61] , \CARRYB[2][60] ,
         \CARRYB[2][59] , \CARRYB[2][58] , \CARRYB[2][57] , \CARRYB[2][56] ,
         \CARRYB[2][55] , \CARRYB[2][54] , \CARRYB[2][53] , \CARRYB[2][52] ,
         \CARRYB[2][51] , \CARRYB[2][50] , \CARRYB[2][49] , \CARRYB[2][48] ,
         \CARRYB[2][47] , \CARRYB[2][46] , \CARRYB[2][45] , \CARRYB[2][44] ,
         \CARRYB[2][43] , \CARRYB[2][42] , \CARRYB[2][41] , \CARRYB[2][40] ,
         \CARRYB[2][39] , \CARRYB[2][38] , \CARRYB[2][37] , \CARRYB[2][36] ,
         \CARRYB[2][35] , \CARRYB[2][34] , \CARRYB[2][33] , \CARRYB[2][32] ,
         \CARRYB[2][31] , \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] ,
         \CARRYB[2][27] , \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] ,
         \CARRYB[2][23] , \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] ,
         \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] ,
         \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[1][94] , \CARRYB[1][93] , \CARRYB[1][92] , \CARRYB[1][91] ,
         \CARRYB[1][90] , \CARRYB[1][89] , \CARRYB[1][88] , \CARRYB[1][87] ,
         \CARRYB[1][86] , \CARRYB[1][85] , \CARRYB[1][84] , \CARRYB[1][83] ,
         \CARRYB[1][82] , \CARRYB[1][81] , \CARRYB[1][80] , \CARRYB[1][79] ,
         \CARRYB[1][78] , \CARRYB[1][77] , \CARRYB[1][76] , \CARRYB[1][75] ,
         \CARRYB[1][74] , \CARRYB[1][73] , \CARRYB[1][72] , \CARRYB[1][71] ,
         \CARRYB[1][70] , \CARRYB[1][69] , \CARRYB[1][68] , \CARRYB[1][67] ,
         \CARRYB[1][66] , \CARRYB[1][65] , \CARRYB[1][64] , \CARRYB[1][63] ,
         \CARRYB[1][62] , \CARRYB[1][61] , \CARRYB[1][60] , \CARRYB[1][59] ,
         \CARRYB[1][58] , \CARRYB[1][57] , \CARRYB[1][56] , \CARRYB[1][55] ,
         \CARRYB[1][54] , \CARRYB[1][53] , \CARRYB[1][52] , \CARRYB[1][51] ,
         \CARRYB[1][50] , \CARRYB[1][49] , \CARRYB[1][48] , \CARRYB[1][47] ,
         \CARRYB[1][46] , \CARRYB[1][45] , \CARRYB[1][44] , \CARRYB[1][43] ,
         \CARRYB[1][42] , \CARRYB[1][41] , \CARRYB[1][40] , \CARRYB[1][39] ,
         \CARRYB[1][38] , \CARRYB[1][37] , \CARRYB[1][36] , \CARRYB[1][35] ,
         \CARRYB[1][34] , \CARRYB[1][33] , \CARRYB[1][32] , \CARRYB[1][31] ,
         \CARRYB[1][30] , \CARRYB[1][29] , \CARRYB[1][28] , \CARRYB[1][27] ,
         \CARRYB[1][26] , \CARRYB[1][25] , \CARRYB[1][24] , \CARRYB[1][23] ,
         \CARRYB[1][22] , \CARRYB[1][21] , \CARRYB[1][20] , \CARRYB[1][19] ,
         \CARRYB[1][18] , \CARRYB[1][17] , \CARRYB[1][16] , \CARRYB[1][15] ,
         \CARRYB[1][14] , \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] ,
         \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] ,
         \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[3][31] ,
         \SUMB[3][30] , \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] ,
         \SUMB[3][26] , \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] ,
         \SUMB[3][22] , \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] ,
         \SUMB[3][18] , \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] ,
         \SUMB[3][14] , \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] ,
         \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \SUMB[2][94] , \SUMB[2][93] , \SUMB[2][92] , \SUMB[2][91] ,
         \SUMB[2][90] , \SUMB[2][89] , \SUMB[2][88] , \SUMB[2][87] ,
         \SUMB[2][86] , \SUMB[2][85] , \SUMB[2][84] , \SUMB[2][83] ,
         \SUMB[2][82] , \SUMB[2][81] , \SUMB[2][80] , \SUMB[2][79] ,
         \SUMB[2][78] , \SUMB[2][77] , \SUMB[2][76] , \SUMB[2][75] ,
         \SUMB[2][74] , \SUMB[2][73] , \SUMB[2][72] , \SUMB[2][71] ,
         \SUMB[2][70] , \SUMB[2][69] , \SUMB[2][68] , \SUMB[2][67] ,
         \SUMB[2][66] , \SUMB[2][65] , \SUMB[2][64] , \SUMB[2][63] ,
         \SUMB[2][62] , \SUMB[2][61] , \SUMB[2][60] , \SUMB[2][59] ,
         \SUMB[2][58] , \SUMB[2][57] , \SUMB[2][56] , \SUMB[2][55] ,
         \SUMB[2][54] , \SUMB[2][53] , \SUMB[2][52] , \SUMB[2][51] ,
         \SUMB[2][50] , \SUMB[2][49] , \SUMB[2][48] , \SUMB[2][47] ,
         \SUMB[2][46] , \SUMB[2][45] , \SUMB[2][44] , \SUMB[2][43] ,
         \SUMB[2][42] , \SUMB[2][41] , \SUMB[2][40] , \SUMB[2][39] ,
         \SUMB[2][38] , \SUMB[2][37] , \SUMB[2][36] , \SUMB[2][35] ,
         \SUMB[2][34] , \SUMB[2][33] , \SUMB[2][32] , \SUMB[2][31] ,
         \SUMB[2][30] , \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] ,
         \SUMB[2][26] , \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] ,
         \SUMB[2][22] , \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] ,
         \SUMB[2][18] , \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][94] , \SUMB[1][93] , \SUMB[1][92] , \SUMB[1][91] ,
         \SUMB[1][90] , \SUMB[1][89] , \SUMB[1][88] , \SUMB[1][87] ,
         \SUMB[1][86] , \SUMB[1][85] , \SUMB[1][84] , \SUMB[1][83] ,
         \SUMB[1][82] , \SUMB[1][81] , \SUMB[1][80] , \SUMB[1][79] ,
         \SUMB[1][78] , \SUMB[1][77] , \SUMB[1][76] , \SUMB[1][75] ,
         \SUMB[1][74] , \SUMB[1][73] , \SUMB[1][72] , \SUMB[1][71] ,
         \SUMB[1][70] , \SUMB[1][69] , \SUMB[1][68] , \SUMB[1][67] ,
         \SUMB[1][66] , \SUMB[1][65] , \SUMB[1][64] , \SUMB[1][63] ,
         \SUMB[1][62] , \SUMB[1][61] , \SUMB[1][60] , \SUMB[1][59] ,
         \SUMB[1][58] , \SUMB[1][57] , \SUMB[1][56] , \SUMB[1][55] ,
         \SUMB[1][54] , \SUMB[1][53] , \SUMB[1][52] , \SUMB[1][51] ,
         \SUMB[1][50] , \SUMB[1][49] , \SUMB[1][48] , \SUMB[1][47] ,
         \SUMB[1][46] , \SUMB[1][45] , \SUMB[1][44] , \SUMB[1][43] ,
         \SUMB[1][42] , \SUMB[1][41] , \SUMB[1][40] , \SUMB[1][39] ,
         \SUMB[1][38] , \SUMB[1][37] , \SUMB[1][36] , \SUMB[1][35] ,
         \SUMB[1][34] , \SUMB[1][33] , \SUMB[1][32] , \SUMB[1][31] ,
         \SUMB[1][30] , \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] ,
         \SUMB[1][26] , \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] ,
         \SUMB[1][22] , \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] ,
         \SUMB[1][18] , \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] ,
         \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[8][63] , \CARRYB[8][62] , \CARRYB[8][61] , \CARRYB[8][60] ,
         \CARRYB[8][59] , \CARRYB[8][58] , \CARRYB[8][57] , \CARRYB[8][56] ,
         \CARRYB[8][55] , \CARRYB[8][54] , \CARRYB[8][53] , \CARRYB[8][52] ,
         \CARRYB[8][51] , \CARRYB[8][50] , \CARRYB[8][49] , \CARRYB[8][48] ,
         \CARRYB[8][47] , \CARRYB[8][46] , \CARRYB[8][45] , \CARRYB[8][44] ,
         \CARRYB[8][43] , \CARRYB[8][42] , \CARRYB[8][41] , \CARRYB[8][40] ,
         \CARRYB[8][39] , \CARRYB[8][38] , \CARRYB[8][37] , \CARRYB[8][36] ,
         \CARRYB[8][35] , \CARRYB[8][34] , \CARRYB[8][33] , \CARRYB[8][32] ,
         \CARRYB[8][31] , \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] ,
         \CARRYB[8][27] , \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] ,
         \CARRYB[8][23] , \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] ,
         \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] ,
         \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][94] , \CARRYB[7][93] , \CARRYB[7][92] , \CARRYB[7][91] ,
         \CARRYB[7][90] , \CARRYB[7][89] , \CARRYB[7][88] , \CARRYB[7][87] ,
         \CARRYB[7][86] , \CARRYB[7][85] , \CARRYB[7][84] , \CARRYB[7][83] ,
         \CARRYB[7][82] , \CARRYB[7][81] , \CARRYB[7][80] , \CARRYB[7][79] ,
         \CARRYB[7][78] , \CARRYB[7][77] , \CARRYB[7][76] , \CARRYB[7][75] ,
         \CARRYB[7][74] , \CARRYB[7][73] , \CARRYB[7][72] , \CARRYB[7][71] ,
         \CARRYB[7][70] , \CARRYB[7][69] , \CARRYB[7][68] , \CARRYB[7][67] ,
         \CARRYB[7][66] , \CARRYB[7][65] , \CARRYB[7][64] , \CARRYB[7][63] ,
         \CARRYB[7][62] , \CARRYB[7][61] , \CARRYB[7][60] , \CARRYB[7][59] ,
         \CARRYB[7][58] , \CARRYB[7][57] , \CARRYB[7][56] , \CARRYB[7][55] ,
         \CARRYB[7][54] , \CARRYB[7][53] , \CARRYB[7][52] , \CARRYB[7][51] ,
         \CARRYB[7][50] , \CARRYB[7][49] , \CARRYB[7][48] , \CARRYB[7][47] ,
         \CARRYB[7][46] , \CARRYB[7][45] , \CARRYB[7][44] , \CARRYB[7][43] ,
         \CARRYB[7][42] , \CARRYB[7][41] , \CARRYB[7][40] , \CARRYB[7][39] ,
         \CARRYB[7][38] , \CARRYB[7][37] , \CARRYB[7][36] , \CARRYB[7][35] ,
         \CARRYB[7][34] , \CARRYB[7][33] , \CARRYB[7][32] , \CARRYB[7][31] ,
         \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] ,
         \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] ,
         \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] ,
         \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] ,
         \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] ,
         \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] ,
         \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] ,
         \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][94] ,
         \CARRYB[6][93] , \CARRYB[6][92] , \CARRYB[6][91] , \CARRYB[6][90] ,
         \CARRYB[6][89] , \CARRYB[6][88] , \CARRYB[6][87] , \CARRYB[6][86] ,
         \CARRYB[6][85] , \CARRYB[6][84] , \CARRYB[6][83] , \CARRYB[6][82] ,
         \CARRYB[6][81] , \CARRYB[6][80] , \CARRYB[6][79] , \CARRYB[6][78] ,
         \CARRYB[6][77] , \CARRYB[6][76] , \CARRYB[6][75] , \CARRYB[6][74] ,
         \CARRYB[6][73] , \CARRYB[6][72] , \CARRYB[6][71] , \CARRYB[6][70] ,
         \CARRYB[6][69] , \CARRYB[6][68] , \CARRYB[6][67] , \CARRYB[6][66] ,
         \CARRYB[6][65] , \CARRYB[6][64] , \CARRYB[6][63] , \CARRYB[6][62] ,
         \CARRYB[6][61] , \CARRYB[6][60] , \CARRYB[6][59] , \CARRYB[6][58] ,
         \CARRYB[6][57] , \CARRYB[6][56] , \CARRYB[6][55] , \CARRYB[6][54] ,
         \CARRYB[6][53] , \CARRYB[6][52] , \CARRYB[6][51] , \CARRYB[6][50] ,
         \CARRYB[6][49] , \CARRYB[6][48] , \CARRYB[6][47] , \CARRYB[6][46] ,
         \CARRYB[6][45] , \CARRYB[6][44] , \CARRYB[6][43] , \CARRYB[6][42] ,
         \CARRYB[6][41] , \CARRYB[6][40] , \CARRYB[6][39] , \CARRYB[6][38] ,
         \CARRYB[6][37] , \CARRYB[6][36] , \CARRYB[6][35] , \CARRYB[6][34] ,
         \CARRYB[6][33] , \CARRYB[6][32] , \CARRYB[6][31] , \CARRYB[6][30] ,
         \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] ,
         \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] ,
         \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] ,
         \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] ,
         \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] ,
         \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][94] , \CARRYB[5][93] ,
         \CARRYB[5][92] , \CARRYB[5][91] , \CARRYB[5][90] , \CARRYB[5][89] ,
         \CARRYB[5][88] , \CARRYB[5][87] , \CARRYB[5][86] , \CARRYB[5][85] ,
         \CARRYB[5][84] , \CARRYB[5][83] , \CARRYB[5][82] , \CARRYB[5][81] ,
         \CARRYB[5][80] , \CARRYB[5][79] , \CARRYB[5][78] , \CARRYB[5][77] ,
         \CARRYB[5][76] , \CARRYB[5][75] , \CARRYB[5][74] , \CARRYB[5][73] ,
         \CARRYB[5][72] , \CARRYB[5][71] , \CARRYB[5][70] , \CARRYB[5][69] ,
         \CARRYB[5][68] , \CARRYB[5][67] , \CARRYB[5][66] , \CARRYB[5][65] ,
         \CARRYB[5][64] , \CARRYB[5][63] , \CARRYB[5][62] , \CARRYB[5][61] ,
         \CARRYB[5][60] , \CARRYB[5][59] , \CARRYB[5][58] , \CARRYB[5][57] ,
         \CARRYB[5][56] , \CARRYB[5][55] , \CARRYB[5][54] , \CARRYB[5][53] ,
         \CARRYB[5][52] , \CARRYB[5][51] , \CARRYB[5][50] , \CARRYB[5][49] ,
         \CARRYB[5][48] , \CARRYB[5][47] , \CARRYB[5][46] , \CARRYB[5][45] ,
         \CARRYB[5][44] , \CARRYB[5][43] , \CARRYB[5][42] , \CARRYB[5][41] ,
         \CARRYB[5][40] , \CARRYB[5][39] , \CARRYB[5][38] , \CARRYB[5][37] ,
         \CARRYB[5][36] , \CARRYB[5][35] , \CARRYB[5][34] , \CARRYB[5][33] ,
         \CARRYB[5][32] , \CARRYB[5][31] , \CARRYB[5][30] , \CARRYB[5][29] ,
         \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] ,
         \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] ,
         \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] ,
         \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][94] , \CARRYB[4][93] , \CARRYB[4][92] ,
         \CARRYB[4][91] , \CARRYB[4][90] , \CARRYB[4][89] , \CARRYB[4][88] ,
         \CARRYB[4][87] , \CARRYB[4][86] , \CARRYB[4][85] , \CARRYB[4][84] ,
         \CARRYB[4][83] , \CARRYB[4][82] , \CARRYB[4][81] , \CARRYB[4][80] ,
         \CARRYB[4][79] , \CARRYB[4][78] , \CARRYB[4][77] , \CARRYB[4][76] ,
         \CARRYB[4][75] , \CARRYB[4][74] , \CARRYB[4][73] , \CARRYB[4][72] ,
         \CARRYB[4][71] , \CARRYB[4][70] , \CARRYB[4][69] , \CARRYB[4][68] ,
         \CARRYB[4][67] , \CARRYB[4][66] , \CARRYB[4][65] , \CARRYB[4][64] ,
         \CARRYB[4][63] , \CARRYB[4][62] , \CARRYB[4][61] , \CARRYB[4][60] ,
         \CARRYB[4][59] , \CARRYB[4][58] , \CARRYB[4][57] , \CARRYB[4][56] ,
         \CARRYB[4][55] , \CARRYB[4][54] , \CARRYB[4][53] , \CARRYB[4][52] ,
         \CARRYB[4][51] , \CARRYB[4][50] , \CARRYB[4][49] , \CARRYB[4][48] ,
         \CARRYB[4][47] , \CARRYB[4][46] , \CARRYB[4][45] , \CARRYB[4][44] ,
         \CARRYB[4][43] , \CARRYB[4][42] , \CARRYB[4][41] , \CARRYB[4][40] ,
         \CARRYB[4][39] , \CARRYB[4][38] , \CARRYB[4][37] , \CARRYB[4][36] ,
         \CARRYB[4][35] , \CARRYB[4][34] , \CARRYB[4][33] , \CARRYB[4][32] ,
         \CARRYB[4][31] , \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] ,
         \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] ,
         \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] ,
         \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] ,
         \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][94] , \CARRYB[3][93] , \CARRYB[3][92] , \CARRYB[3][91] ,
         \CARRYB[3][90] , \CARRYB[3][89] , \CARRYB[3][88] , \CARRYB[3][87] ,
         \CARRYB[3][86] , \CARRYB[3][85] , \CARRYB[3][84] , \CARRYB[3][83] ,
         \CARRYB[3][82] , \CARRYB[3][81] , \CARRYB[3][80] , \CARRYB[3][79] ,
         \CARRYB[3][78] , \CARRYB[3][77] , \CARRYB[3][76] , \CARRYB[3][75] ,
         \CARRYB[3][74] , \CARRYB[3][73] , \CARRYB[3][72] , \CARRYB[3][71] ,
         \CARRYB[3][70] , \CARRYB[3][69] , \CARRYB[3][68] , \CARRYB[3][67] ,
         \CARRYB[3][66] , \CARRYB[3][65] , \CARRYB[3][64] , \CARRYB[3][63] ,
         \CARRYB[3][62] , \CARRYB[3][61] , \CARRYB[3][60] , \CARRYB[3][59] ,
         \CARRYB[3][58] , \CARRYB[3][57] , \CARRYB[3][56] , \CARRYB[3][55] ,
         \CARRYB[3][54] , \CARRYB[3][53] , \CARRYB[3][52] , \CARRYB[3][51] ,
         \CARRYB[3][50] , \CARRYB[3][49] , \CARRYB[3][48] , \CARRYB[3][47] ,
         \CARRYB[3][46] , \CARRYB[3][45] , \CARRYB[3][44] , \CARRYB[3][43] ,
         \CARRYB[3][42] , \CARRYB[3][41] , \CARRYB[3][40] , \CARRYB[3][39] ,
         \CARRYB[3][38] , \CARRYB[3][37] , \CARRYB[3][36] , \CARRYB[3][35] ,
         \CARRYB[3][34] , \CARRYB[3][33] , \CARRYB[3][32] , \SUMB[8][63] ,
         \SUMB[8][62] , \SUMB[8][61] , \SUMB[8][60] , \SUMB[8][59] ,
         \SUMB[8][58] , \SUMB[8][57] , \SUMB[8][56] , \SUMB[8][55] ,
         \SUMB[8][54] , \SUMB[8][53] , \SUMB[8][52] , \SUMB[8][51] ,
         \SUMB[8][50] , \SUMB[8][49] , \SUMB[8][48] , \SUMB[8][47] ,
         \SUMB[8][46] , \SUMB[8][45] , \SUMB[8][44] , \SUMB[8][43] ,
         \SUMB[8][42] , \SUMB[8][41] , \SUMB[8][40] , \SUMB[8][39] ,
         \SUMB[8][38] , \SUMB[8][37] , \SUMB[8][36] , \SUMB[8][35] ,
         \SUMB[8][34] , \SUMB[8][33] , \SUMB[8][32] , \SUMB[8][31] ,
         \SUMB[8][30] , \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] ,
         \SUMB[8][26] , \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] ,
         \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][94] , \SUMB[7][93] , \SUMB[7][92] , \SUMB[7][91] ,
         \SUMB[7][90] , \SUMB[7][89] , \SUMB[7][88] , \SUMB[7][87] ,
         \SUMB[7][86] , \SUMB[7][85] , \SUMB[7][84] , \SUMB[7][83] ,
         \SUMB[7][82] , \SUMB[7][81] , \SUMB[7][80] , \SUMB[7][79] ,
         \SUMB[7][78] , \SUMB[7][77] , \SUMB[7][76] , \SUMB[7][75] ,
         \SUMB[7][74] , \SUMB[7][73] , \SUMB[7][72] , \SUMB[7][71] ,
         \SUMB[7][70] , \SUMB[7][69] , \SUMB[7][68] , \SUMB[7][67] ,
         \SUMB[7][66] , \SUMB[7][65] , \SUMB[7][64] , \SUMB[7][63] ,
         \SUMB[7][62] , \SUMB[7][61] , \SUMB[7][60] , \SUMB[7][59] ,
         \SUMB[7][58] , \SUMB[7][57] , \SUMB[7][56] , \SUMB[7][55] ,
         \SUMB[7][54] , \SUMB[7][53] , \SUMB[7][52] , \SUMB[7][51] ,
         \SUMB[7][50] , \SUMB[7][49] , \SUMB[7][48] , \SUMB[7][47] ,
         \SUMB[7][46] , \SUMB[7][45] , \SUMB[7][44] , \SUMB[7][43] ,
         \SUMB[7][42] , \SUMB[7][41] , \SUMB[7][40] , \SUMB[7][39] ,
         \SUMB[7][38] , \SUMB[7][37] , \SUMB[7][36] , \SUMB[7][35] ,
         \SUMB[7][34] , \SUMB[7][33] , \SUMB[7][32] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][94] , \SUMB[6][93] , \SUMB[6][92] , \SUMB[6][91] ,
         \SUMB[6][90] , \SUMB[6][89] , \SUMB[6][88] , \SUMB[6][87] ,
         \SUMB[6][86] , \SUMB[6][85] , \SUMB[6][84] , \SUMB[6][83] ,
         \SUMB[6][82] , \SUMB[6][81] , \SUMB[6][80] , \SUMB[6][79] ,
         \SUMB[6][78] , \SUMB[6][77] , \SUMB[6][76] , \SUMB[6][75] ,
         \SUMB[6][74] , \SUMB[6][73] , \SUMB[6][72] , \SUMB[6][71] ,
         \SUMB[6][70] , \SUMB[6][69] , \SUMB[6][68] , \SUMB[6][67] ,
         \SUMB[6][66] , \SUMB[6][65] , \SUMB[6][64] , \SUMB[6][63] ,
         \SUMB[6][62] , \SUMB[6][61] , \SUMB[6][60] , \SUMB[6][59] ,
         \SUMB[6][58] , \SUMB[6][57] , \SUMB[6][56] , \SUMB[6][55] ,
         \SUMB[6][54] , \SUMB[6][53] , \SUMB[6][52] , \SUMB[6][51] ,
         \SUMB[6][50] , \SUMB[6][49] , \SUMB[6][48] , \SUMB[6][47] ,
         \SUMB[6][46] , \SUMB[6][45] , \SUMB[6][44] , \SUMB[6][43] ,
         \SUMB[6][42] , \SUMB[6][41] , \SUMB[6][40] , \SUMB[6][39] ,
         \SUMB[6][38] , \SUMB[6][37] , \SUMB[6][36] , \SUMB[6][35] ,
         \SUMB[6][34] , \SUMB[6][33] , \SUMB[6][32] , \SUMB[6][31] ,
         \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] ,
         \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] ,
         \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] ,
         \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][94] , \SUMB[5][93] , \SUMB[5][92] , \SUMB[5][91] ,
         \SUMB[5][90] , \SUMB[5][89] , \SUMB[5][88] , \SUMB[5][87] ,
         \SUMB[5][86] , \SUMB[5][85] , \SUMB[5][84] , \SUMB[5][83] ,
         \SUMB[5][82] , \SUMB[5][81] , \SUMB[5][80] , \SUMB[5][79] ,
         \SUMB[5][78] , \SUMB[5][77] , \SUMB[5][76] , \SUMB[5][75] ,
         \SUMB[5][74] , \SUMB[5][73] , \SUMB[5][72] , \SUMB[5][71] ,
         \SUMB[5][70] , \SUMB[5][69] , \SUMB[5][68] , \SUMB[5][67] ,
         \SUMB[5][66] , \SUMB[5][65] , \SUMB[5][64] , \SUMB[5][63] ,
         \SUMB[5][62] , \SUMB[5][61] , \SUMB[5][60] , \SUMB[5][59] ,
         \SUMB[5][58] , \SUMB[5][57] , \SUMB[5][56] , \SUMB[5][55] ,
         \SUMB[5][54] , \SUMB[5][53] , \SUMB[5][52] , \SUMB[5][51] ,
         \SUMB[5][50] , \SUMB[5][49] , \SUMB[5][48] , \SUMB[5][47] ,
         \SUMB[5][46] , \SUMB[5][45] , \SUMB[5][44] , \SUMB[5][43] ,
         \SUMB[5][42] , \SUMB[5][41] , \SUMB[5][40] , \SUMB[5][39] ,
         \SUMB[5][38] , \SUMB[5][37] , \SUMB[5][36] , \SUMB[5][35] ,
         \SUMB[5][34] , \SUMB[5][33] , \SUMB[5][32] , \SUMB[5][31] ,
         \SUMB[5][30] , \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] ,
         \SUMB[5][26] , \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] ,
         \SUMB[5][22] , \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] ,
         \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][94] , \SUMB[4][93] , \SUMB[4][92] , \SUMB[4][91] ,
         \SUMB[4][90] , \SUMB[4][89] , \SUMB[4][88] , \SUMB[4][87] ,
         \SUMB[4][86] , \SUMB[4][85] , \SUMB[4][84] , \SUMB[4][83] ,
         \SUMB[4][82] , \SUMB[4][81] , \SUMB[4][80] , \SUMB[4][79] ,
         \SUMB[4][78] , \SUMB[4][77] , \SUMB[4][76] , \SUMB[4][75] ,
         \SUMB[4][74] , \SUMB[4][73] , \SUMB[4][72] , \SUMB[4][71] ,
         \SUMB[4][70] , \SUMB[4][69] , \SUMB[4][68] , \SUMB[4][67] ,
         \SUMB[4][66] , \SUMB[4][65] , \SUMB[4][64] , \SUMB[4][63] ,
         \SUMB[4][62] , \SUMB[4][61] , \SUMB[4][60] , \SUMB[4][59] ,
         \SUMB[4][58] , \SUMB[4][57] , \SUMB[4][56] , \SUMB[4][55] ,
         \SUMB[4][54] , \SUMB[4][53] , \SUMB[4][52] , \SUMB[4][51] ,
         \SUMB[4][50] , \SUMB[4][49] , \SUMB[4][48] , \SUMB[4][47] ,
         \SUMB[4][46] , \SUMB[4][45] , \SUMB[4][44] , \SUMB[4][43] ,
         \SUMB[4][42] , \SUMB[4][41] , \SUMB[4][40] , \SUMB[4][39] ,
         \SUMB[4][38] , \SUMB[4][37] , \SUMB[4][36] , \SUMB[4][35] ,
         \SUMB[4][34] , \SUMB[4][33] , \SUMB[4][32] , \SUMB[4][31] ,
         \SUMB[4][30] , \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] ,
         \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][94] , \SUMB[3][93] , \SUMB[3][92] , \SUMB[3][91] ,
         \SUMB[3][90] , \SUMB[3][89] , \SUMB[3][88] , \SUMB[3][87] ,
         \SUMB[3][86] , \SUMB[3][85] , \SUMB[3][84] , \SUMB[3][83] ,
         \SUMB[3][82] , \SUMB[3][81] , \SUMB[3][80] , \SUMB[3][79] ,
         \SUMB[3][78] , \SUMB[3][77] , \SUMB[3][76] , \SUMB[3][75] ,
         \SUMB[3][74] , \SUMB[3][73] , \SUMB[3][72] , \SUMB[3][71] ,
         \SUMB[3][70] , \SUMB[3][69] , \SUMB[3][68] , \SUMB[3][67] ,
         \SUMB[3][66] , \SUMB[3][65] , \SUMB[3][64] , \SUMB[3][63] ,
         \SUMB[3][62] , \SUMB[3][61] , \SUMB[3][60] , \SUMB[3][59] ,
         \SUMB[3][58] , \SUMB[3][57] , \SUMB[3][56] , \SUMB[3][55] ,
         \SUMB[3][54] , \SUMB[3][53] , \SUMB[3][52] , \SUMB[3][51] ,
         \SUMB[3][50] , \SUMB[3][49] , \SUMB[3][48] , \SUMB[3][47] ,
         \SUMB[3][46] , \SUMB[3][45] , \SUMB[3][44] , \SUMB[3][43] ,
         \SUMB[3][42] , \SUMB[3][41] , \SUMB[3][40] , \SUMB[3][39] ,
         \SUMB[3][38] , \SUMB[3][37] , \SUMB[3][36] , \SUMB[3][35] ,
         \SUMB[3][34] , \SUMB[3][33] , \SUMB[3][32] , \CARRYB[13][94] ,
         \CARRYB[13][93] , \CARRYB[13][92] , \CARRYB[13][91] ,
         \CARRYB[13][90] , \CARRYB[13][89] , \CARRYB[13][88] ,
         \CARRYB[13][87] , \CARRYB[13][86] , \CARRYB[13][85] ,
         \CARRYB[13][84] , \CARRYB[13][83] , \CARRYB[13][82] ,
         \CARRYB[13][81] , \CARRYB[13][80] , \CARRYB[13][79] ,
         \CARRYB[13][78] , \CARRYB[13][77] , \CARRYB[13][76] ,
         \CARRYB[13][75] , \CARRYB[13][74] , \CARRYB[13][73] ,
         \CARRYB[13][72] , \CARRYB[13][71] , \CARRYB[13][70] ,
         \CARRYB[13][69] , \CARRYB[13][68] , \CARRYB[13][67] ,
         \CARRYB[13][66] , \CARRYB[13][65] , \CARRYB[13][64] ,
         \CARRYB[13][63] , \CARRYB[13][62] , \CARRYB[13][61] ,
         \CARRYB[13][60] , \CARRYB[13][59] , \CARRYB[13][58] ,
         \CARRYB[13][57] , \CARRYB[13][56] , \CARRYB[13][55] ,
         \CARRYB[13][54] , \CARRYB[13][53] , \CARRYB[13][52] ,
         \CARRYB[13][51] , \CARRYB[13][50] , \CARRYB[13][49] ,
         \CARRYB[13][48] , \CARRYB[13][47] , \CARRYB[13][46] ,
         \CARRYB[13][45] , \CARRYB[13][44] , \CARRYB[13][43] ,
         \CARRYB[13][42] , \CARRYB[13][41] , \CARRYB[13][40] ,
         \CARRYB[13][39] , \CARRYB[13][38] , \CARRYB[13][37] ,
         \CARRYB[13][36] , \CARRYB[13][35] , \CARRYB[13][34] ,
         \CARRYB[13][33] , \CARRYB[13][32] , \CARRYB[13][31] ,
         \CARRYB[13][30] , \CARRYB[13][29] , \CARRYB[13][28] ,
         \CARRYB[13][27] , \CARRYB[13][26] , \CARRYB[13][25] ,
         \CARRYB[13][24] , \CARRYB[13][23] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][94] , \CARRYB[12][93] , \CARRYB[12][92] ,
         \CARRYB[12][91] , \CARRYB[12][90] , \CARRYB[12][89] ,
         \CARRYB[12][88] , \CARRYB[12][87] , \CARRYB[12][86] ,
         \CARRYB[12][85] , \CARRYB[12][84] , \CARRYB[12][83] ,
         \CARRYB[12][82] , \CARRYB[12][81] , \CARRYB[12][80] ,
         \CARRYB[12][79] , \CARRYB[12][78] , \CARRYB[12][77] ,
         \CARRYB[12][76] , \CARRYB[12][75] , \CARRYB[12][74] ,
         \CARRYB[12][73] , \CARRYB[12][72] , \CARRYB[12][71] ,
         \CARRYB[12][70] , \CARRYB[12][69] , \CARRYB[12][68] ,
         \CARRYB[12][67] , \CARRYB[12][66] , \CARRYB[12][65] ,
         \CARRYB[12][64] , \CARRYB[12][63] , \CARRYB[12][62] ,
         \CARRYB[12][61] , \CARRYB[12][60] , \CARRYB[12][59] ,
         \CARRYB[12][58] , \CARRYB[12][57] , \CARRYB[12][56] ,
         \CARRYB[12][55] , \CARRYB[12][54] , \CARRYB[12][53] ,
         \CARRYB[12][52] , \CARRYB[12][51] , \CARRYB[12][50] ,
         \CARRYB[12][49] , \CARRYB[12][48] , \CARRYB[12][47] ,
         \CARRYB[12][46] , \CARRYB[12][45] , \CARRYB[12][44] ,
         \CARRYB[12][43] , \CARRYB[12][42] , \CARRYB[12][41] ,
         \CARRYB[12][40] , \CARRYB[12][39] , \CARRYB[12][38] ,
         \CARRYB[12][37] , \CARRYB[12][36] , \CARRYB[12][35] ,
         \CARRYB[12][34] , \CARRYB[12][33] , \CARRYB[12][32] ,
         \CARRYB[12][31] , \CARRYB[12][30] , \CARRYB[12][29] ,
         \CARRYB[12][28] , \CARRYB[12][27] , \CARRYB[12][26] ,
         \CARRYB[12][25] , \CARRYB[12][24] , \CARRYB[12][23] ,
         \CARRYB[12][22] , \CARRYB[12][21] , \CARRYB[12][20] ,
         \CARRYB[12][19] , \CARRYB[12][18] , \CARRYB[12][17] ,
         \CARRYB[12][16] , \CARRYB[12][15] , \CARRYB[12][14] ,
         \CARRYB[12][13] , \CARRYB[12][12] , \CARRYB[12][11] ,
         \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] , \CARRYB[12][7] ,
         \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] , \CARRYB[11][94] ,
         \CARRYB[11][93] , \CARRYB[11][92] , \CARRYB[11][91] ,
         \CARRYB[11][90] , \CARRYB[11][89] , \CARRYB[11][88] ,
         \CARRYB[11][87] , \CARRYB[11][86] , \CARRYB[11][85] ,
         \CARRYB[11][84] , \CARRYB[11][83] , \CARRYB[11][82] ,
         \CARRYB[11][81] , \CARRYB[11][80] , \CARRYB[11][79] ,
         \CARRYB[11][78] , \CARRYB[11][77] , \CARRYB[11][76] ,
         \CARRYB[11][75] , \CARRYB[11][74] , \CARRYB[11][73] ,
         \CARRYB[11][72] , \CARRYB[11][71] , \CARRYB[11][70] ,
         \CARRYB[11][69] , \CARRYB[11][68] , \CARRYB[11][67] ,
         \CARRYB[11][66] , \CARRYB[11][65] , \CARRYB[11][64] ,
         \CARRYB[11][63] , \CARRYB[11][62] , \CARRYB[11][61] ,
         \CARRYB[11][60] , \CARRYB[11][59] , \CARRYB[11][58] ,
         \CARRYB[11][57] , \CARRYB[11][56] , \CARRYB[11][55] ,
         \CARRYB[11][54] , \CARRYB[11][53] , \CARRYB[11][52] ,
         \CARRYB[11][51] , \CARRYB[11][50] , \CARRYB[11][49] ,
         \CARRYB[11][48] , \CARRYB[11][47] , \CARRYB[11][46] ,
         \CARRYB[11][45] , \CARRYB[11][44] , \CARRYB[11][43] ,
         \CARRYB[11][42] , \CARRYB[11][41] , \CARRYB[11][40] ,
         \CARRYB[11][39] , \CARRYB[11][38] , \CARRYB[11][37] ,
         \CARRYB[11][36] , \CARRYB[11][35] , \CARRYB[11][34] ,
         \CARRYB[11][33] , \CARRYB[11][32] , \CARRYB[11][31] ,
         \CARRYB[11][30] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][23] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][94] , \CARRYB[10][93] , \CARRYB[10][92] ,
         \CARRYB[10][91] , \CARRYB[10][90] , \CARRYB[10][89] ,
         \CARRYB[10][88] , \CARRYB[10][87] , \CARRYB[10][86] ,
         \CARRYB[10][85] , \CARRYB[10][84] , \CARRYB[10][83] ,
         \CARRYB[10][82] , \CARRYB[10][81] , \CARRYB[10][80] ,
         \CARRYB[10][79] , \CARRYB[10][78] , \CARRYB[10][77] ,
         \CARRYB[10][76] , \CARRYB[10][75] , \CARRYB[10][74] ,
         \CARRYB[10][73] , \CARRYB[10][72] , \CARRYB[10][71] ,
         \CARRYB[10][70] , \CARRYB[10][69] , \CARRYB[10][68] ,
         \CARRYB[10][67] , \CARRYB[10][66] , \CARRYB[10][65] ,
         \CARRYB[10][64] , \CARRYB[10][63] , \CARRYB[10][62] ,
         \CARRYB[10][61] , \CARRYB[10][60] , \CARRYB[10][59] ,
         \CARRYB[10][58] , \CARRYB[10][57] , \CARRYB[10][56] ,
         \CARRYB[10][55] , \CARRYB[10][54] , \CARRYB[10][53] ,
         \CARRYB[10][52] , \CARRYB[10][51] , \CARRYB[10][50] ,
         \CARRYB[10][49] , \CARRYB[10][48] , \CARRYB[10][47] ,
         \CARRYB[10][46] , \CARRYB[10][45] , \CARRYB[10][44] ,
         \CARRYB[10][43] , \CARRYB[10][42] , \CARRYB[10][41] ,
         \CARRYB[10][40] , \CARRYB[10][39] , \CARRYB[10][38] ,
         \CARRYB[10][37] , \CARRYB[10][36] , \CARRYB[10][35] ,
         \CARRYB[10][34] , \CARRYB[10][33] , \CARRYB[10][32] ,
         \CARRYB[10][31] , \CARRYB[10][30] , \CARRYB[10][29] ,
         \CARRYB[10][28] , \CARRYB[10][27] , \CARRYB[10][26] ,
         \CARRYB[10][25] , \CARRYB[10][24] , \CARRYB[10][23] ,
         \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][94] ,
         \CARRYB[9][93] , \CARRYB[9][92] , \CARRYB[9][91] , \CARRYB[9][90] ,
         \CARRYB[9][89] , \CARRYB[9][88] , \CARRYB[9][87] , \CARRYB[9][86] ,
         \CARRYB[9][85] , \CARRYB[9][84] , \CARRYB[9][83] , \CARRYB[9][82] ,
         \CARRYB[9][81] , \CARRYB[9][80] , \CARRYB[9][79] , \CARRYB[9][78] ,
         \CARRYB[9][77] , \CARRYB[9][76] , \CARRYB[9][75] , \CARRYB[9][74] ,
         \CARRYB[9][73] , \CARRYB[9][72] , \CARRYB[9][71] , \CARRYB[9][70] ,
         \CARRYB[9][69] , \CARRYB[9][68] , \CARRYB[9][67] , \CARRYB[9][66] ,
         \CARRYB[9][65] , \CARRYB[9][64] , \CARRYB[9][63] , \CARRYB[9][62] ,
         \CARRYB[9][61] , \CARRYB[9][60] , \CARRYB[9][59] , \CARRYB[9][58] ,
         \CARRYB[9][57] , \CARRYB[9][56] , \CARRYB[9][55] , \CARRYB[9][54] ,
         \CARRYB[9][53] , \CARRYB[9][52] , \CARRYB[9][51] , \CARRYB[9][50] ,
         \CARRYB[9][49] , \CARRYB[9][48] , \CARRYB[9][47] , \CARRYB[9][46] ,
         \CARRYB[9][45] , \CARRYB[9][44] , \CARRYB[9][43] , \CARRYB[9][42] ,
         \CARRYB[9][41] , \CARRYB[9][40] , \CARRYB[9][39] , \CARRYB[9][38] ,
         \CARRYB[9][37] , \CARRYB[9][36] , \CARRYB[9][35] , \CARRYB[9][34] ,
         \CARRYB[9][33] , \CARRYB[9][32] , \CARRYB[9][31] , \CARRYB[9][30] ,
         \CARRYB[9][29] , \CARRYB[9][28] , \CARRYB[9][27] , \CARRYB[9][26] ,
         \CARRYB[9][25] , \CARRYB[9][24] , \CARRYB[9][23] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][94] , \CARRYB[8][93] ,
         \CARRYB[8][92] , \CARRYB[8][91] , \CARRYB[8][90] , \CARRYB[8][89] ,
         \CARRYB[8][88] , \CARRYB[8][87] , \CARRYB[8][86] , \CARRYB[8][85] ,
         \CARRYB[8][84] , \CARRYB[8][83] , \CARRYB[8][82] , \CARRYB[8][81] ,
         \CARRYB[8][80] , \CARRYB[8][79] , \CARRYB[8][78] , \CARRYB[8][77] ,
         \CARRYB[8][76] , \CARRYB[8][75] , \CARRYB[8][74] , \CARRYB[8][73] ,
         \CARRYB[8][72] , \CARRYB[8][71] , \CARRYB[8][70] , \CARRYB[8][69] ,
         \CARRYB[8][68] , \CARRYB[8][67] , \CARRYB[8][66] , \CARRYB[8][65] ,
         \CARRYB[8][64] , \SUMB[13][94] , \SUMB[13][93] , \SUMB[13][92] ,
         \SUMB[13][91] , \SUMB[13][90] , \SUMB[13][89] , \SUMB[13][88] ,
         \SUMB[13][87] , \SUMB[13][86] , \SUMB[13][85] , \SUMB[13][84] ,
         \SUMB[13][83] , \SUMB[13][82] , \SUMB[13][81] , \SUMB[13][80] ,
         \SUMB[13][79] , \SUMB[13][78] , \SUMB[13][77] , \SUMB[13][76] ,
         \SUMB[13][75] , \SUMB[13][74] , \SUMB[13][73] , \SUMB[13][72] ,
         \SUMB[13][71] , \SUMB[13][70] , \SUMB[13][69] , \SUMB[13][68] ,
         \SUMB[13][67] , \SUMB[13][66] , \SUMB[13][65] , \SUMB[13][64] ,
         \SUMB[13][63] , \SUMB[13][62] , \SUMB[13][61] , \SUMB[13][60] ,
         \SUMB[13][59] , \SUMB[13][58] , \SUMB[13][57] , \SUMB[13][56] ,
         \SUMB[13][55] , \SUMB[13][54] , \SUMB[13][53] , \SUMB[13][52] ,
         \SUMB[13][51] , \SUMB[13][50] , \SUMB[13][49] , \SUMB[13][48] ,
         \SUMB[13][47] , \SUMB[13][46] , \SUMB[13][45] , \SUMB[13][44] ,
         \SUMB[13][43] , \SUMB[13][42] , \SUMB[13][41] , \SUMB[13][40] ,
         \SUMB[13][39] , \SUMB[13][38] , \SUMB[13][37] , \SUMB[13][36] ,
         \SUMB[13][35] , \SUMB[13][34] , \SUMB[13][33] , \SUMB[13][32] ,
         \SUMB[13][31] , \SUMB[13][30] , \SUMB[13][29] , \SUMB[13][28] ,
         \SUMB[13][27] , \SUMB[13][26] , \SUMB[13][25] , \SUMB[13][24] ,
         \SUMB[13][23] , \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] ,
         \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] ,
         \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][94] ,
         \SUMB[12][93] , \SUMB[12][92] , \SUMB[12][91] , \SUMB[12][90] ,
         \SUMB[12][89] , \SUMB[12][88] , \SUMB[12][87] , \SUMB[12][86] ,
         \SUMB[12][85] , \SUMB[12][84] , \SUMB[12][83] , \SUMB[12][82] ,
         \SUMB[12][81] , \SUMB[12][80] , \SUMB[12][79] , \SUMB[12][78] ,
         \SUMB[12][77] , \SUMB[12][76] , \SUMB[12][75] , \SUMB[12][74] ,
         \SUMB[12][73] , \SUMB[12][72] , \SUMB[12][71] , \SUMB[12][70] ,
         \SUMB[12][69] , \SUMB[12][68] , \SUMB[12][67] , \SUMB[12][66] ,
         \SUMB[12][65] , \SUMB[12][64] , \SUMB[12][63] , \SUMB[12][62] ,
         \SUMB[12][61] , \SUMB[12][60] , \SUMB[12][59] , \SUMB[12][58] ,
         \SUMB[12][57] , \SUMB[12][56] , \SUMB[12][55] , \SUMB[12][54] ,
         \SUMB[12][53] , \SUMB[12][52] , \SUMB[12][51] , \SUMB[12][50] ,
         \SUMB[12][49] , \SUMB[12][48] , \SUMB[12][47] , \SUMB[12][46] ,
         \SUMB[12][45] , \SUMB[12][44] , \SUMB[12][43] , \SUMB[12][42] ,
         \SUMB[12][41] , \SUMB[12][40] , \SUMB[12][39] , \SUMB[12][38] ,
         \SUMB[12][37] , \SUMB[12][36] , \SUMB[12][35] , \SUMB[12][34] ,
         \SUMB[12][33] , \SUMB[12][32] , \SUMB[12][31] , \SUMB[12][30] ,
         \SUMB[12][29] , \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] ,
         \SUMB[12][25] , \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] ,
         \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] ,
         \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][94] , \SUMB[11][93] , \SUMB[11][92] ,
         \SUMB[11][91] , \SUMB[11][90] , \SUMB[11][89] , \SUMB[11][88] ,
         \SUMB[11][87] , \SUMB[11][86] , \SUMB[11][85] , \SUMB[11][84] ,
         \SUMB[11][83] , \SUMB[11][82] , \SUMB[11][81] , \SUMB[11][80] ,
         \SUMB[11][79] , \SUMB[11][78] , \SUMB[11][77] , \SUMB[11][76] ,
         \SUMB[11][75] , \SUMB[11][74] , \SUMB[11][73] , \SUMB[11][72] ,
         \SUMB[11][71] , \SUMB[11][70] , \SUMB[11][69] , \SUMB[11][68] ,
         \SUMB[11][67] , \SUMB[11][66] , \SUMB[11][65] , \SUMB[11][64] ,
         \SUMB[11][63] , \SUMB[11][62] , \SUMB[11][61] , \SUMB[11][60] ,
         \SUMB[11][59] , \SUMB[11][58] , \SUMB[11][57] , \SUMB[11][56] ,
         \SUMB[11][55] , \SUMB[11][54] , \SUMB[11][53] , \SUMB[11][52] ,
         \SUMB[11][51] , \SUMB[11][50] , \SUMB[11][49] , \SUMB[11][48] ,
         \SUMB[11][47] , \SUMB[11][46] , \SUMB[11][45] , \SUMB[11][44] ,
         \SUMB[11][43] , \SUMB[11][42] , \SUMB[11][41] , \SUMB[11][40] ,
         \SUMB[11][39] , \SUMB[11][38] , \SUMB[11][37] , \SUMB[11][36] ,
         \SUMB[11][35] , \SUMB[11][34] , \SUMB[11][33] , \SUMB[11][32] ,
         \SUMB[11][31] , \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] ,
         \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] ,
         \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][94] ,
         \SUMB[10][93] , \SUMB[10][92] , \SUMB[10][91] , \SUMB[10][90] ,
         \SUMB[10][89] , \SUMB[10][88] , \SUMB[10][87] , \SUMB[10][86] ,
         \SUMB[10][85] , \SUMB[10][84] , \SUMB[10][83] , \SUMB[10][82] ,
         \SUMB[10][81] , \SUMB[10][80] , \SUMB[10][79] , \SUMB[10][78] ,
         \SUMB[10][77] , \SUMB[10][76] , \SUMB[10][75] , \SUMB[10][74] ,
         \SUMB[10][73] , \SUMB[10][72] , \SUMB[10][71] , \SUMB[10][70] ,
         \SUMB[10][69] , \SUMB[10][68] , \SUMB[10][67] , \SUMB[10][66] ,
         \SUMB[10][65] , \SUMB[10][64] , \SUMB[10][63] , \SUMB[10][62] ,
         \SUMB[10][61] , \SUMB[10][60] , \SUMB[10][59] , \SUMB[10][58] ,
         \SUMB[10][57] , \SUMB[10][56] , \SUMB[10][55] , \SUMB[10][54] ,
         \SUMB[10][53] , \SUMB[10][52] , \SUMB[10][51] , \SUMB[10][50] ,
         \SUMB[10][49] , \SUMB[10][48] , \SUMB[10][47] , \SUMB[10][46] ,
         \SUMB[10][45] , \SUMB[10][44] , \SUMB[10][43] , \SUMB[10][42] ,
         \SUMB[10][41] , \SUMB[10][40] , \SUMB[10][39] , \SUMB[10][38] ,
         \SUMB[10][37] , \SUMB[10][36] , \SUMB[10][35] , \SUMB[10][34] ,
         \SUMB[10][33] , \SUMB[10][32] , \SUMB[10][31] , \SUMB[10][30] ,
         \SUMB[10][29] , \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] ,
         \SUMB[10][25] , \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] ,
         \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] ,
         \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][94] , \SUMB[9][93] , \SUMB[9][92] ,
         \SUMB[9][91] , \SUMB[9][90] , \SUMB[9][89] , \SUMB[9][88] ,
         \SUMB[9][87] , \SUMB[9][86] , \SUMB[9][85] , \SUMB[9][84] ,
         \SUMB[9][83] , \SUMB[9][82] , \SUMB[9][81] , \SUMB[9][80] ,
         \SUMB[9][79] , \SUMB[9][78] , \SUMB[9][77] , \SUMB[9][76] ,
         \SUMB[9][75] , \SUMB[9][74] , \SUMB[9][73] , \SUMB[9][72] ,
         \SUMB[9][71] , \SUMB[9][70] , \SUMB[9][69] , \SUMB[9][68] ,
         \SUMB[9][67] , \SUMB[9][66] , \SUMB[9][65] , \SUMB[9][64] ,
         \SUMB[9][63] , \SUMB[9][62] , \SUMB[9][61] , \SUMB[9][60] ,
         \SUMB[9][59] , \SUMB[9][58] , \SUMB[9][57] , \SUMB[9][56] ,
         \SUMB[9][55] , \SUMB[9][54] , \SUMB[9][53] , \SUMB[9][52] ,
         \SUMB[9][51] , \SUMB[9][50] , \SUMB[9][49] , \SUMB[9][48] ,
         \SUMB[9][47] , \SUMB[9][46] , \SUMB[9][45] , \SUMB[9][44] ,
         \SUMB[9][43] , \SUMB[9][42] , \SUMB[9][41] , \SUMB[9][40] ,
         \SUMB[9][39] , \SUMB[9][38] , \SUMB[9][37] , \SUMB[9][36] ,
         \SUMB[9][35] , \SUMB[9][34] , \SUMB[9][33] , \SUMB[9][32] ,
         \SUMB[9][31] , \SUMB[9][30] , \SUMB[9][29] , \SUMB[9][28] ,
         \SUMB[9][27] , \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] ,
         \SUMB[9][23] , \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] ,
         \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] ,
         \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][94] , \SUMB[8][93] ,
         \SUMB[8][92] , \SUMB[8][91] , \SUMB[8][90] , \SUMB[8][89] ,
         \SUMB[8][88] , \SUMB[8][87] , \SUMB[8][86] , \SUMB[8][85] ,
         \SUMB[8][84] , \SUMB[8][83] , \SUMB[8][82] , \SUMB[8][81] ,
         \SUMB[8][80] , \SUMB[8][79] , \SUMB[8][78] , \SUMB[8][77] ,
         \SUMB[8][76] , \SUMB[8][75] , \SUMB[8][74] , \SUMB[8][73] ,
         \SUMB[8][72] , \SUMB[8][71] , \SUMB[8][70] , \SUMB[8][69] ,
         \SUMB[8][68] , \SUMB[8][67] , \SUMB[8][66] , \SUMB[8][65] ,
         \SUMB[8][64] , \CARRYB[19][31] , \CARRYB[19][30] , \CARRYB[19][29] ,
         \CARRYB[19][28] , \CARRYB[19][27] , \CARRYB[19][26] ,
         \CARRYB[19][25] , \CARRYB[19][24] , \CARRYB[19][23] ,
         \CARRYB[19][22] , \CARRYB[19][21] , \CARRYB[19][20] ,
         \CARRYB[19][19] , \CARRYB[19][18] , \CARRYB[19][17] ,
         \CARRYB[19][16] , \CARRYB[19][15] , \CARRYB[19][14] ,
         \CARRYB[19][13] , \CARRYB[19][12] , \CARRYB[19][11] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][94] ,
         \CARRYB[18][93] , \CARRYB[18][92] , \CARRYB[18][91] ,
         \CARRYB[18][90] , \CARRYB[18][89] , \CARRYB[18][88] ,
         \CARRYB[18][87] , \CARRYB[18][86] , \CARRYB[18][85] ,
         \CARRYB[18][84] , \CARRYB[18][83] , \CARRYB[18][82] ,
         \CARRYB[18][81] , \CARRYB[18][80] , \CARRYB[18][79] ,
         \CARRYB[18][78] , \CARRYB[18][77] , \CARRYB[18][76] ,
         \CARRYB[18][75] , \CARRYB[18][74] , \CARRYB[18][73] ,
         \CARRYB[18][72] , \CARRYB[18][71] , \CARRYB[18][70] ,
         \CARRYB[18][69] , \CARRYB[18][68] , \CARRYB[18][67] ,
         \CARRYB[18][66] , \CARRYB[18][65] , \CARRYB[18][64] ,
         \CARRYB[18][63] , \CARRYB[18][62] , \CARRYB[18][61] ,
         \CARRYB[18][60] , \CARRYB[18][59] , \CARRYB[18][58] ,
         \CARRYB[18][57] , \CARRYB[18][56] , \CARRYB[18][55] ,
         \CARRYB[18][54] , \CARRYB[18][53] , \CARRYB[18][52] ,
         \CARRYB[18][51] , \CARRYB[18][50] , \CARRYB[18][49] ,
         \CARRYB[18][48] , \CARRYB[18][47] , \CARRYB[18][46] ,
         \CARRYB[18][45] , \CARRYB[18][44] , \CARRYB[18][43] ,
         \CARRYB[18][42] , \CARRYB[18][41] , \CARRYB[18][40] ,
         \CARRYB[18][39] , \CARRYB[18][38] , \CARRYB[18][37] ,
         \CARRYB[18][36] , \CARRYB[18][35] , \CARRYB[18][34] ,
         \CARRYB[18][33] , \CARRYB[18][32] , \CARRYB[18][31] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][94] , \CARRYB[17][93] , \CARRYB[17][92] ,
         \CARRYB[17][91] , \CARRYB[17][90] , \CARRYB[17][89] ,
         \CARRYB[17][88] , \CARRYB[17][87] , \CARRYB[17][86] ,
         \CARRYB[17][85] , \CARRYB[17][84] , \CARRYB[17][83] ,
         \CARRYB[17][82] , \CARRYB[17][81] , \CARRYB[17][80] ,
         \CARRYB[17][79] , \CARRYB[17][78] , \CARRYB[17][77] ,
         \CARRYB[17][76] , \CARRYB[17][75] , \CARRYB[17][74] ,
         \CARRYB[17][73] , \CARRYB[17][72] , \CARRYB[17][71] ,
         \CARRYB[17][70] , \CARRYB[17][69] , \CARRYB[17][68] ,
         \CARRYB[17][67] , \CARRYB[17][66] , \CARRYB[17][65] ,
         \CARRYB[17][64] , \CARRYB[17][63] , \CARRYB[17][62] ,
         \CARRYB[17][61] , \CARRYB[17][60] , \CARRYB[17][59] ,
         \CARRYB[17][58] , \CARRYB[17][57] , \CARRYB[17][56] ,
         \CARRYB[17][55] , \CARRYB[17][54] , \CARRYB[17][53] ,
         \CARRYB[17][52] , \CARRYB[17][51] , \CARRYB[17][50] ,
         \CARRYB[17][49] , \CARRYB[17][48] , \CARRYB[17][47] ,
         \CARRYB[17][46] , \CARRYB[17][45] , \CARRYB[17][44] ,
         \CARRYB[17][43] , \CARRYB[17][42] , \CARRYB[17][41] ,
         \CARRYB[17][40] , \CARRYB[17][39] , \CARRYB[17][38] ,
         \CARRYB[17][37] , \CARRYB[17][36] , \CARRYB[17][35] ,
         \CARRYB[17][34] , \CARRYB[17][33] , \CARRYB[17][32] ,
         \CARRYB[17][31] , \CARRYB[17][30] , \CARRYB[17][29] ,
         \CARRYB[17][28] , \CARRYB[17][27] , \CARRYB[17][26] ,
         \CARRYB[17][25] , \CARRYB[17][24] , \CARRYB[17][23] ,
         \CARRYB[17][22] , \CARRYB[17][21] , \CARRYB[17][20] ,
         \CARRYB[17][19] , \CARRYB[17][18] , \CARRYB[17][17] ,
         \CARRYB[17][16] , \CARRYB[17][15] , \CARRYB[17][14] ,
         \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][94] ,
         \CARRYB[16][93] , \CARRYB[16][92] , \CARRYB[16][91] ,
         \CARRYB[16][90] , \CARRYB[16][89] , \CARRYB[16][88] ,
         \CARRYB[16][87] , \CARRYB[16][86] , \CARRYB[16][85] ,
         \CARRYB[16][84] , \CARRYB[16][83] , \CARRYB[16][82] ,
         \CARRYB[16][81] , \CARRYB[16][80] , \CARRYB[16][79] ,
         \CARRYB[16][78] , \CARRYB[16][77] , \CARRYB[16][76] ,
         \CARRYB[16][75] , \CARRYB[16][74] , \CARRYB[16][73] ,
         \CARRYB[16][72] , \CARRYB[16][71] , \CARRYB[16][70] ,
         \CARRYB[16][69] , \CARRYB[16][68] , \CARRYB[16][67] ,
         \CARRYB[16][66] , \CARRYB[16][65] , \CARRYB[16][64] ,
         \CARRYB[16][63] , \CARRYB[16][62] , \CARRYB[16][61] ,
         \CARRYB[16][60] , \CARRYB[16][59] , \CARRYB[16][58] ,
         \CARRYB[16][57] , \CARRYB[16][56] , \CARRYB[16][55] ,
         \CARRYB[16][54] , \CARRYB[16][53] , \CARRYB[16][52] ,
         \CARRYB[16][51] , \CARRYB[16][50] , \CARRYB[16][49] ,
         \CARRYB[16][48] , \CARRYB[16][47] , \CARRYB[16][46] ,
         \CARRYB[16][45] , \CARRYB[16][44] , \CARRYB[16][43] ,
         \CARRYB[16][42] , \CARRYB[16][41] , \CARRYB[16][40] ,
         \CARRYB[16][39] , \CARRYB[16][38] , \CARRYB[16][37] ,
         \CARRYB[16][36] , \CARRYB[16][35] , \CARRYB[16][34] ,
         \CARRYB[16][33] , \CARRYB[16][32] , \CARRYB[16][31] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \CARRYB[15][94] , \CARRYB[15][93] , \CARRYB[15][92] ,
         \CARRYB[15][91] , \CARRYB[15][90] , \CARRYB[15][89] ,
         \CARRYB[15][88] , \CARRYB[15][87] , \CARRYB[15][86] ,
         \CARRYB[15][85] , \CARRYB[15][84] , \CARRYB[15][83] ,
         \CARRYB[15][82] , \CARRYB[15][81] , \CARRYB[15][80] ,
         \CARRYB[15][79] , \CARRYB[15][78] , \CARRYB[15][77] ,
         \CARRYB[15][76] , \CARRYB[15][75] , \CARRYB[15][74] ,
         \CARRYB[15][73] , \CARRYB[15][72] , \CARRYB[15][71] ,
         \CARRYB[15][70] , \CARRYB[15][69] , \CARRYB[15][68] ,
         \CARRYB[15][67] , \CARRYB[15][66] , \CARRYB[15][65] ,
         \CARRYB[15][64] , \CARRYB[15][63] , \CARRYB[15][62] ,
         \CARRYB[15][61] , \CARRYB[15][60] , \CARRYB[15][59] ,
         \CARRYB[15][58] , \CARRYB[15][57] , \CARRYB[15][56] ,
         \CARRYB[15][55] , \CARRYB[15][54] , \CARRYB[15][53] ,
         \CARRYB[15][52] , \CARRYB[15][51] , \CARRYB[15][50] ,
         \CARRYB[15][49] , \CARRYB[15][48] , \CARRYB[15][47] ,
         \CARRYB[15][46] , \CARRYB[15][45] , \CARRYB[15][44] ,
         \CARRYB[15][43] , \CARRYB[15][42] , \CARRYB[15][41] ,
         \CARRYB[15][40] , \CARRYB[15][39] , \CARRYB[15][38] ,
         \CARRYB[15][37] , \CARRYB[15][36] , \CARRYB[15][35] ,
         \CARRYB[15][34] , \CARRYB[15][33] , \CARRYB[15][32] ,
         \CARRYB[15][31] , \CARRYB[15][30] , \CARRYB[15][29] ,
         \CARRYB[15][28] , \CARRYB[15][27] , \CARRYB[15][26] ,
         \CARRYB[15][25] , \CARRYB[15][24] , \CARRYB[15][23] ,
         \CARRYB[15][22] , \CARRYB[15][21] , \CARRYB[15][20] ,
         \CARRYB[15][19] , \CARRYB[15][18] , \CARRYB[15][17] ,
         \CARRYB[15][16] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][94] ,
         \CARRYB[14][93] , \CARRYB[14][92] , \CARRYB[14][91] ,
         \CARRYB[14][90] , \CARRYB[14][89] , \CARRYB[14][88] ,
         \CARRYB[14][87] , \CARRYB[14][86] , \CARRYB[14][85] ,
         \CARRYB[14][84] , \CARRYB[14][83] , \CARRYB[14][82] ,
         \CARRYB[14][81] , \CARRYB[14][80] , \CARRYB[14][79] ,
         \CARRYB[14][78] , \CARRYB[14][77] , \CARRYB[14][76] ,
         \CARRYB[14][75] , \CARRYB[14][74] , \CARRYB[14][73] ,
         \CARRYB[14][72] , \CARRYB[14][71] , \CARRYB[14][70] ,
         \CARRYB[14][69] , \CARRYB[14][68] , \CARRYB[14][67] ,
         \CARRYB[14][66] , \CARRYB[14][65] , \CARRYB[14][64] ,
         \CARRYB[14][63] , \CARRYB[14][62] , \CARRYB[14][61] ,
         \CARRYB[14][60] , \CARRYB[14][59] , \CARRYB[14][58] ,
         \CARRYB[14][57] , \CARRYB[14][56] , \CARRYB[14][55] ,
         \CARRYB[14][54] , \CARRYB[14][53] , \CARRYB[14][52] ,
         \CARRYB[14][51] , \CARRYB[14][50] , \CARRYB[14][49] ,
         \CARRYB[14][48] , \CARRYB[14][47] , \CARRYB[14][46] ,
         \CARRYB[14][45] , \CARRYB[14][44] , \CARRYB[14][43] ,
         \CARRYB[14][42] , \CARRYB[14][41] , \CARRYB[14][40] ,
         \CARRYB[14][39] , \CARRYB[14][38] , \CARRYB[14][37] ,
         \CARRYB[14][36] , \CARRYB[14][35] , \CARRYB[14][34] ,
         \CARRYB[14][33] , \CARRYB[14][32] , \CARRYB[14][31] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \SUMB[19][31] , \SUMB[19][30] , \SUMB[19][29] ,
         \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] , \SUMB[19][25] ,
         \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] , \SUMB[19][21] ,
         \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] ,
         \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] ,
         \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] ,
         \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] ,
         \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] ,
         \SUMB[18][94] , \SUMB[18][93] , \SUMB[18][92] , \SUMB[18][91] ,
         \SUMB[18][90] , \SUMB[18][89] , \SUMB[18][88] , \SUMB[18][87] ,
         \SUMB[18][86] , \SUMB[18][85] , \SUMB[18][84] , \SUMB[18][83] ,
         \SUMB[18][82] , \SUMB[18][81] , \SUMB[18][80] , \SUMB[18][79] ,
         \SUMB[18][78] , \SUMB[18][77] , \SUMB[18][76] , \SUMB[18][75] ,
         \SUMB[18][74] , \SUMB[18][73] , \SUMB[18][72] , \SUMB[18][71] ,
         \SUMB[18][70] , \SUMB[18][69] , \SUMB[18][68] , \SUMB[18][67] ,
         \SUMB[18][66] , \SUMB[18][65] , \SUMB[18][64] , \SUMB[18][63] ,
         \SUMB[18][62] , \SUMB[18][61] , \SUMB[18][60] , \SUMB[18][59] ,
         \SUMB[18][58] , \SUMB[18][57] , \SUMB[18][56] , \SUMB[18][55] ,
         \SUMB[18][54] , \SUMB[18][53] , \SUMB[18][52] , \SUMB[18][51] ,
         \SUMB[18][50] , \SUMB[18][49] , \SUMB[18][48] , \SUMB[18][47] ,
         \SUMB[18][46] , \SUMB[18][45] , \SUMB[18][44] , \SUMB[18][43] ,
         \SUMB[18][42] , \SUMB[18][41] , \SUMB[18][40] , \SUMB[18][39] ,
         \SUMB[18][38] , \SUMB[18][37] , \SUMB[18][36] , \SUMB[18][35] ,
         \SUMB[18][34] , \SUMB[18][33] , \SUMB[18][32] , \SUMB[18][31] ,
         \SUMB[18][30] , \SUMB[18][29] , \SUMB[18][28] , \SUMB[18][27] ,
         \SUMB[18][26] , \SUMB[18][25] , \SUMB[18][24] , \SUMB[18][23] ,
         \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] ,
         \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] ,
         \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] ,
         \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] ,
         \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][94] , \SUMB[17][93] ,
         \SUMB[17][92] , \SUMB[17][91] , \SUMB[17][90] , \SUMB[17][89] ,
         \SUMB[17][88] , \SUMB[17][87] , \SUMB[17][86] , \SUMB[17][85] ,
         \SUMB[17][84] , \SUMB[17][83] , \SUMB[17][82] , \SUMB[17][81] ,
         \SUMB[17][80] , \SUMB[17][79] , \SUMB[17][78] , \SUMB[17][77] ,
         \SUMB[17][76] , \SUMB[17][75] , \SUMB[17][74] , \SUMB[17][73] ,
         \SUMB[17][72] , \SUMB[17][71] , \SUMB[17][70] , \SUMB[17][69] ,
         \SUMB[17][68] , \SUMB[17][67] , \SUMB[17][66] , \SUMB[17][65] ,
         \SUMB[17][64] , \SUMB[17][63] , \SUMB[17][62] , \SUMB[17][61] ,
         \SUMB[17][60] , \SUMB[17][59] , \SUMB[17][58] , \SUMB[17][57] ,
         \SUMB[17][56] , \SUMB[17][55] , \SUMB[17][54] , \SUMB[17][53] ,
         \SUMB[17][52] , \SUMB[17][51] , \SUMB[17][50] , \SUMB[17][49] ,
         \SUMB[17][48] , \SUMB[17][47] , \SUMB[17][46] , \SUMB[17][45] ,
         \SUMB[17][44] , \SUMB[17][43] , \SUMB[17][42] , \SUMB[17][41] ,
         \SUMB[17][40] , \SUMB[17][39] , \SUMB[17][38] , \SUMB[17][37] ,
         \SUMB[17][36] , \SUMB[17][35] , \SUMB[17][34] , \SUMB[17][33] ,
         \SUMB[17][32] , \SUMB[17][31] , \SUMB[17][30] , \SUMB[17][29] ,
         \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] , \SUMB[17][25] ,
         \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] , \SUMB[17][21] ,
         \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] ,
         \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][94] , \SUMB[16][93] , \SUMB[16][92] , \SUMB[16][91] ,
         \SUMB[16][90] , \SUMB[16][89] , \SUMB[16][88] , \SUMB[16][87] ,
         \SUMB[16][86] , \SUMB[16][85] , \SUMB[16][84] , \SUMB[16][83] ,
         \SUMB[16][82] , \SUMB[16][81] , \SUMB[16][80] , \SUMB[16][79] ,
         \SUMB[16][78] , \SUMB[16][77] , \SUMB[16][76] , \SUMB[16][75] ,
         \SUMB[16][74] , \SUMB[16][73] , \SUMB[16][72] , \SUMB[16][71] ,
         \SUMB[16][70] , \SUMB[16][69] , \SUMB[16][68] , \SUMB[16][67] ,
         \SUMB[16][66] , \SUMB[16][65] , \SUMB[16][64] , \SUMB[16][63] ,
         \SUMB[16][62] , \SUMB[16][61] , \SUMB[16][60] , \SUMB[16][59] ,
         \SUMB[16][58] , \SUMB[16][57] , \SUMB[16][56] , \SUMB[16][55] ,
         \SUMB[16][54] , \SUMB[16][53] , \SUMB[16][52] , \SUMB[16][51] ,
         \SUMB[16][50] , \SUMB[16][49] , \SUMB[16][48] , \SUMB[16][47] ,
         \SUMB[16][46] , \SUMB[16][45] , \SUMB[16][44] , \SUMB[16][43] ,
         \SUMB[16][42] , \SUMB[16][41] , \SUMB[16][40] , \SUMB[16][39] ,
         \SUMB[16][38] , \SUMB[16][37] , \SUMB[16][36] , \SUMB[16][35] ,
         \SUMB[16][34] , \SUMB[16][33] , \SUMB[16][32] , \SUMB[16][31] ,
         \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] , \SUMB[16][27] ,
         \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] , \SUMB[16][23] ,
         \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][19] ,
         \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] , \SUMB[16][15] ,
         \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] ,
         \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] ,
         \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] ,
         \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][94] , \SUMB[15][93] ,
         \SUMB[15][92] , \SUMB[15][91] , \SUMB[15][90] , \SUMB[15][89] ,
         \SUMB[15][88] , \SUMB[15][87] , \SUMB[15][86] , \SUMB[15][85] ,
         \SUMB[15][84] , \SUMB[15][83] , \SUMB[15][82] , \SUMB[15][81] ,
         \SUMB[15][80] , \SUMB[15][79] , \SUMB[15][78] , \SUMB[15][77] ,
         \SUMB[15][76] , \SUMB[15][75] , \SUMB[15][74] , \SUMB[15][73] ,
         \SUMB[15][72] , \SUMB[15][71] , \SUMB[15][70] , \SUMB[15][69] ,
         \SUMB[15][68] , \SUMB[15][67] , \SUMB[15][66] , \SUMB[15][65] ,
         \SUMB[15][64] , \SUMB[15][63] , \SUMB[15][62] , \SUMB[15][61] ,
         \SUMB[15][60] , \SUMB[15][59] , \SUMB[15][58] , \SUMB[15][57] ,
         \SUMB[15][56] , \SUMB[15][55] , \SUMB[15][54] , \SUMB[15][53] ,
         \SUMB[15][52] , \SUMB[15][51] , \SUMB[15][50] , \SUMB[15][49] ,
         \SUMB[15][48] , \SUMB[15][47] , \SUMB[15][46] , \SUMB[15][45] ,
         \SUMB[15][44] , \SUMB[15][43] , \SUMB[15][42] , \SUMB[15][41] ,
         \SUMB[15][40] , \SUMB[15][39] , \SUMB[15][38] , \SUMB[15][37] ,
         \SUMB[15][36] , \SUMB[15][35] , \SUMB[15][34] , \SUMB[15][33] ,
         \SUMB[15][32] , \SUMB[15][31] , \SUMB[15][30] , \SUMB[15][29] ,
         \SUMB[15][28] , \SUMB[15][27] , \SUMB[15][26] , \SUMB[15][25] ,
         \SUMB[15][24] , \SUMB[15][23] , \SUMB[15][22] , \SUMB[15][21] ,
         \SUMB[15][20] , \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] ,
         \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][94] , \SUMB[14][93] , \SUMB[14][92] , \SUMB[14][91] ,
         \SUMB[14][90] , \SUMB[14][89] , \SUMB[14][88] , \SUMB[14][87] ,
         \SUMB[14][86] , \SUMB[14][85] , \SUMB[14][84] , \SUMB[14][83] ,
         \SUMB[14][82] , \SUMB[14][81] , \SUMB[14][80] , \SUMB[14][79] ,
         \SUMB[14][78] , \SUMB[14][77] , \SUMB[14][76] , \SUMB[14][75] ,
         \SUMB[14][74] , \SUMB[14][73] , \SUMB[14][72] , \SUMB[14][71] ,
         \SUMB[14][70] , \SUMB[14][69] , \SUMB[14][68] , \SUMB[14][67] ,
         \SUMB[14][66] , \SUMB[14][65] , \SUMB[14][64] , \SUMB[14][63] ,
         \SUMB[14][62] , \SUMB[14][61] , \SUMB[14][60] , \SUMB[14][59] ,
         \SUMB[14][58] , \SUMB[14][57] , \SUMB[14][56] , \SUMB[14][55] ,
         \SUMB[14][54] , \SUMB[14][53] , \SUMB[14][52] , \SUMB[14][51] ,
         \SUMB[14][50] , \SUMB[14][49] , \SUMB[14][48] , \SUMB[14][47] ,
         \SUMB[14][46] , \SUMB[14][45] , \SUMB[14][44] , \SUMB[14][43] ,
         \SUMB[14][42] , \SUMB[14][41] , \SUMB[14][40] , \SUMB[14][39] ,
         \SUMB[14][38] , \SUMB[14][37] , \SUMB[14][36] , \SUMB[14][35] ,
         \SUMB[14][34] , \SUMB[14][33] , \SUMB[14][32] , \SUMB[14][31] ,
         \SUMB[14][30] , \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] ,
         \SUMB[14][26] , \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] ,
         \SUMB[14][22] , \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] ,
         \SUMB[14][18] , \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] ,
         \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] ,
         \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] ,
         \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] ,
         \SUMB[14][2] , \SUMB[14][1] , \CARRYB[24][63] , \CARRYB[24][62] ,
         \CARRYB[24][61] , \CARRYB[24][60] , \CARRYB[24][59] ,
         \CARRYB[24][58] , \CARRYB[24][57] , \CARRYB[24][56] ,
         \CARRYB[24][55] , \CARRYB[24][54] , \CARRYB[24][53] ,
         \CARRYB[24][52] , \CARRYB[24][51] , \CARRYB[24][50] ,
         \CARRYB[24][49] , \CARRYB[24][48] , \CARRYB[24][47] ,
         \CARRYB[24][46] , \CARRYB[24][45] , \CARRYB[24][44] ,
         \CARRYB[24][43] , \CARRYB[24][42] , \CARRYB[24][41] ,
         \CARRYB[24][40] , \CARRYB[24][39] , \CARRYB[24][38] ,
         \CARRYB[24][37] , \CARRYB[24][36] , \CARRYB[24][35] ,
         \CARRYB[24][34] , \CARRYB[24][33] , \CARRYB[24][32] ,
         \CARRYB[24][31] , \CARRYB[24][30] , \CARRYB[24][29] ,
         \CARRYB[24][28] , \CARRYB[24][27] , \CARRYB[24][26] ,
         \CARRYB[24][25] , \CARRYB[24][24] , \CARRYB[24][23] ,
         \CARRYB[24][22] , \CARRYB[24][21] , \CARRYB[24][20] ,
         \CARRYB[24][19] , \CARRYB[24][18] , \CARRYB[24][17] ,
         \CARRYB[24][16] , \CARRYB[24][15] , \CARRYB[24][14] ,
         \CARRYB[24][13] , \CARRYB[24][12] , \CARRYB[24][11] ,
         \CARRYB[24][10] , \CARRYB[24][9] , \CARRYB[24][8] , \CARRYB[24][7] ,
         \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][3] ,
         \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] , \CARRYB[23][94] ,
         \CARRYB[23][93] , \CARRYB[23][92] , \CARRYB[23][91] ,
         \CARRYB[23][90] , \CARRYB[23][89] , \CARRYB[23][88] ,
         \CARRYB[23][87] , \CARRYB[23][86] , \CARRYB[23][85] ,
         \CARRYB[23][84] , \CARRYB[23][83] , \CARRYB[23][82] ,
         \CARRYB[23][81] , \CARRYB[23][80] , \CARRYB[23][79] ,
         \CARRYB[23][78] , \CARRYB[23][77] , \CARRYB[23][76] ,
         \CARRYB[23][75] , \CARRYB[23][74] , \CARRYB[23][73] ,
         \CARRYB[23][72] , \CARRYB[23][71] , \CARRYB[23][70] ,
         \CARRYB[23][69] , \CARRYB[23][68] , \CARRYB[23][67] ,
         \CARRYB[23][66] , \CARRYB[23][65] , \CARRYB[23][64] ,
         \CARRYB[23][63] , \CARRYB[23][62] , \CARRYB[23][61] ,
         \CARRYB[23][60] , \CARRYB[23][59] , \CARRYB[23][58] ,
         \CARRYB[23][57] , \CARRYB[23][56] , \CARRYB[23][55] ,
         \CARRYB[23][54] , \CARRYB[23][53] , \CARRYB[23][52] ,
         \CARRYB[23][51] , \CARRYB[23][50] , \CARRYB[23][49] ,
         \CARRYB[23][48] , \CARRYB[23][47] , \CARRYB[23][46] ,
         \CARRYB[23][45] , \CARRYB[23][44] , \CARRYB[23][43] ,
         \CARRYB[23][42] , \CARRYB[23][41] , \CARRYB[23][40] ,
         \CARRYB[23][39] , \CARRYB[23][38] , \CARRYB[23][37] ,
         \CARRYB[23][36] , \CARRYB[23][35] , \CARRYB[23][34] ,
         \CARRYB[23][33] , \CARRYB[23][32] , \CARRYB[23][31] ,
         \CARRYB[23][30] , \CARRYB[23][29] , \CARRYB[23][28] ,
         \CARRYB[23][27] , \CARRYB[23][26] , \CARRYB[23][25] ,
         \CARRYB[23][24] , \CARRYB[23][23] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][94] , \CARRYB[22][93] , \CARRYB[22][92] ,
         \CARRYB[22][91] , \CARRYB[22][90] , \CARRYB[22][89] ,
         \CARRYB[22][88] , \CARRYB[22][87] , \CARRYB[22][86] ,
         \CARRYB[22][85] , \CARRYB[22][84] , \CARRYB[22][83] ,
         \CARRYB[22][82] , \CARRYB[22][81] , \CARRYB[22][80] ,
         \CARRYB[22][79] , \CARRYB[22][78] , \CARRYB[22][77] ,
         \CARRYB[22][76] , \CARRYB[22][75] , \CARRYB[22][74] ,
         \CARRYB[22][73] , \CARRYB[22][72] , \CARRYB[22][71] ,
         \CARRYB[22][70] , \CARRYB[22][69] , \CARRYB[22][68] ,
         \CARRYB[22][67] , \CARRYB[22][66] , \CARRYB[22][65] ,
         \CARRYB[22][64] , \CARRYB[22][63] , \CARRYB[22][62] ,
         \CARRYB[22][61] , \CARRYB[22][60] , \CARRYB[22][59] ,
         \CARRYB[22][58] , \CARRYB[22][57] , \CARRYB[22][56] ,
         \CARRYB[22][55] , \CARRYB[22][54] , \CARRYB[22][53] ,
         \CARRYB[22][52] , \CARRYB[22][51] , \CARRYB[22][50] ,
         \CARRYB[22][49] , \CARRYB[22][48] , \CARRYB[22][47] ,
         \CARRYB[22][46] , \CARRYB[22][45] , \CARRYB[22][44] ,
         \CARRYB[22][43] , \CARRYB[22][42] , \CARRYB[22][41] ,
         \CARRYB[22][40] , \CARRYB[22][39] , \CARRYB[22][38] ,
         \CARRYB[22][37] , \CARRYB[22][36] , \CARRYB[22][35] ,
         \CARRYB[22][34] , \CARRYB[22][33] , \CARRYB[22][32] ,
         \CARRYB[22][31] , \CARRYB[22][30] , \CARRYB[22][29] ,
         \CARRYB[22][28] , \CARRYB[22][27] , \CARRYB[22][26] ,
         \CARRYB[22][25] , \CARRYB[22][24] , \CARRYB[22][23] ,
         \CARRYB[22][22] , \CARRYB[22][21] , \CARRYB[22][20] ,
         \CARRYB[22][19] , \CARRYB[22][18] , \CARRYB[22][17] ,
         \CARRYB[22][16] , \CARRYB[22][15] , \CARRYB[22][14] ,
         \CARRYB[22][13] , \CARRYB[22][12] , \CARRYB[22][11] ,
         \CARRYB[22][10] , \CARRYB[22][9] , \CARRYB[22][8] , \CARRYB[22][7] ,
         \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][94] ,
         \CARRYB[21][93] , \CARRYB[21][92] , \CARRYB[21][91] ,
         \CARRYB[21][90] , \CARRYB[21][89] , \CARRYB[21][88] ,
         \CARRYB[21][87] , \CARRYB[21][86] , \CARRYB[21][85] ,
         \CARRYB[21][84] , \CARRYB[21][83] , \CARRYB[21][82] ,
         \CARRYB[21][81] , \CARRYB[21][80] , \CARRYB[21][79] ,
         \CARRYB[21][78] , \CARRYB[21][77] , \CARRYB[21][76] ,
         \CARRYB[21][75] , \CARRYB[21][74] , \CARRYB[21][73] ,
         \CARRYB[21][72] , \CARRYB[21][71] , \CARRYB[21][70] ,
         \CARRYB[21][69] , \CARRYB[21][68] , \CARRYB[21][67] ,
         \CARRYB[21][66] , \CARRYB[21][65] , \CARRYB[21][64] ,
         \CARRYB[21][63] , \CARRYB[21][62] , \CARRYB[21][61] ,
         \CARRYB[21][60] , \CARRYB[21][59] , \CARRYB[21][58] ,
         \CARRYB[21][57] , \CARRYB[21][56] , \CARRYB[21][55] ,
         \CARRYB[21][54] , \CARRYB[21][53] , \CARRYB[21][52] ,
         \CARRYB[21][51] , \CARRYB[21][50] , \CARRYB[21][49] ,
         \CARRYB[21][48] , \CARRYB[21][47] , \CARRYB[21][46] ,
         \CARRYB[21][45] , \CARRYB[21][44] , \CARRYB[21][43] ,
         \CARRYB[21][42] , \CARRYB[21][41] , \CARRYB[21][40] ,
         \CARRYB[21][39] , \CARRYB[21][38] , \CARRYB[21][37] ,
         \CARRYB[21][36] , \CARRYB[21][35] , \CARRYB[21][34] ,
         \CARRYB[21][33] , \CARRYB[21][32] , \CARRYB[21][31] ,
         \CARRYB[21][30] , \CARRYB[21][29] , \CARRYB[21][28] ,
         \CARRYB[21][27] , \CARRYB[21][26] , \CARRYB[21][25] ,
         \CARRYB[21][24] , \CARRYB[21][23] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][94] , \CARRYB[20][93] , \CARRYB[20][92] ,
         \CARRYB[20][91] , \CARRYB[20][90] , \CARRYB[20][89] ,
         \CARRYB[20][88] , \CARRYB[20][87] , \CARRYB[20][86] ,
         \CARRYB[20][85] , \CARRYB[20][84] , \CARRYB[20][83] ,
         \CARRYB[20][82] , \CARRYB[20][81] , \CARRYB[20][80] ,
         \CARRYB[20][79] , \CARRYB[20][78] , \CARRYB[20][77] ,
         \CARRYB[20][76] , \CARRYB[20][75] , \CARRYB[20][74] ,
         \CARRYB[20][73] , \CARRYB[20][72] , \CARRYB[20][71] ,
         \CARRYB[20][70] , \CARRYB[20][69] , \CARRYB[20][68] ,
         \CARRYB[20][67] , \CARRYB[20][66] , \CARRYB[20][65] ,
         \CARRYB[20][64] , \CARRYB[20][63] , \CARRYB[20][62] ,
         \CARRYB[20][61] , \CARRYB[20][60] , \CARRYB[20][59] ,
         \CARRYB[20][58] , \CARRYB[20][57] , \CARRYB[20][56] ,
         \CARRYB[20][55] , \CARRYB[20][54] , \CARRYB[20][53] ,
         \CARRYB[20][52] , \CARRYB[20][51] , \CARRYB[20][50] ,
         \CARRYB[20][49] , \CARRYB[20][48] , \CARRYB[20][47] ,
         \CARRYB[20][46] , \CARRYB[20][45] , \CARRYB[20][44] ,
         \CARRYB[20][43] , \CARRYB[20][42] , \CARRYB[20][41] ,
         \CARRYB[20][40] , \CARRYB[20][39] , \CARRYB[20][38] ,
         \CARRYB[20][37] , \CARRYB[20][36] , \CARRYB[20][35] ,
         \CARRYB[20][34] , \CARRYB[20][33] , \CARRYB[20][32] ,
         \CARRYB[20][31] , \CARRYB[20][30] , \CARRYB[20][29] ,
         \CARRYB[20][28] , \CARRYB[20][27] , \CARRYB[20][26] ,
         \CARRYB[20][25] , \CARRYB[20][24] , \CARRYB[20][23] ,
         \CARRYB[20][22] , \CARRYB[20][21] , \CARRYB[20][20] ,
         \CARRYB[20][19] , \CARRYB[20][18] , \CARRYB[20][17] ,
         \CARRYB[20][16] , \CARRYB[20][15] , \CARRYB[20][14] ,
         \CARRYB[20][13] , \CARRYB[20][12] , \CARRYB[20][11] ,
         \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] , \CARRYB[20][7] ,
         \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] , \CARRYB[20][3] ,
         \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] , \CARRYB[19][94] ,
         \CARRYB[19][93] , \CARRYB[19][92] , \CARRYB[19][91] ,
         \CARRYB[19][90] , \CARRYB[19][89] , \CARRYB[19][88] ,
         \CARRYB[19][87] , \CARRYB[19][86] , \CARRYB[19][85] ,
         \CARRYB[19][84] , \CARRYB[19][83] , \CARRYB[19][82] ,
         \CARRYB[19][81] , \CARRYB[19][80] , \CARRYB[19][79] ,
         \CARRYB[19][78] , \CARRYB[19][77] , \CARRYB[19][76] ,
         \CARRYB[19][75] , \CARRYB[19][74] , \CARRYB[19][73] ,
         \CARRYB[19][72] , \CARRYB[19][71] , \CARRYB[19][70] ,
         \CARRYB[19][69] , \CARRYB[19][68] , \CARRYB[19][67] ,
         \CARRYB[19][66] , \CARRYB[19][65] , \CARRYB[19][64] ,
         \CARRYB[19][63] , \CARRYB[19][62] , \CARRYB[19][61] ,
         \CARRYB[19][60] , \CARRYB[19][59] , \CARRYB[19][58] ,
         \CARRYB[19][57] , \CARRYB[19][56] , \CARRYB[19][55] ,
         \CARRYB[19][54] , \CARRYB[19][53] , \CARRYB[19][52] ,
         \CARRYB[19][51] , \CARRYB[19][50] , \CARRYB[19][49] ,
         \CARRYB[19][48] , \CARRYB[19][47] , \CARRYB[19][46] ,
         \CARRYB[19][45] , \CARRYB[19][44] , \CARRYB[19][43] ,
         \CARRYB[19][42] , \CARRYB[19][41] , \CARRYB[19][40] ,
         \CARRYB[19][39] , \CARRYB[19][38] , \CARRYB[19][37] ,
         \CARRYB[19][36] , \CARRYB[19][35] , \CARRYB[19][34] ,
         \CARRYB[19][33] , \CARRYB[19][32] , \SUMB[24][63] , \SUMB[24][62] ,
         \SUMB[24][61] , \SUMB[24][60] , \SUMB[24][59] , \SUMB[24][58] ,
         \SUMB[24][57] , \SUMB[24][56] , \SUMB[24][55] , \SUMB[24][54] ,
         \SUMB[24][53] , \SUMB[24][52] , \SUMB[24][51] , \SUMB[24][50] ,
         \SUMB[24][49] , \SUMB[24][48] , \SUMB[24][47] , \SUMB[24][46] ,
         \SUMB[24][45] , \SUMB[24][44] , \SUMB[24][43] , \SUMB[24][42] ,
         \SUMB[24][41] , \SUMB[24][40] , \SUMB[24][39] , \SUMB[24][38] ,
         \SUMB[24][37] , \SUMB[24][36] , \SUMB[24][35] , \SUMB[24][34] ,
         \SUMB[24][33] , \SUMB[24][32] , \SUMB[24][31] , \SUMB[24][30] ,
         \SUMB[24][29] , \SUMB[24][28] , \SUMB[24][27] , \SUMB[24][26] ,
         \SUMB[24][25] , \SUMB[24][24] , \SUMB[24][23] , \SUMB[24][22] ,
         \SUMB[24][21] , \SUMB[24][20] , \SUMB[24][19] , \SUMB[24][18] ,
         \SUMB[24][17] , \SUMB[24][16] , \SUMB[24][15] , \SUMB[24][14] ,
         \SUMB[24][13] , \SUMB[24][12] , \SUMB[24][11] , \SUMB[24][10] ,
         \SUMB[24][9] , \SUMB[24][8] , \SUMB[24][7] , \SUMB[24][6] ,
         \SUMB[24][5] , \SUMB[24][4] , \SUMB[24][3] , \SUMB[24][2] ,
         \SUMB[24][1] , \SUMB[23][94] , \SUMB[23][93] , \SUMB[23][92] ,
         \SUMB[23][91] , \SUMB[23][90] , \SUMB[23][89] , \SUMB[23][88] ,
         \SUMB[23][87] , \SUMB[23][86] , \SUMB[23][85] , \SUMB[23][84] ,
         \SUMB[23][83] , \SUMB[23][82] , \SUMB[23][81] , \SUMB[23][80] ,
         \SUMB[23][79] , \SUMB[23][78] , \SUMB[23][77] , \SUMB[23][76] ,
         \SUMB[23][75] , \SUMB[23][74] , \SUMB[23][73] , \SUMB[23][72] ,
         \SUMB[23][71] , \SUMB[23][70] , \SUMB[23][69] , \SUMB[23][68] ,
         \SUMB[23][67] , \SUMB[23][66] , \SUMB[23][65] , \SUMB[23][64] ,
         \SUMB[23][63] , \SUMB[23][62] , \SUMB[23][61] , \SUMB[23][60] ,
         \SUMB[23][59] , \SUMB[23][58] , \SUMB[23][57] , \SUMB[23][56] ,
         \SUMB[23][55] , \SUMB[23][54] , \SUMB[23][53] , \SUMB[23][52] ,
         \SUMB[23][51] , \SUMB[23][50] , \SUMB[23][49] , \SUMB[23][48] ,
         \SUMB[23][47] , \SUMB[23][46] , \SUMB[23][45] , \SUMB[23][44] ,
         \SUMB[23][43] , \SUMB[23][42] , \SUMB[23][41] , \SUMB[23][40] ,
         \SUMB[23][39] , \SUMB[23][38] , \SUMB[23][37] , \SUMB[23][36] ,
         \SUMB[23][35] , \SUMB[23][34] , \SUMB[23][33] , \SUMB[23][32] ,
         \SUMB[23][31] , \SUMB[23][30] , \SUMB[23][29] , \SUMB[23][28] ,
         \SUMB[23][27] , \SUMB[23][26] , \SUMB[23][25] , \SUMB[23][24] ,
         \SUMB[23][23] , \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] ,
         \SUMB[23][19] , \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] ,
         \SUMB[23][15] , \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] ,
         \SUMB[23][11] , \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] ,
         \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] ,
         \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][94] ,
         \SUMB[22][93] , \SUMB[22][92] , \SUMB[22][91] , \SUMB[22][90] ,
         \SUMB[22][89] , \SUMB[22][88] , \SUMB[22][87] , \SUMB[22][86] ,
         \SUMB[22][85] , \SUMB[22][84] , \SUMB[22][83] , \SUMB[22][82] ,
         \SUMB[22][81] , \SUMB[22][80] , \SUMB[22][79] , \SUMB[22][78] ,
         \SUMB[22][77] , \SUMB[22][76] , \SUMB[22][75] , \SUMB[22][74] ,
         \SUMB[22][73] , \SUMB[22][72] , \SUMB[22][71] , \SUMB[22][70] ,
         \SUMB[22][69] , \SUMB[22][68] , \SUMB[22][67] , \SUMB[22][66] ,
         \SUMB[22][65] , \SUMB[22][64] , \SUMB[22][63] , \SUMB[22][62] ,
         \SUMB[22][61] , \SUMB[22][60] , \SUMB[22][59] , \SUMB[22][58] ,
         \SUMB[22][57] , \SUMB[22][56] , \SUMB[22][55] , \SUMB[22][54] ,
         \SUMB[22][53] , \SUMB[22][52] , \SUMB[22][51] , \SUMB[22][50] ,
         \SUMB[22][49] , \SUMB[22][48] , \SUMB[22][47] , \SUMB[22][46] ,
         \SUMB[22][45] , \SUMB[22][44] , \SUMB[22][43] , \SUMB[22][42] ,
         \SUMB[22][41] , \SUMB[22][40] , \SUMB[22][39] , \SUMB[22][38] ,
         \SUMB[22][37] , \SUMB[22][36] , \SUMB[22][35] , \SUMB[22][34] ,
         \SUMB[22][33] , \SUMB[22][32] , \SUMB[22][31] , \SUMB[22][30] ,
         \SUMB[22][29] , \SUMB[22][28] , \SUMB[22][27] , \SUMB[22][26] ,
         \SUMB[22][25] , \SUMB[22][24] , \SUMB[22][23] , \SUMB[22][22] ,
         \SUMB[22][21] , \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] ,
         \SUMB[22][17] , \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] ,
         \SUMB[22][13] , \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] ,
         \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] ,
         \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] ,
         \SUMB[22][1] , \SUMB[21][94] , \SUMB[21][93] , \SUMB[21][92] ,
         \SUMB[21][91] , \SUMB[21][90] , \SUMB[21][89] , \SUMB[21][88] ,
         \SUMB[21][87] , \SUMB[21][86] , \SUMB[21][85] , \SUMB[21][84] ,
         \SUMB[21][83] , \SUMB[21][82] , \SUMB[21][81] , \SUMB[21][80] ,
         \SUMB[21][79] , \SUMB[21][78] , \SUMB[21][77] , \SUMB[21][76] ,
         \SUMB[21][75] , \SUMB[21][74] , \SUMB[21][73] , \SUMB[21][72] ,
         \SUMB[21][71] , \SUMB[21][70] , \SUMB[21][69] , \SUMB[21][68] ,
         \SUMB[21][67] , \SUMB[21][66] , \SUMB[21][65] , \SUMB[21][64] ,
         \SUMB[21][63] , \SUMB[21][62] , \SUMB[21][61] , \SUMB[21][60] ,
         \SUMB[21][59] , \SUMB[21][58] , \SUMB[21][57] , \SUMB[21][56] ,
         \SUMB[21][55] , \SUMB[21][54] , \SUMB[21][53] , \SUMB[21][52] ,
         \SUMB[21][51] , \SUMB[21][50] , \SUMB[21][49] , \SUMB[21][48] ,
         \SUMB[21][47] , \SUMB[21][46] , \SUMB[21][45] , \SUMB[21][44] ,
         \SUMB[21][43] , \SUMB[21][42] , \SUMB[21][41] , \SUMB[21][40] ,
         \SUMB[21][39] , \SUMB[21][38] , \SUMB[21][37] , \SUMB[21][36] ,
         \SUMB[21][35] , \SUMB[21][34] , \SUMB[21][33] , \SUMB[21][32] ,
         \SUMB[21][31] , \SUMB[21][30] , \SUMB[21][29] , \SUMB[21][28] ,
         \SUMB[21][27] , \SUMB[21][26] , \SUMB[21][25] , \SUMB[21][24] ,
         \SUMB[21][23] , \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] ,
         \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] ,
         \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] ,
         \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] ,
         \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] ,
         \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][94] ,
         \SUMB[20][93] , \SUMB[20][92] , \SUMB[20][91] , \SUMB[20][90] ,
         \SUMB[20][89] , \SUMB[20][88] , \SUMB[20][87] , \SUMB[20][86] ,
         \SUMB[20][85] , \SUMB[20][84] , \SUMB[20][83] , \SUMB[20][82] ,
         \SUMB[20][81] , \SUMB[20][80] , \SUMB[20][79] , \SUMB[20][78] ,
         \SUMB[20][77] , \SUMB[20][76] , \SUMB[20][75] , \SUMB[20][74] ,
         \SUMB[20][73] , \SUMB[20][72] , \SUMB[20][71] , \SUMB[20][70] ,
         \SUMB[20][69] , \SUMB[20][68] , \SUMB[20][67] , \SUMB[20][66] ,
         \SUMB[20][65] , \SUMB[20][64] , \SUMB[20][63] , \SUMB[20][62] ,
         \SUMB[20][61] , \SUMB[20][60] , \SUMB[20][59] , \SUMB[20][58] ,
         \SUMB[20][57] , \SUMB[20][56] , \SUMB[20][55] , \SUMB[20][54] ,
         \SUMB[20][53] , \SUMB[20][52] , \SUMB[20][51] , \SUMB[20][50] ,
         \SUMB[20][49] , \SUMB[20][48] , \SUMB[20][47] , \SUMB[20][46] ,
         \SUMB[20][45] , \SUMB[20][44] , \SUMB[20][43] , \SUMB[20][42] ,
         \SUMB[20][41] , \SUMB[20][40] , \SUMB[20][39] , \SUMB[20][38] ,
         \SUMB[20][37] , \SUMB[20][36] , \SUMB[20][35] , \SUMB[20][34] ,
         \SUMB[20][33] , \SUMB[20][32] , \SUMB[20][31] , \SUMB[20][30] ,
         \SUMB[20][29] , \SUMB[20][28] , \SUMB[20][27] , \SUMB[20][26] ,
         \SUMB[20][25] , \SUMB[20][24] , \SUMB[20][23] , \SUMB[20][22] ,
         \SUMB[20][21] , \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] ,
         \SUMB[20][17] , \SUMB[20][16] , \SUMB[20][15] , \SUMB[20][14] ,
         \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] , \SUMB[20][10] ,
         \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] ,
         \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] ,
         \SUMB[20][1] , \SUMB[19][94] , \SUMB[19][93] , \SUMB[19][92] ,
         \SUMB[19][91] , \SUMB[19][90] , \SUMB[19][89] , \SUMB[19][88] ,
         \SUMB[19][87] , \SUMB[19][86] , \SUMB[19][85] , \SUMB[19][84] ,
         \SUMB[19][83] , \SUMB[19][82] , \SUMB[19][81] , \SUMB[19][80] ,
         \SUMB[19][79] , \SUMB[19][78] , \SUMB[19][77] , \SUMB[19][76] ,
         \SUMB[19][75] , \SUMB[19][74] , \SUMB[19][73] , \SUMB[19][72] ,
         \SUMB[19][71] , \SUMB[19][70] , \SUMB[19][69] , \SUMB[19][68] ,
         \SUMB[19][67] , \SUMB[19][66] , \SUMB[19][65] , \SUMB[19][64] ,
         \SUMB[19][63] , \SUMB[19][62] , \SUMB[19][61] , \SUMB[19][60] ,
         \SUMB[19][59] , \SUMB[19][58] , \SUMB[19][57] , \SUMB[19][56] ,
         \SUMB[19][55] , \SUMB[19][54] , \SUMB[19][53] , \SUMB[19][52] ,
         \SUMB[19][51] , \SUMB[19][50] , \SUMB[19][49] , \SUMB[19][48] ,
         \SUMB[19][47] , \SUMB[19][46] , \SUMB[19][45] , \SUMB[19][44] ,
         \SUMB[19][43] , \SUMB[19][42] , \SUMB[19][41] , \SUMB[19][40] ,
         \SUMB[19][39] , \SUMB[19][38] , \SUMB[19][37] , \SUMB[19][36] ,
         \SUMB[19][35] , \SUMB[19][34] , \SUMB[19][33] , \SUMB[19][32] ,
         \CARRYB[29][94] , \CARRYB[29][93] , \CARRYB[29][92] ,
         \CARRYB[29][91] , \CARRYB[29][90] , \CARRYB[29][89] ,
         \CARRYB[29][88] , \CARRYB[29][87] , \CARRYB[29][86] ,
         \CARRYB[29][85] , \CARRYB[29][84] , \CARRYB[29][83] ,
         \CARRYB[29][82] , \CARRYB[29][81] , \CARRYB[29][80] ,
         \CARRYB[29][79] , \CARRYB[29][78] , \CARRYB[29][77] ,
         \CARRYB[29][76] , \CARRYB[29][75] , \CARRYB[29][74] ,
         \CARRYB[29][73] , \CARRYB[29][72] , \CARRYB[29][71] ,
         \CARRYB[29][70] , \CARRYB[29][69] , \CARRYB[29][68] ,
         \CARRYB[29][67] , \CARRYB[29][66] , \CARRYB[29][65] ,
         \CARRYB[29][64] , \CARRYB[29][63] , \CARRYB[29][62] ,
         \CARRYB[29][61] , \CARRYB[29][60] , \CARRYB[29][59] ,
         \CARRYB[29][58] , \CARRYB[29][57] , \CARRYB[29][56] ,
         \CARRYB[29][55] , \CARRYB[29][54] , \CARRYB[29][53] ,
         \CARRYB[29][52] , \CARRYB[29][51] , \CARRYB[29][50] ,
         \CARRYB[29][49] , \CARRYB[29][48] , \CARRYB[29][47] ,
         \CARRYB[29][46] , \CARRYB[29][45] , \CARRYB[29][44] ,
         \CARRYB[29][43] , \CARRYB[29][42] , \CARRYB[29][41] ,
         \CARRYB[29][40] , \CARRYB[29][39] , \CARRYB[29][38] ,
         \CARRYB[29][37] , \CARRYB[29][36] , \CARRYB[29][35] ,
         \CARRYB[29][34] , \CARRYB[29][33] , \CARRYB[29][32] ,
         \CARRYB[29][31] , \CARRYB[29][30] , \CARRYB[29][29] ,
         \CARRYB[29][28] , \CARRYB[29][27] , \CARRYB[29][26] ,
         \CARRYB[29][25] , \CARRYB[29][24] , \CARRYB[29][23] ,
         \CARRYB[29][22] , \CARRYB[29][21] , \CARRYB[29][20] ,
         \CARRYB[29][19] , \CARRYB[29][18] , \CARRYB[29][17] ,
         \CARRYB[29][16] , \CARRYB[29][15] , \CARRYB[29][14] ,
         \CARRYB[29][13] , \CARRYB[29][12] , \CARRYB[29][11] ,
         \CARRYB[29][10] , \CARRYB[29][9] , \CARRYB[29][8] , \CARRYB[29][7] ,
         \CARRYB[29][6] , \CARRYB[29][5] , \CARRYB[29][4] , \CARRYB[29][3] ,
         \CARRYB[29][2] , \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][94] ,
         \CARRYB[28][93] , \CARRYB[28][92] , \CARRYB[28][91] ,
         \CARRYB[28][90] , \CARRYB[28][89] , \CARRYB[28][88] ,
         \CARRYB[28][87] , \CARRYB[28][86] , \CARRYB[28][85] ,
         \CARRYB[28][84] , \CARRYB[28][83] , \CARRYB[28][82] ,
         \CARRYB[28][81] , \CARRYB[28][80] , \CARRYB[28][79] ,
         \CARRYB[28][78] , \CARRYB[28][77] , \CARRYB[28][76] ,
         \CARRYB[28][75] , \CARRYB[28][74] , \CARRYB[28][73] ,
         \CARRYB[28][72] , \CARRYB[28][71] , \CARRYB[28][70] ,
         \CARRYB[28][69] , \CARRYB[28][68] , \CARRYB[28][67] ,
         \CARRYB[28][66] , \CARRYB[28][65] , \CARRYB[28][64] ,
         \CARRYB[28][63] , \CARRYB[28][62] , \CARRYB[28][61] ,
         \CARRYB[28][60] , \CARRYB[28][59] , \CARRYB[28][58] ,
         \CARRYB[28][57] , \CARRYB[28][56] , \CARRYB[28][55] ,
         \CARRYB[28][54] , \CARRYB[28][53] , \CARRYB[28][52] ,
         \CARRYB[28][51] , \CARRYB[28][50] , \CARRYB[28][49] ,
         \CARRYB[28][48] , \CARRYB[28][47] , \CARRYB[28][46] ,
         \CARRYB[28][45] , \CARRYB[28][44] , \CARRYB[28][43] ,
         \CARRYB[28][42] , \CARRYB[28][41] , \CARRYB[28][40] ,
         \CARRYB[28][39] , \CARRYB[28][38] , \CARRYB[28][37] ,
         \CARRYB[28][36] , \CARRYB[28][35] , \CARRYB[28][34] ,
         \CARRYB[28][33] , \CARRYB[28][32] , \CARRYB[28][31] ,
         \CARRYB[28][30] , \CARRYB[28][29] , \CARRYB[28][28] ,
         \CARRYB[28][27] , \CARRYB[28][26] , \CARRYB[28][25] ,
         \CARRYB[28][24] , \CARRYB[28][23] , \CARRYB[28][22] ,
         \CARRYB[28][21] , \CARRYB[28][20] , \CARRYB[28][19] ,
         \CARRYB[28][18] , \CARRYB[28][17] , \CARRYB[28][16] ,
         \CARRYB[28][15] , \CARRYB[28][14] , \CARRYB[28][13] ,
         \CARRYB[28][12] , \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] ,
         \CARRYB[28][8] , \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] ,
         \CARRYB[28][4] , \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][94] , \CARRYB[27][93] , \CARRYB[27][92] ,
         \CARRYB[27][91] , \CARRYB[27][90] , \CARRYB[27][89] ,
         \CARRYB[27][88] , \CARRYB[27][87] , \CARRYB[27][86] ,
         \CARRYB[27][85] , \CARRYB[27][84] , \CARRYB[27][83] ,
         \CARRYB[27][82] , \CARRYB[27][81] , \CARRYB[27][80] ,
         \CARRYB[27][79] , \CARRYB[27][78] , \CARRYB[27][77] ,
         \CARRYB[27][76] , \CARRYB[27][75] , \CARRYB[27][74] ,
         \CARRYB[27][73] , \CARRYB[27][72] , \CARRYB[27][71] ,
         \CARRYB[27][70] , \CARRYB[27][69] , \CARRYB[27][68] ,
         \CARRYB[27][67] , \CARRYB[27][66] , \CARRYB[27][65] ,
         \CARRYB[27][64] , \CARRYB[27][63] , \CARRYB[27][62] ,
         \CARRYB[27][61] , \CARRYB[27][60] , \CARRYB[27][59] ,
         \CARRYB[27][58] , \CARRYB[27][57] , \CARRYB[27][56] ,
         \CARRYB[27][55] , \CARRYB[27][54] , \CARRYB[27][53] ,
         \CARRYB[27][52] , \CARRYB[27][51] , \CARRYB[27][50] ,
         \CARRYB[27][49] , \CARRYB[27][48] , \CARRYB[27][47] ,
         \CARRYB[27][46] , \CARRYB[27][45] , \CARRYB[27][44] ,
         \CARRYB[27][43] , \CARRYB[27][42] , \CARRYB[27][41] ,
         \CARRYB[27][40] , \CARRYB[27][39] , \CARRYB[27][38] ,
         \CARRYB[27][37] , \CARRYB[27][36] , \CARRYB[27][35] ,
         \CARRYB[27][34] , \CARRYB[27][33] , \CARRYB[27][32] ,
         \CARRYB[27][31] , \CARRYB[27][30] , \CARRYB[27][29] ,
         \CARRYB[27][28] , \CARRYB[27][27] , \CARRYB[27][26] ,
         \CARRYB[27][25] , \CARRYB[27][24] , \CARRYB[27][23] ,
         \CARRYB[27][22] , \CARRYB[27][21] , \CARRYB[27][20] ,
         \CARRYB[27][19] , \CARRYB[27][18] , \CARRYB[27][17] ,
         \CARRYB[27][16] , \CARRYB[27][15] , \CARRYB[27][14] ,
         \CARRYB[27][13] , \CARRYB[27][12] , \CARRYB[27][11] ,
         \CARRYB[27][10] , \CARRYB[27][9] , \CARRYB[27][8] , \CARRYB[27][7] ,
         \CARRYB[27][6] , \CARRYB[27][5] , \CARRYB[27][4] , \CARRYB[27][3] ,
         \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] , \CARRYB[26][94] ,
         \CARRYB[26][93] , \CARRYB[26][92] , \CARRYB[26][91] ,
         \CARRYB[26][90] , \CARRYB[26][89] , \CARRYB[26][88] ,
         \CARRYB[26][87] , \CARRYB[26][86] , \CARRYB[26][85] ,
         \CARRYB[26][84] , \CARRYB[26][83] , \CARRYB[26][82] ,
         \CARRYB[26][81] , \CARRYB[26][80] , \CARRYB[26][79] ,
         \CARRYB[26][78] , \CARRYB[26][77] , \CARRYB[26][76] ,
         \CARRYB[26][75] , \CARRYB[26][74] , \CARRYB[26][73] ,
         \CARRYB[26][72] , \CARRYB[26][71] , \CARRYB[26][70] ,
         \CARRYB[26][69] , \CARRYB[26][68] , \CARRYB[26][67] ,
         \CARRYB[26][66] , \CARRYB[26][65] , \CARRYB[26][64] ,
         \CARRYB[26][63] , \CARRYB[26][62] , \CARRYB[26][61] ,
         \CARRYB[26][60] , \CARRYB[26][59] , \CARRYB[26][58] ,
         \CARRYB[26][57] , \CARRYB[26][56] , \CARRYB[26][55] ,
         \CARRYB[26][54] , \CARRYB[26][53] , \CARRYB[26][52] ,
         \CARRYB[26][51] , \CARRYB[26][50] , \CARRYB[26][49] ,
         \CARRYB[26][48] , \CARRYB[26][47] , \CARRYB[26][46] ,
         \CARRYB[26][45] , \CARRYB[26][44] , \CARRYB[26][43] ,
         \CARRYB[26][42] , \CARRYB[26][41] , \CARRYB[26][40] ,
         \CARRYB[26][39] , \CARRYB[26][38] , \CARRYB[26][37] ,
         \CARRYB[26][36] , \CARRYB[26][35] , \CARRYB[26][34] ,
         \CARRYB[26][33] , \CARRYB[26][32] , \CARRYB[26][31] ,
         \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][94] , \CARRYB[25][93] , \CARRYB[25][92] ,
         \CARRYB[25][91] , \CARRYB[25][90] , \CARRYB[25][89] ,
         \CARRYB[25][88] , \CARRYB[25][87] , \CARRYB[25][86] ,
         \CARRYB[25][85] , \CARRYB[25][84] , \CARRYB[25][83] ,
         \CARRYB[25][82] , \CARRYB[25][81] , \CARRYB[25][80] ,
         \CARRYB[25][79] , \CARRYB[25][78] , \CARRYB[25][77] ,
         \CARRYB[25][76] , \CARRYB[25][75] , \CARRYB[25][74] ,
         \CARRYB[25][73] , \CARRYB[25][72] , \CARRYB[25][71] ,
         \CARRYB[25][70] , \CARRYB[25][69] , \CARRYB[25][68] ,
         \CARRYB[25][67] , \CARRYB[25][66] , \CARRYB[25][65] ,
         \CARRYB[25][64] , \CARRYB[25][63] , \CARRYB[25][62] ,
         \CARRYB[25][61] , \CARRYB[25][60] , \CARRYB[25][59] ,
         \CARRYB[25][58] , \CARRYB[25][57] , \CARRYB[25][56] ,
         \CARRYB[25][55] , \CARRYB[25][54] , \CARRYB[25][53] ,
         \CARRYB[25][52] , \CARRYB[25][51] , \CARRYB[25][50] ,
         \CARRYB[25][49] , \CARRYB[25][48] , \CARRYB[25][47] ,
         \CARRYB[25][46] , \CARRYB[25][45] , \CARRYB[25][44] ,
         \CARRYB[25][43] , \CARRYB[25][42] , \CARRYB[25][41] ,
         \CARRYB[25][40] , \CARRYB[25][39] , \CARRYB[25][38] ,
         \CARRYB[25][37] , \CARRYB[25][36] , \CARRYB[25][35] ,
         \CARRYB[25][34] , \CARRYB[25][33] , \CARRYB[25][32] ,
         \CARRYB[25][31] , \CARRYB[25][30] , \CARRYB[25][29] ,
         \CARRYB[25][28] , \CARRYB[25][27] , \CARRYB[25][26] ,
         \CARRYB[25][25] , \CARRYB[25][24] , \CARRYB[25][23] ,
         \CARRYB[25][22] , \CARRYB[25][21] , \CARRYB[25][20] ,
         \CARRYB[25][19] , \CARRYB[25][18] , \CARRYB[25][17] ,
         \CARRYB[25][16] , \CARRYB[25][15] , \CARRYB[25][14] ,
         \CARRYB[25][13] , \CARRYB[25][12] , \CARRYB[25][11] ,
         \CARRYB[25][10] , \CARRYB[25][9] , \CARRYB[25][8] , \CARRYB[25][7] ,
         \CARRYB[25][6] , \CARRYB[25][5] , \CARRYB[25][4] , \CARRYB[25][3] ,
         \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] , \CARRYB[24][94] ,
         \CARRYB[24][93] , \CARRYB[24][92] , \CARRYB[24][91] ,
         \CARRYB[24][90] , \CARRYB[24][89] , \CARRYB[24][88] ,
         \CARRYB[24][87] , \CARRYB[24][86] , \CARRYB[24][85] ,
         \CARRYB[24][84] , \CARRYB[24][83] , \CARRYB[24][82] ,
         \CARRYB[24][81] , \CARRYB[24][80] , \CARRYB[24][79] ,
         \CARRYB[24][78] , \CARRYB[24][77] , \CARRYB[24][76] ,
         \CARRYB[24][75] , \CARRYB[24][74] , \CARRYB[24][73] ,
         \CARRYB[24][72] , \CARRYB[24][71] , \CARRYB[24][70] ,
         \CARRYB[24][69] , \CARRYB[24][68] , \CARRYB[24][67] ,
         \CARRYB[24][66] , \CARRYB[24][65] , \CARRYB[24][64] , \SUMB[29][94] ,
         \SUMB[29][93] , \SUMB[29][92] , \SUMB[29][91] , \SUMB[29][90] ,
         \SUMB[29][89] , \SUMB[29][88] , \SUMB[29][87] , \SUMB[29][86] ,
         \SUMB[29][85] , \SUMB[29][84] , \SUMB[29][83] , \SUMB[29][82] ,
         \SUMB[29][81] , \SUMB[29][80] , \SUMB[29][79] , \SUMB[29][78] ,
         \SUMB[29][77] , \SUMB[29][76] , \SUMB[29][75] , \SUMB[29][74] ,
         \SUMB[29][73] , \SUMB[29][72] , \SUMB[29][71] , \SUMB[29][70] ,
         \SUMB[29][69] , \SUMB[29][68] , \SUMB[29][67] , \SUMB[29][66] ,
         \SUMB[29][65] , \SUMB[29][64] , \SUMB[29][63] , \SUMB[29][62] ,
         \SUMB[29][61] , \SUMB[29][60] , \SUMB[29][59] , \SUMB[29][58] ,
         \SUMB[29][57] , \SUMB[29][56] , \SUMB[29][55] , \SUMB[29][54] ,
         \SUMB[29][53] , \SUMB[29][52] , \SUMB[29][51] , \SUMB[29][50] ,
         \SUMB[29][49] , \SUMB[29][48] , \SUMB[29][47] , \SUMB[29][46] ,
         \SUMB[29][45] , \SUMB[29][44] , \SUMB[29][43] , \SUMB[29][42] ,
         \SUMB[29][41] , \SUMB[29][40] , \SUMB[29][39] , \SUMB[29][38] ,
         \SUMB[29][37] , \SUMB[29][36] , \SUMB[29][35] , \SUMB[29][34] ,
         \SUMB[29][33] , \SUMB[29][32] , \SUMB[29][31] , \SUMB[29][30] ,
         \SUMB[29][29] , \SUMB[29][28] , \SUMB[29][27] , \SUMB[29][26] ,
         \SUMB[29][25] , \SUMB[29][24] , \SUMB[29][23] , \SUMB[29][22] ,
         \SUMB[29][21] , \SUMB[29][20] , \SUMB[29][19] , \SUMB[29][18] ,
         \SUMB[29][17] , \SUMB[29][16] , \SUMB[29][15] , \SUMB[29][14] ,
         \SUMB[29][13] , \SUMB[29][12] , \SUMB[29][11] , \SUMB[29][10] ,
         \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] , \SUMB[29][6] ,
         \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] , \SUMB[29][2] ,
         \SUMB[29][1] , \SUMB[29][0] , \SUMB[28][94] , \SUMB[28][93] ,
         \SUMB[28][92] , \SUMB[28][91] , \SUMB[28][90] , \SUMB[28][89] ,
         \SUMB[28][88] , \SUMB[28][87] , \SUMB[28][86] , \SUMB[28][85] ,
         \SUMB[28][84] , \SUMB[28][83] , \SUMB[28][82] , \SUMB[28][81] ,
         \SUMB[28][80] , \SUMB[28][79] , \SUMB[28][78] , \SUMB[28][77] ,
         \SUMB[28][76] , \SUMB[28][75] , \SUMB[28][74] , \SUMB[28][73] ,
         \SUMB[28][72] , \SUMB[28][71] , \SUMB[28][70] , \SUMB[28][69] ,
         \SUMB[28][68] , \SUMB[28][67] , \SUMB[28][66] , \SUMB[28][65] ,
         \SUMB[28][64] , \SUMB[28][63] , \SUMB[28][62] , \SUMB[28][61] ,
         \SUMB[28][60] , \SUMB[28][59] , \SUMB[28][58] , \SUMB[28][57] ,
         \SUMB[28][56] , \SUMB[28][55] , \SUMB[28][54] , \SUMB[28][53] ,
         \SUMB[28][52] , \SUMB[28][51] , \SUMB[28][50] , \SUMB[28][49] ,
         \SUMB[28][48] , \SUMB[28][47] , \SUMB[28][46] , \SUMB[28][45] ,
         \SUMB[28][44] , \SUMB[28][43] , \SUMB[28][42] , \SUMB[28][41] ,
         \SUMB[28][40] , \SUMB[28][39] , \SUMB[28][38] , \SUMB[28][37] ,
         \SUMB[28][36] , \SUMB[28][35] , \SUMB[28][34] , \SUMB[28][33] ,
         \SUMB[28][32] , \SUMB[28][31] , \SUMB[28][30] , \SUMB[28][29] ,
         \SUMB[28][28] , \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] ,
         \SUMB[28][24] , \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] ,
         \SUMB[28][20] , \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] ,
         \SUMB[28][16] , \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] ,
         \SUMB[28][12] , \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] ,
         \SUMB[28][8] , \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] ,
         \SUMB[28][4] , \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] ,
         \SUMB[27][94] , \SUMB[27][93] , \SUMB[27][92] , \SUMB[27][91] ,
         \SUMB[27][90] , \SUMB[27][89] , \SUMB[27][88] , \SUMB[27][87] ,
         \SUMB[27][86] , \SUMB[27][85] , \SUMB[27][84] , \SUMB[27][83] ,
         \SUMB[27][82] , \SUMB[27][81] , \SUMB[27][80] , \SUMB[27][79] ,
         \SUMB[27][78] , \SUMB[27][77] , \SUMB[27][76] , \SUMB[27][75] ,
         \SUMB[27][74] , \SUMB[27][73] , \SUMB[27][72] , \SUMB[27][71] ,
         \SUMB[27][70] , \SUMB[27][69] , \SUMB[27][68] , \SUMB[27][67] ,
         \SUMB[27][66] , \SUMB[27][65] , \SUMB[27][64] , \SUMB[27][63] ,
         \SUMB[27][62] , \SUMB[27][61] , \SUMB[27][60] , \SUMB[27][59] ,
         \SUMB[27][58] , \SUMB[27][57] , \SUMB[27][56] , \SUMB[27][55] ,
         \SUMB[27][54] , \SUMB[27][53] , \SUMB[27][52] , \SUMB[27][51] ,
         \SUMB[27][50] , \SUMB[27][49] , \SUMB[27][48] , \SUMB[27][47] ,
         \SUMB[27][46] , \SUMB[27][45] , \SUMB[27][44] , \SUMB[27][43] ,
         \SUMB[27][42] , \SUMB[27][41] , \SUMB[27][40] , \SUMB[27][39] ,
         \SUMB[27][38] , \SUMB[27][37] , \SUMB[27][36] , \SUMB[27][35] ,
         \SUMB[27][34] , \SUMB[27][33] , \SUMB[27][32] , \SUMB[27][31] ,
         \SUMB[27][30] , \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] ,
         \SUMB[27][26] , \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] ,
         \SUMB[27][22] , \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] ,
         \SUMB[27][18] , \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] ,
         \SUMB[27][14] , \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] ,
         \SUMB[27][10] , \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] ,
         \SUMB[27][6] , \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][94] , \SUMB[26][93] ,
         \SUMB[26][92] , \SUMB[26][91] , \SUMB[26][90] , \SUMB[26][89] ,
         \SUMB[26][88] , \SUMB[26][87] , \SUMB[26][86] , \SUMB[26][85] ,
         \SUMB[26][84] , \SUMB[26][83] , \SUMB[26][82] , \SUMB[26][81] ,
         \SUMB[26][80] , \SUMB[26][79] , \SUMB[26][78] , \SUMB[26][77] ,
         \SUMB[26][76] , \SUMB[26][75] , \SUMB[26][74] , \SUMB[26][73] ,
         \SUMB[26][72] , \SUMB[26][71] , \SUMB[26][70] , \SUMB[26][69] ,
         \SUMB[26][68] , \SUMB[26][67] , \SUMB[26][66] , \SUMB[26][65] ,
         \SUMB[26][64] , \SUMB[26][63] , \SUMB[26][62] , \SUMB[26][61] ,
         \SUMB[26][60] , \SUMB[26][59] , \SUMB[26][58] , \SUMB[26][57] ,
         \SUMB[26][56] , \SUMB[26][55] , \SUMB[26][54] , \SUMB[26][53] ,
         \SUMB[26][52] , \SUMB[26][51] , \SUMB[26][50] , \SUMB[26][49] ,
         \SUMB[26][48] , \SUMB[26][47] , \SUMB[26][46] , \SUMB[26][45] ,
         \SUMB[26][44] , \SUMB[26][43] , \SUMB[26][42] , \SUMB[26][41] ,
         \SUMB[26][40] , \SUMB[26][39] , \SUMB[26][38] , \SUMB[26][37] ,
         \SUMB[26][36] , \SUMB[26][35] , \SUMB[26][34] , \SUMB[26][33] ,
         \SUMB[26][32] , \SUMB[26][31] , \SUMB[26][30] , \SUMB[26][29] ,
         \SUMB[26][28] , \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] ,
         \SUMB[26][24] , \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] ,
         \SUMB[26][20] , \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] ,
         \SUMB[26][16] , \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] ,
         \SUMB[26][12] , \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] ,
         \SUMB[26][8] , \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] ,
         \SUMB[26][4] , \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] ,
         \SUMB[25][94] , \SUMB[25][93] , \SUMB[25][92] , \SUMB[25][91] ,
         \SUMB[25][90] , \SUMB[25][89] , \SUMB[25][88] , \SUMB[25][87] ,
         \SUMB[25][86] , \SUMB[25][85] , \SUMB[25][84] , \SUMB[25][83] ,
         \SUMB[25][82] , \SUMB[25][81] , \SUMB[25][80] , \SUMB[25][79] ,
         \SUMB[25][78] , \SUMB[25][77] , \SUMB[25][76] , \SUMB[25][75] ,
         \SUMB[25][74] , \SUMB[25][73] , \SUMB[25][72] , \SUMB[25][71] ,
         \SUMB[25][70] , \SUMB[25][69] , \SUMB[25][68] , \SUMB[25][67] ,
         \SUMB[25][66] , \SUMB[25][65] , \SUMB[25][64] , \SUMB[25][63] ,
         \SUMB[25][62] , \SUMB[25][61] , \SUMB[25][60] , \SUMB[25][59] ,
         \SUMB[25][58] , \SUMB[25][57] , \SUMB[25][56] , \SUMB[25][55] ,
         \SUMB[25][54] , \SUMB[25][53] , \SUMB[25][52] , \SUMB[25][51] ,
         \SUMB[25][50] , \SUMB[25][49] , \SUMB[25][48] , \SUMB[25][47] ,
         \SUMB[25][46] , \SUMB[25][45] , \SUMB[25][44] , \SUMB[25][43] ,
         \SUMB[25][42] , \SUMB[25][41] , \SUMB[25][40] , \SUMB[25][39] ,
         \SUMB[25][38] , \SUMB[25][37] , \SUMB[25][36] , \SUMB[25][35] ,
         \SUMB[25][34] , \SUMB[25][33] , \SUMB[25][32] , \SUMB[25][31] ,
         \SUMB[25][30] , \SUMB[25][29] , \SUMB[25][28] , \SUMB[25][27] ,
         \SUMB[25][26] , \SUMB[25][25] , \SUMB[25][24] , \SUMB[25][23] ,
         \SUMB[25][22] , \SUMB[25][21] , \SUMB[25][20] , \SUMB[25][19] ,
         \SUMB[25][18] , \SUMB[25][17] , \SUMB[25][16] , \SUMB[25][15] ,
         \SUMB[25][14] , \SUMB[25][13] , \SUMB[25][12] , \SUMB[25][11] ,
         \SUMB[25][10] , \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] ,
         \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] ,
         \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][94] , \SUMB[24][93] ,
         \SUMB[24][92] , \SUMB[24][91] , \SUMB[24][90] , \SUMB[24][89] ,
         \SUMB[24][88] , \SUMB[24][87] , \SUMB[24][86] , \SUMB[24][85] ,
         \SUMB[24][84] , \SUMB[24][83] , \SUMB[24][82] , \SUMB[24][81] ,
         \SUMB[24][80] , \SUMB[24][79] , \SUMB[24][78] , \SUMB[24][77] ,
         \SUMB[24][76] , \SUMB[24][75] , \SUMB[24][74] , \SUMB[24][73] ,
         \SUMB[24][72] , \SUMB[24][71] , \SUMB[24][70] , \SUMB[24][69] ,
         \SUMB[24][68] , \SUMB[24][67] , \SUMB[24][66] , \SUMB[24][65] ,
         \SUMB[24][64] , \A1[122] , \A1[121] , \A1[120] , \A1[119] , \A1[118] ,
         \A1[117] , \A1[116] , \A1[115] , \A1[114] , \A1[113] , \A1[112] ,
         \A1[111] , \A1[110] , \A1[109] , \A1[108] , \A1[107] , \A1[106] ,
         \A1[105] , \A1[104] , \A1[103] , \A1[102] , \A1[101] , \A1[100] ,
         \A1[99] , \A1[98] , \A1[97] , \A1[96] , \A1[95] , \A1[94] , \A1[93] ,
         \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] ,
         \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] ,
         \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] ,
         \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] ,
         \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] ,
         \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] ,
         \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] ,
         \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] ,
         \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] ,
         \A1[29] , \A1[28] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[123] , \A2[122] , \A2[121] , \A2[120] , \A2[119] ,
         \A2[118] , \A2[117] , \A2[116] , \A2[115] , \A2[114] , \A2[113] ,
         \A2[112] , \A2[111] , \A2[110] , \A2[109] , \A2[108] , \A2[107] ,
         \A2[106] , \A2[105] , \A2[104] , \A2[103] , \A2[102] , \A2[101] ,
         \A2[100] , \A2[99] , \A2[98] , \A2[97] , \A2[96] , \A2[95] , \A2[94] ,
         \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] ,
         \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] ,
         \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] ,
         \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] ,
         \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] ,
         \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] ,
         \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         \A2[30] , \A2[29] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93;

  LOG_POLY_DW01_add_6 FS_1 ( .A({1'b0, \A1[122] , \A1[121] , \A1[120] , 
        \A1[119] , \A1[118] , \A1[117] , \A1[116] , \A1[115] , \A1[114] , 
        \A1[113] , \A1[112] , \A1[111] , \A1[110] , \A1[109] , \A1[108] , 
        \A1[107] , \A1[106] , \A1[105] , \A1[104] , \A1[103] , \A1[102] , 
        \A1[101] , \A1[100] , \A1[99] , \A1[98] , \A1[97] , \A1[96] , \A1[95] , 
        \A1[94] , \A1[93] , \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , 
        \A1[87] , \A1[86] , \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , 
        \A1[80] , \A1[79] , \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , 
        \A1[73] , \A1[72] , \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , 
        \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , 
        \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , 
        \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , 
        \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , 
        \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , 
        \A1[31] , \A1[30] , \A1[29] , \A1[28] , \SUMB[29][0] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[123] , 
        \A2[122] , \A2[121] , \A2[120] , \A2[119] , \A2[118] , \A2[117] , 
        \A2[116] , \A2[115] , \A2[114] , \A2[113] , \A2[112] , \A2[111] , 
        \A2[110] , \A2[109] , \A2[108] , \A2[107] , \A2[106] , \A2[105] , 
        \A2[104] , \A2[103] , \A2[102] , \A2[101] , \A2[100] , \A2[99] , 
        \A2[98] , \A2[97] , \A2[96] , \A2[95] , \A2[94] , \A2[93] , \A2[92] , 
        \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] , \A2[86] , \A2[85] , 
        \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] , \A2[79] , \A2[78] , 
        \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] , \A2[72] , \A2[71] , 
        \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] , \A2[65] , \A2[64] , 
        \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , \A2[57] , 
        \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , 
        \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] , \A2[44] , \A2[43] , 
        \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , 
        \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , \A2[29] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, PRODUCT[118:89], SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93}) );
  FA1A S2_14_57 ( .A(\ab[14][57] ), .B(\CARRYB[13][57] ), .CI(\SUMB[13][58] ), 
        .CO(\CARRYB[14][57] ), .S(\SUMB[14][57] ) );
  FA1A S2_13_57 ( .A(\ab[13][57] ), .B(\CARRYB[12][57] ), .CI(\SUMB[12][58] ), 
        .CO(\CARRYB[13][57] ), .S(\SUMB[13][57] ) );
  FA1A S2_12_57 ( .A(\ab[12][57] ), .B(\CARRYB[11][57] ), .CI(\SUMB[11][58] ), 
        .CO(\CARRYB[12][57] ), .S(\SUMB[12][57] ) );
  FA1A S2_11_57 ( .A(\ab[11][57] ), .B(\CARRYB[10][57] ), .CI(\SUMB[10][58] ), 
        .CO(\CARRYB[11][57] ), .S(\SUMB[11][57] ) );
  FA1A S2_10_57 ( .A(\ab[10][57] ), .B(\CARRYB[9][57] ), .CI(\SUMB[9][58] ), 
        .CO(\CARRYB[10][57] ), .S(\SUMB[10][57] ) );
  FA1A S2_9_57 ( .A(\ab[9][57] ), .B(\CARRYB[8][57] ), .CI(\SUMB[8][58] ), 
        .CO(\CARRYB[9][57] ), .S(\SUMB[9][57] ) );
  FA1A S2_8_57 ( .A(\ab[8][57] ), .B(\CARRYB[7][57] ), .CI(\SUMB[7][58] ), 
        .CO(\CARRYB[8][57] ), .S(\SUMB[8][57] ) );
  FA1A S2_7_57 ( .A(\ab[7][57] ), .B(\CARRYB[6][57] ), .CI(\SUMB[6][58] ), 
        .CO(\CARRYB[7][57] ), .S(\SUMB[7][57] ) );
  FA1A S2_6_57 ( .A(\ab[6][57] ), .B(\CARRYB[5][57] ), .CI(\SUMB[5][58] ), 
        .CO(\CARRYB[6][57] ), .S(\SUMB[6][57] ) );
  FA1A S2_5_57 ( .A(\ab[5][57] ), .B(\CARRYB[4][57] ), .CI(\SUMB[4][58] ), 
        .CO(\CARRYB[5][57] ), .S(\SUMB[5][57] ) );
  FA1A S2_4_57 ( .A(\ab[4][57] ), .B(\CARRYB[3][57] ), .CI(\SUMB[3][58] ), 
        .CO(\CARRYB[4][57] ), .S(\SUMB[4][57] ) );
  FA1A S2_3_57 ( .A(\ab[3][57] ), .B(\CARRYB[2][57] ), .CI(\SUMB[2][58] ), 
        .CO(\CARRYB[3][57] ), .S(\SUMB[3][57] ) );
  FA1A S2_2_57 ( .A(\ab[2][57] ), .B(\CARRYB[1][57] ), .CI(\SUMB[1][58] ), 
        .CO(\CARRYB[2][57] ), .S(\SUMB[2][57] ) );
  FA1A S2_14_56 ( .A(\ab[14][56] ), .B(\CARRYB[13][56] ), .CI(\SUMB[13][57] ), 
        .CO(\CARRYB[14][56] ), .S(\SUMB[14][56] ) );
  FA1A S2_14_54 ( .A(\ab[14][54] ), .B(\CARRYB[13][54] ), .CI(\SUMB[13][55] ), 
        .CO(\CARRYB[14][54] ), .S(\SUMB[14][54] ) );
  FA1A S2_14_53 ( .A(\ab[14][53] ), .B(\CARRYB[13][53] ), .CI(\SUMB[13][54] ), 
        .CO(\CARRYB[14][53] ), .S(\SUMB[14][53] ) );
  FA1A S2_14_59 ( .A(\ab[14][59] ), .B(\CARRYB[13][59] ), .CI(\SUMB[13][60] ), 
        .CO(\CARRYB[14][59] ), .S(\SUMB[14][59] ) );
  FA1A S2_14_58 ( .A(\ab[14][58] ), .B(\CARRYB[13][58] ), .CI(\SUMB[13][59] ), 
        .CO(\CARRYB[14][58] ), .S(\SUMB[14][58] ) );
  FA1A S2_13_58 ( .A(\ab[13][58] ), .B(\CARRYB[12][58] ), .CI(\SUMB[12][59] ), 
        .CO(\CARRYB[13][58] ), .S(\SUMB[13][58] ) );
  FA1A S2_13_56 ( .A(\ab[13][56] ), .B(\CARRYB[12][56] ), .CI(\SUMB[12][57] ), 
        .CO(\CARRYB[13][56] ), .S(\SUMB[13][56] ) );
  FA1A S2_13_54 ( .A(\ab[13][54] ), .B(\CARRYB[12][54] ), .CI(\SUMB[12][55] ), 
        .CO(\CARRYB[13][54] ), .S(\SUMB[13][54] ) );
  FA1A S2_13_53 ( .A(\ab[13][53] ), .B(\CARRYB[12][53] ), .CI(\SUMB[12][54] ), 
        .CO(\CARRYB[13][53] ), .S(\SUMB[13][53] ) );
  FA1A S2_13_59 ( .A(\ab[13][59] ), .B(\CARRYB[12][59] ), .CI(\SUMB[12][60] ), 
        .CO(\CARRYB[13][59] ), .S(\SUMB[13][59] ) );
  FA1A S2_12_59 ( .A(\ab[12][59] ), .B(\CARRYB[11][59] ), .CI(\SUMB[11][60] ), 
        .CO(\CARRYB[12][59] ), .S(\SUMB[12][59] ) );
  FA1A S2_12_58 ( .A(\ab[12][58] ), .B(\CARRYB[11][58] ), .CI(\SUMB[11][59] ), 
        .CO(\CARRYB[12][58] ), .S(\SUMB[12][58] ) );
  FA1A S2_12_56 ( .A(\ab[12][56] ), .B(\CARRYB[11][56] ), .CI(\SUMB[11][57] ), 
        .CO(\CARRYB[12][56] ), .S(\SUMB[12][56] ) );
  FA1A S2_12_54 ( .A(\ab[12][54] ), .B(\CARRYB[11][54] ), .CI(\SUMB[11][55] ), 
        .CO(\CARRYB[12][54] ), .S(\SUMB[12][54] ) );
  FA1A S2_12_53 ( .A(\ab[12][53] ), .B(\CARRYB[11][53] ), .CI(\SUMB[11][54] ), 
        .CO(\CARRYB[12][53] ), .S(\SUMB[12][53] ) );
  FA1A S2_11_59 ( .A(\ab[11][59] ), .B(\CARRYB[10][59] ), .CI(\SUMB[10][60] ), 
        .CO(\CARRYB[11][59] ), .S(\SUMB[11][59] ) );
  FA1A S2_11_58 ( .A(\ab[11][58] ), .B(\CARRYB[10][58] ), .CI(\SUMB[10][59] ), 
        .CO(\CARRYB[11][58] ), .S(\SUMB[11][58] ) );
  FA1A S2_11_56 ( .A(\ab[11][56] ), .B(\CARRYB[10][56] ), .CI(\SUMB[10][57] ), 
        .CO(\CARRYB[11][56] ), .S(\SUMB[11][56] ) );
  FA1A S2_11_54 ( .A(\ab[11][54] ), .B(\CARRYB[10][54] ), .CI(\SUMB[10][55] ), 
        .CO(\CARRYB[11][54] ), .S(\SUMB[11][54] ) );
  FA1A S2_11_53 ( .A(\ab[11][53] ), .B(\CARRYB[10][53] ), .CI(\SUMB[10][54] ), 
        .CO(\CARRYB[11][53] ), .S(\SUMB[11][53] ) );
  FA1A S2_10_59 ( .A(\ab[10][59] ), .B(\CARRYB[9][59] ), .CI(\SUMB[9][60] ), 
        .CO(\CARRYB[10][59] ), .S(\SUMB[10][59] ) );
  FA1A S2_10_58 ( .A(\ab[10][58] ), .B(\CARRYB[9][58] ), .CI(\SUMB[9][59] ), 
        .CO(\CARRYB[10][58] ), .S(\SUMB[10][58] ) );
  FA1A S2_10_56 ( .A(\ab[10][56] ), .B(\CARRYB[9][56] ), .CI(\SUMB[9][57] ), 
        .CO(\CARRYB[10][56] ), .S(\SUMB[10][56] ) );
  FA1A S2_10_54 ( .A(\ab[10][54] ), .B(\CARRYB[9][54] ), .CI(\SUMB[9][55] ), 
        .CO(\CARRYB[10][54] ), .S(\SUMB[10][54] ) );
  FA1A S2_10_53 ( .A(\ab[10][53] ), .B(\CARRYB[9][53] ), .CI(\SUMB[9][54] ), 
        .CO(\CARRYB[10][53] ), .S(\SUMB[10][53] ) );
  FA1A S2_9_59 ( .A(\ab[9][59] ), .B(\CARRYB[8][59] ), .CI(\SUMB[8][60] ), 
        .CO(\CARRYB[9][59] ), .S(\SUMB[9][59] ) );
  FA1A S2_9_58 ( .A(\ab[9][58] ), .B(\CARRYB[8][58] ), .CI(\SUMB[8][59] ), 
        .CO(\CARRYB[9][58] ), .S(\SUMB[9][58] ) );
  FA1A S2_9_56 ( .A(\ab[9][56] ), .B(\CARRYB[8][56] ), .CI(\SUMB[8][57] ), 
        .CO(\CARRYB[9][56] ), .S(\SUMB[9][56] ) );
  FA1A S2_9_54 ( .A(\ab[9][54] ), .B(\CARRYB[8][54] ), .CI(\SUMB[8][55] ), 
        .CO(\CARRYB[9][54] ), .S(\SUMB[9][54] ) );
  FA1A S2_9_53 ( .A(\ab[9][53] ), .B(\CARRYB[8][53] ), .CI(\SUMB[8][54] ), 
        .CO(\CARRYB[9][53] ), .S(\SUMB[9][53] ) );
  FA1A S2_8_59 ( .A(\ab[8][59] ), .B(\CARRYB[7][59] ), .CI(\SUMB[7][60] ), 
        .CO(\CARRYB[8][59] ), .S(\SUMB[8][59] ) );
  FA1A S2_8_58 ( .A(\ab[8][58] ), .B(\CARRYB[7][58] ), .CI(\SUMB[7][59] ), 
        .CO(\CARRYB[8][58] ), .S(\SUMB[8][58] ) );
  FA1A S2_8_56 ( .A(\ab[8][56] ), .B(\CARRYB[7][56] ), .CI(\SUMB[7][57] ), 
        .CO(\CARRYB[8][56] ), .S(\SUMB[8][56] ) );
  FA1A S2_8_54 ( .A(\ab[8][54] ), .B(\CARRYB[7][54] ), .CI(\SUMB[7][55] ), 
        .CO(\CARRYB[8][54] ), .S(\SUMB[8][54] ) );
  FA1A S2_8_53 ( .A(\ab[8][53] ), .B(\CARRYB[7][53] ), .CI(\SUMB[7][54] ), 
        .CO(\CARRYB[8][53] ), .S(\SUMB[8][53] ) );
  FA1A S2_7_59 ( .A(\ab[7][59] ), .B(\CARRYB[6][59] ), .CI(\SUMB[6][60] ), 
        .CO(\CARRYB[7][59] ), .S(\SUMB[7][59] ) );
  FA1A S2_7_58 ( .A(\ab[7][58] ), .B(\CARRYB[6][58] ), .CI(\SUMB[6][59] ), 
        .CO(\CARRYB[7][58] ), .S(\SUMB[7][58] ) );
  FA1A S2_7_56 ( .A(\ab[7][56] ), .B(\CARRYB[6][56] ), .CI(\SUMB[6][57] ), 
        .CO(\CARRYB[7][56] ), .S(\SUMB[7][56] ) );
  FA1A S2_7_54 ( .A(\ab[7][54] ), .B(\CARRYB[6][54] ), .CI(\SUMB[6][55] ), 
        .CO(\CARRYB[7][54] ), .S(\SUMB[7][54] ) );
  FA1A S2_7_53 ( .A(\ab[7][53] ), .B(\CARRYB[6][53] ), .CI(\SUMB[6][54] ), 
        .CO(\CARRYB[7][53] ), .S(\SUMB[7][53] ) );
  FA1A S2_6_59 ( .A(\ab[6][59] ), .B(\CARRYB[5][59] ), .CI(\SUMB[5][60] ), 
        .CO(\CARRYB[6][59] ), .S(\SUMB[6][59] ) );
  FA1A S2_6_58 ( .A(\ab[6][58] ), .B(\CARRYB[5][58] ), .CI(\SUMB[5][59] ), 
        .CO(\CARRYB[6][58] ), .S(\SUMB[6][58] ) );
  FA1A S2_6_56 ( .A(\ab[6][56] ), .B(\CARRYB[5][56] ), .CI(\SUMB[5][57] ), 
        .CO(\CARRYB[6][56] ), .S(\SUMB[6][56] ) );
  FA1A S2_6_54 ( .A(\ab[6][54] ), .B(\CARRYB[5][54] ), .CI(\SUMB[5][55] ), 
        .CO(\CARRYB[6][54] ), .S(\SUMB[6][54] ) );
  FA1A S2_6_53 ( .A(\ab[6][53] ), .B(\CARRYB[5][53] ), .CI(\SUMB[5][54] ), 
        .CO(\CARRYB[6][53] ), .S(\SUMB[6][53] ) );
  FA1A S2_5_59 ( .A(\ab[5][59] ), .B(\CARRYB[4][59] ), .CI(\SUMB[4][60] ), 
        .CO(\CARRYB[5][59] ), .S(\SUMB[5][59] ) );
  FA1A S2_5_58 ( .A(\ab[5][58] ), .B(\CARRYB[4][58] ), .CI(\SUMB[4][59] ), 
        .CO(\CARRYB[5][58] ), .S(\SUMB[5][58] ) );
  FA1A S2_5_56 ( .A(\ab[5][56] ), .B(\CARRYB[4][56] ), .CI(\SUMB[4][57] ), 
        .CO(\CARRYB[5][56] ), .S(\SUMB[5][56] ) );
  FA1A S2_5_54 ( .A(\ab[5][54] ), .B(\CARRYB[4][54] ), .CI(\SUMB[4][55] ), 
        .CO(\CARRYB[5][54] ), .S(\SUMB[5][54] ) );
  FA1A S2_5_53 ( .A(\ab[5][53] ), .B(\CARRYB[4][53] ), .CI(\SUMB[4][54] ), 
        .CO(\CARRYB[5][53] ), .S(\SUMB[5][53] ) );
  FA1A S2_4_59 ( .A(\ab[4][59] ), .B(\CARRYB[3][59] ), .CI(\SUMB[3][60] ), 
        .CO(\CARRYB[4][59] ), .S(\SUMB[4][59] ) );
  FA1A S2_4_58 ( .A(\ab[4][58] ), .B(\CARRYB[3][58] ), .CI(\SUMB[3][59] ), 
        .CO(\CARRYB[4][58] ), .S(\SUMB[4][58] ) );
  FA1A S2_4_56 ( .A(\ab[4][56] ), .B(\CARRYB[3][56] ), .CI(\SUMB[3][57] ), 
        .CO(\CARRYB[4][56] ), .S(\SUMB[4][56] ) );
  FA1A S2_4_54 ( .A(\ab[4][54] ), .B(\CARRYB[3][54] ), .CI(\SUMB[3][55] ), 
        .CO(\CARRYB[4][54] ), .S(\SUMB[4][54] ) );
  FA1A S2_4_53 ( .A(\ab[4][53] ), .B(\CARRYB[3][53] ), .CI(\SUMB[3][54] ), 
        .CO(\CARRYB[4][53] ), .S(\SUMB[4][53] ) );
  FA1A S2_3_59 ( .A(\ab[3][59] ), .B(\CARRYB[2][59] ), .CI(\SUMB[2][60] ), 
        .CO(\CARRYB[3][59] ), .S(\SUMB[3][59] ) );
  FA1A S2_3_58 ( .A(\ab[3][58] ), .B(\CARRYB[2][58] ), .CI(\SUMB[2][59] ), 
        .CO(\CARRYB[3][58] ), .S(\SUMB[3][58] ) );
  FA1A S2_3_56 ( .A(\ab[3][56] ), .B(\CARRYB[2][56] ), .CI(\SUMB[2][57] ), 
        .CO(\CARRYB[3][56] ), .S(\SUMB[3][56] ) );
  FA1A S2_3_54 ( .A(\ab[3][54] ), .B(\CARRYB[2][54] ), .CI(\SUMB[2][55] ), 
        .CO(\CARRYB[3][54] ), .S(\SUMB[3][54] ) );
  FA1A S2_3_53 ( .A(\ab[3][53] ), .B(\CARRYB[2][53] ), .CI(\SUMB[2][54] ), 
        .CO(\CARRYB[3][53] ), .S(\SUMB[3][53] ) );
  FA1A S2_2_59 ( .A(\ab[2][59] ), .B(\CARRYB[1][59] ), .CI(\SUMB[1][60] ), 
        .CO(\CARRYB[2][59] ), .S(\SUMB[2][59] ) );
  FA1A S2_2_58 ( .A(\ab[2][58] ), .B(\CARRYB[1][58] ), .CI(\SUMB[1][59] ), 
        .CO(\CARRYB[2][58] ), .S(\SUMB[2][58] ) );
  FA1A S2_2_56 ( .A(\ab[2][56] ), .B(\CARRYB[1][56] ), .CI(\SUMB[1][57] ), 
        .CO(\CARRYB[2][56] ), .S(\SUMB[2][56] ) );
  FA1A S2_2_54 ( .A(\ab[2][54] ), .B(\CARRYB[1][54] ), .CI(\SUMB[1][55] ), 
        .CO(\CARRYB[2][54] ), .S(\SUMB[2][54] ) );
  FA1A S2_2_53 ( .A(\ab[2][53] ), .B(\CARRYB[1][53] ), .CI(\SUMB[1][54] ), 
        .CO(\CARRYB[2][53] ), .S(\SUMB[2][53] ) );
  FA1A S2_14_52 ( .A(\ab[14][52] ), .B(\CARRYB[13][52] ), .CI(\SUMB[13][53] ), 
        .CO(\CARRYB[14][52] ), .S(\SUMB[14][52] ) );
  FA1A S2_14_44 ( .A(\ab[14][44] ), .B(\CARRYB[13][44] ), .CI(\SUMB[13][45] ), 
        .CO(\CARRYB[14][44] ), .S(\SUMB[14][44] ) );
  FA1A S2_14_43 ( .A(\ab[14][43] ), .B(\CARRYB[13][43] ), .CI(\SUMB[13][44] ), 
        .CO(\CARRYB[14][43] ), .S(\SUMB[14][43] ) );
  FA1A S2_14_42 ( .A(\ab[14][42] ), .B(\CARRYB[13][42] ), .CI(\SUMB[13][43] ), 
        .CO(\CARRYB[14][42] ), .S(\SUMB[14][42] ) );
  FA1A S2_14_41 ( .A(\ab[14][41] ), .B(\CARRYB[13][41] ), .CI(\SUMB[13][42] ), 
        .CO(\CARRYB[14][41] ), .S(\SUMB[14][41] ) );
  FA1A S2_13_52 ( .A(\ab[13][52] ), .B(\CARRYB[12][52] ), .CI(\SUMB[12][53] ), 
        .CO(\CARRYB[13][52] ), .S(\SUMB[13][52] ) );
  FA1A S2_13_44 ( .A(\ab[13][44] ), .B(\CARRYB[12][44] ), .CI(\SUMB[12][45] ), 
        .CO(\CARRYB[13][44] ), .S(\SUMB[13][44] ) );
  FA1A S2_13_43 ( .A(\ab[13][43] ), .B(\CARRYB[12][43] ), .CI(\SUMB[12][44] ), 
        .CO(\CARRYB[13][43] ), .S(\SUMB[13][43] ) );
  FA1A S2_13_42 ( .A(\ab[13][42] ), .B(\CARRYB[12][42] ), .CI(\SUMB[12][43] ), 
        .CO(\CARRYB[13][42] ), .S(\SUMB[13][42] ) );
  FA1A S2_14_39 ( .A(\ab[14][39] ), .B(\CARRYB[13][39] ), .CI(\SUMB[13][40] ), 
        .CO(\CARRYB[14][39] ), .S(\SUMB[14][39] ) );
  FA1A S2_14_40 ( .A(\ab[14][40] ), .B(\CARRYB[13][40] ), .CI(\SUMB[13][41] ), 
        .CO(\CARRYB[14][40] ), .S(\SUMB[14][40] ) );
  FA1A S2_12_52 ( .A(\ab[12][52] ), .B(\CARRYB[11][52] ), .CI(\SUMB[11][53] ), 
        .CO(\CARRYB[12][52] ), .S(\SUMB[12][52] ) );
  FA1A S2_12_44 ( .A(\ab[12][44] ), .B(\CARRYB[11][44] ), .CI(\SUMB[11][45] ), 
        .CO(\CARRYB[12][44] ), .S(\SUMB[12][44] ) );
  FA1A S2_12_43 ( .A(\ab[12][43] ), .B(\CARRYB[11][43] ), .CI(\SUMB[11][44] ), 
        .CO(\CARRYB[12][43] ), .S(\SUMB[12][43] ) );
  FA1A S2_13_40 ( .A(\ab[13][40] ), .B(\CARRYB[12][40] ), .CI(\SUMB[12][41] ), 
        .CO(\CARRYB[13][40] ), .S(\SUMB[13][40] ) );
  FA1A S2_13_41 ( .A(\ab[13][41] ), .B(\CARRYB[12][41] ), .CI(\SUMB[12][42] ), 
        .CO(\CARRYB[13][41] ), .S(\SUMB[13][41] ) );
  FA1A S2_11_52 ( .A(\ab[11][52] ), .B(\CARRYB[10][52] ), .CI(\SUMB[10][53] ), 
        .CO(\CARRYB[11][52] ), .S(\SUMB[11][52] ) );
  FA1A S2_11_44 ( .A(\ab[11][44] ), .B(\CARRYB[10][44] ), .CI(\SUMB[10][45] ), 
        .CO(\CARRYB[11][44] ), .S(\SUMB[11][44] ) );
  FA1A S2_12_41 ( .A(\ab[12][41] ), .B(\CARRYB[11][41] ), .CI(\SUMB[11][42] ), 
        .CO(\CARRYB[12][41] ), .S(\SUMB[12][41] ) );
  FA1A S2_12_42 ( .A(\ab[12][42] ), .B(\CARRYB[11][42] ), .CI(\SUMB[11][43] ), 
        .CO(\CARRYB[12][42] ), .S(\SUMB[12][42] ) );
  FA1A S2_13_39 ( .A(\ab[13][39] ), .B(\CARRYB[12][39] ), .CI(\SUMB[12][40] ), 
        .CO(\CARRYB[13][39] ), .S(\SUMB[13][39] ) );
  FA1A S2_10_52 ( .A(\ab[10][52] ), .B(\CARRYB[9][52] ), .CI(\SUMB[9][53] ), 
        .CO(\CARRYB[10][52] ), .S(\SUMB[10][52] ) );
  FA1A S2_11_42 ( .A(\ab[11][42] ), .B(\CARRYB[10][42] ), .CI(\SUMB[10][43] ), 
        .CO(\CARRYB[11][42] ), .S(\SUMB[11][42] ) );
  FA1A S2_11_43 ( .A(\ab[11][43] ), .B(\CARRYB[10][43] ), .CI(\SUMB[10][44] ), 
        .CO(\CARRYB[11][43] ), .S(\SUMB[11][43] ) );
  FA1A S2_12_40 ( .A(\ab[12][40] ), .B(\CARRYB[11][40] ), .CI(\SUMB[11][41] ), 
        .CO(\CARRYB[12][40] ), .S(\SUMB[12][40] ) );
  FA1A S2_12_39 ( .A(\ab[12][39] ), .B(\CARRYB[11][39] ), .CI(\SUMB[11][40] ), 
        .CO(\CARRYB[12][39] ), .S(\SUMB[12][39] ) );
  FA1A S2_9_52 ( .A(\ab[9][52] ), .B(\CARRYB[8][52] ), .CI(\SUMB[8][53] ), 
        .CO(\CARRYB[9][52] ), .S(\SUMB[9][52] ) );
  FA1A S2_10_43 ( .A(\ab[10][43] ), .B(\CARRYB[9][43] ), .CI(\SUMB[9][44] ), 
        .CO(\CARRYB[10][43] ), .S(\SUMB[10][43] ) );
  FA1A S2_10_44 ( .A(\ab[10][44] ), .B(\CARRYB[9][44] ), .CI(\SUMB[9][45] ), 
        .CO(\CARRYB[10][44] ), .S(\SUMB[10][44] ) );
  FA1A S2_11_41 ( .A(\ab[11][41] ), .B(\CARRYB[10][41] ), .CI(\SUMB[10][42] ), 
        .CO(\CARRYB[11][41] ), .S(\SUMB[11][41] ) );
  FA1A S2_11_40 ( .A(\ab[11][40] ), .B(\CARRYB[10][40] ), .CI(\SUMB[10][41] ), 
        .CO(\CARRYB[11][40] ), .S(\SUMB[11][40] ) );
  FA1A S2_11_39 ( .A(\ab[11][39] ), .B(\CARRYB[10][39] ), .CI(\SUMB[10][40] ), 
        .CO(\CARRYB[11][39] ), .S(\SUMB[11][39] ) );
  FA1A S2_8_52 ( .A(\ab[8][52] ), .B(\CARRYB[7][52] ), .CI(\SUMB[7][53] ), 
        .CO(\CARRYB[8][52] ), .S(\SUMB[8][52] ) );
  FA1A S2_9_44 ( .A(\ab[9][44] ), .B(\CARRYB[8][44] ), .CI(\SUMB[8][45] ), 
        .CO(\CARRYB[9][44] ), .S(\SUMB[9][44] ) );
  FA1A S2_10_42 ( .A(\ab[10][42] ), .B(\CARRYB[9][42] ), .CI(\SUMB[9][43] ), 
        .CO(\CARRYB[10][42] ), .S(\SUMB[10][42] ) );
  FA1A S2_10_41 ( .A(\ab[10][41] ), .B(\CARRYB[9][41] ), .CI(\SUMB[9][42] ), 
        .CO(\CARRYB[10][41] ), .S(\SUMB[10][41] ) );
  FA1A S2_10_40 ( .A(\ab[10][40] ), .B(\CARRYB[9][40] ), .CI(\SUMB[9][41] ), 
        .CO(\CARRYB[10][40] ), .S(\SUMB[10][40] ) );
  FA1A S2_10_39 ( .A(\ab[10][39] ), .B(\CARRYB[9][39] ), .CI(\SUMB[9][40] ), 
        .CO(\CARRYB[10][39] ), .S(\SUMB[10][39] ) );
  FA1A S2_7_52 ( .A(\ab[7][52] ), .B(\CARRYB[6][52] ), .CI(\SUMB[6][53] ), 
        .CO(\CARRYB[7][52] ), .S(\SUMB[7][52] ) );
  FA1A S2_9_43 ( .A(\ab[9][43] ), .B(\CARRYB[8][43] ), .CI(\SUMB[8][44] ), 
        .CO(\CARRYB[9][43] ), .S(\SUMB[9][43] ) );
  FA1A S2_9_42 ( .A(\ab[9][42] ), .B(\CARRYB[8][42] ), .CI(\SUMB[8][43] ), 
        .CO(\CARRYB[9][42] ), .S(\SUMB[9][42] ) );
  FA1A S2_9_41 ( .A(\ab[9][41] ), .B(\CARRYB[8][41] ), .CI(\SUMB[8][42] ), 
        .CO(\CARRYB[9][41] ), .S(\SUMB[9][41] ) );
  FA1A S2_9_40 ( .A(\ab[9][40] ), .B(\CARRYB[8][40] ), .CI(\SUMB[8][41] ), 
        .CO(\CARRYB[9][40] ), .S(\SUMB[9][40] ) );
  FA1A S2_9_39 ( .A(\ab[9][39] ), .B(\CARRYB[8][39] ), .CI(\SUMB[8][40] ), 
        .CO(\CARRYB[9][39] ), .S(\SUMB[9][39] ) );
  FA1A S2_6_52 ( .A(\ab[6][52] ), .B(\CARRYB[5][52] ), .CI(\SUMB[5][53] ), 
        .CO(\CARRYB[6][52] ), .S(\SUMB[6][52] ) );
  FA1A S2_8_44 ( .A(\ab[8][44] ), .B(\CARRYB[7][44] ), .CI(\SUMB[7][45] ), 
        .CO(\CARRYB[8][44] ), .S(\SUMB[8][44] ) );
  FA1A S2_8_43 ( .A(\ab[8][43] ), .B(\CARRYB[7][43] ), .CI(\SUMB[7][44] ), 
        .CO(\CARRYB[8][43] ), .S(\SUMB[8][43] ) );
  FA1A S2_8_42 ( .A(\ab[8][42] ), .B(\CARRYB[7][42] ), .CI(\SUMB[7][43] ), 
        .CO(\CARRYB[8][42] ), .S(\SUMB[8][42] ) );
  FA1A S2_8_41 ( .A(\ab[8][41] ), .B(\CARRYB[7][41] ), .CI(\SUMB[7][42] ), 
        .CO(\CARRYB[8][41] ), .S(\SUMB[8][41] ) );
  FA1A S2_8_40 ( .A(\ab[8][40] ), .B(\CARRYB[7][40] ), .CI(\SUMB[7][41] ), 
        .CO(\CARRYB[8][40] ), .S(\SUMB[8][40] ) );
  FA1A S2_8_39 ( .A(\ab[8][39] ), .B(\CARRYB[7][39] ), .CI(\SUMB[7][40] ), 
        .CO(\CARRYB[8][39] ), .S(\SUMB[8][39] ) );
  FA1A S2_5_52 ( .A(\ab[5][52] ), .B(\CARRYB[4][52] ), .CI(\SUMB[4][53] ), 
        .CO(\CARRYB[5][52] ), .S(\SUMB[5][52] ) );
  FA1A S2_7_44 ( .A(\ab[7][44] ), .B(\CARRYB[6][44] ), .CI(\SUMB[6][45] ), 
        .CO(\CARRYB[7][44] ), .S(\SUMB[7][44] ) );
  FA1A S2_7_43 ( .A(\ab[7][43] ), .B(\CARRYB[6][43] ), .CI(\SUMB[6][44] ), 
        .CO(\CARRYB[7][43] ), .S(\SUMB[7][43] ) );
  FA1A S2_7_42 ( .A(\ab[7][42] ), .B(\CARRYB[6][42] ), .CI(\SUMB[6][43] ), 
        .CO(\CARRYB[7][42] ), .S(\SUMB[7][42] ) );
  FA1A S2_7_41 ( .A(\ab[7][41] ), .B(\CARRYB[6][41] ), .CI(\SUMB[6][42] ), 
        .CO(\CARRYB[7][41] ), .S(\SUMB[7][41] ) );
  FA1A S2_7_40 ( .A(\ab[7][40] ), .B(\CARRYB[6][40] ), .CI(\SUMB[6][41] ), 
        .CO(\CARRYB[7][40] ), .S(\SUMB[7][40] ) );
  FA1A S2_7_39 ( .A(\ab[7][39] ), .B(\CARRYB[6][39] ), .CI(\SUMB[6][40] ), 
        .CO(\CARRYB[7][39] ), .S(\SUMB[7][39] ) );
  FA1A S2_4_52 ( .A(\ab[4][52] ), .B(\CARRYB[3][52] ), .CI(\SUMB[3][53] ), 
        .CO(\CARRYB[4][52] ), .S(\SUMB[4][52] ) );
  FA1A S2_6_44 ( .A(\ab[6][44] ), .B(\CARRYB[5][44] ), .CI(\SUMB[5][45] ), 
        .CO(\CARRYB[6][44] ), .S(\SUMB[6][44] ) );
  FA1A S2_6_43 ( .A(\ab[6][43] ), .B(\CARRYB[5][43] ), .CI(\SUMB[5][44] ), 
        .CO(\CARRYB[6][43] ), .S(\SUMB[6][43] ) );
  FA1A S2_6_42 ( .A(\ab[6][42] ), .B(\CARRYB[5][42] ), .CI(\SUMB[5][43] ), 
        .CO(\CARRYB[6][42] ), .S(\SUMB[6][42] ) );
  FA1A S2_6_41 ( .A(\ab[6][41] ), .B(\CARRYB[5][41] ), .CI(\SUMB[5][42] ), 
        .CO(\CARRYB[6][41] ), .S(\SUMB[6][41] ) );
  FA1A S2_6_40 ( .A(\ab[6][40] ), .B(\CARRYB[5][40] ), .CI(\SUMB[5][41] ), 
        .CO(\CARRYB[6][40] ), .S(\SUMB[6][40] ) );
  FA1A S2_6_39 ( .A(\ab[6][39] ), .B(\CARRYB[5][39] ), .CI(\SUMB[5][40] ), 
        .CO(\CARRYB[6][39] ), .S(\SUMB[6][39] ) );
  FA1A S2_3_52 ( .A(\ab[3][52] ), .B(\CARRYB[2][52] ), .CI(\SUMB[2][53] ), 
        .CO(\CARRYB[3][52] ), .S(\SUMB[3][52] ) );
  FA1A S2_5_44 ( .A(\ab[5][44] ), .B(\CARRYB[4][44] ), .CI(\SUMB[4][45] ), 
        .CO(\CARRYB[5][44] ), .S(\SUMB[5][44] ) );
  FA1A S2_5_43 ( .A(\ab[5][43] ), .B(\CARRYB[4][43] ), .CI(\SUMB[4][44] ), 
        .CO(\CARRYB[5][43] ), .S(\SUMB[5][43] ) );
  FA1A S2_5_42 ( .A(\ab[5][42] ), .B(\CARRYB[4][42] ), .CI(\SUMB[4][43] ), 
        .CO(\CARRYB[5][42] ), .S(\SUMB[5][42] ) );
  FA1A S2_5_41 ( .A(\ab[5][41] ), .B(\CARRYB[4][41] ), .CI(\SUMB[4][42] ), 
        .CO(\CARRYB[5][41] ), .S(\SUMB[5][41] ) );
  FA1A S2_5_40 ( .A(\ab[5][40] ), .B(\CARRYB[4][40] ), .CI(\SUMB[4][41] ), 
        .CO(\CARRYB[5][40] ), .S(\SUMB[5][40] ) );
  FA1A S2_5_39 ( .A(\ab[5][39] ), .B(\CARRYB[4][39] ), .CI(\SUMB[4][40] ), 
        .CO(\CARRYB[5][39] ), .S(\SUMB[5][39] ) );
  FA1A S2_4_44 ( .A(\ab[4][44] ), .B(\CARRYB[3][44] ), .CI(\SUMB[3][45] ), 
        .CO(\CARRYB[4][44] ), .S(\SUMB[4][44] ) );
  FA1A S2_4_43 ( .A(\ab[4][43] ), .B(\CARRYB[3][43] ), .CI(\SUMB[3][44] ), 
        .CO(\CARRYB[4][43] ), .S(\SUMB[4][43] ) );
  FA1A S2_4_42 ( .A(\ab[4][42] ), .B(\CARRYB[3][42] ), .CI(\SUMB[3][43] ), 
        .CO(\CARRYB[4][42] ), .S(\SUMB[4][42] ) );
  FA1A S2_4_41 ( .A(\ab[4][41] ), .B(\CARRYB[3][41] ), .CI(\SUMB[3][42] ), 
        .CO(\CARRYB[4][41] ), .S(\SUMB[4][41] ) );
  FA1A S2_4_40 ( .A(\ab[4][40] ), .B(\CARRYB[3][40] ), .CI(\SUMB[3][41] ), 
        .CO(\CARRYB[4][40] ), .S(\SUMB[4][40] ) );
  FA1A S2_4_39 ( .A(\ab[4][39] ), .B(\CARRYB[3][39] ), .CI(\SUMB[3][40] ), 
        .CO(\CARRYB[4][39] ), .S(\SUMB[4][39] ) );
  FA1A S2_2_52 ( .A(\ab[2][52] ), .B(\CARRYB[1][52] ), .CI(\SUMB[1][53] ), 
        .CO(\CARRYB[2][52] ), .S(\SUMB[2][52] ) );
  FA1A S2_3_44 ( .A(\ab[3][44] ), .B(\CARRYB[2][44] ), .CI(\SUMB[2][45] ), 
        .CO(\CARRYB[3][44] ), .S(\SUMB[3][44] ) );
  FA1A S2_3_43 ( .A(\ab[3][43] ), .B(\CARRYB[2][43] ), .CI(\SUMB[2][44] ), 
        .CO(\CARRYB[3][43] ), .S(\SUMB[3][43] ) );
  FA1A S2_3_42 ( .A(\ab[3][42] ), .B(\CARRYB[2][42] ), .CI(\SUMB[2][43] ), 
        .CO(\CARRYB[3][42] ), .S(\SUMB[3][42] ) );
  FA1A S2_3_41 ( .A(\ab[3][41] ), .B(\CARRYB[2][41] ), .CI(\SUMB[2][42] ), 
        .CO(\CARRYB[3][41] ), .S(\SUMB[3][41] ) );
  FA1A S2_3_40 ( .A(\ab[3][40] ), .B(\CARRYB[2][40] ), .CI(\SUMB[2][41] ), 
        .CO(\CARRYB[3][40] ), .S(\SUMB[3][40] ) );
  FA1A S2_3_39 ( .A(\ab[3][39] ), .B(\CARRYB[2][39] ), .CI(\SUMB[2][40] ), 
        .CO(\CARRYB[3][39] ), .S(\SUMB[3][39] ) );
  FA1A S2_2_44 ( .A(\ab[2][44] ), .B(\CARRYB[1][44] ), .CI(\SUMB[1][45] ), 
        .CO(\CARRYB[2][44] ), .S(\SUMB[2][44] ) );
  FA1A S2_2_43 ( .A(\ab[2][43] ), .B(\CARRYB[1][43] ), .CI(\SUMB[1][44] ), 
        .CO(\CARRYB[2][43] ), .S(\SUMB[2][43] ) );
  FA1A S2_2_42 ( .A(\ab[2][42] ), .B(\CARRYB[1][42] ), .CI(\SUMB[1][43] ), 
        .CO(\CARRYB[2][42] ), .S(\SUMB[2][42] ) );
  FA1A S2_2_41 ( .A(\ab[2][41] ), .B(\CARRYB[1][41] ), .CI(\SUMB[1][42] ), 
        .CO(\CARRYB[2][41] ), .S(\SUMB[2][41] ) );
  FA1A S2_2_40 ( .A(\ab[2][40] ), .B(\CARRYB[1][40] ), .CI(\SUMB[1][41] ), 
        .CO(\CARRYB[2][40] ), .S(\SUMB[2][40] ) );
  FA1A S2_2_39 ( .A(\ab[2][39] ), .B(\CARRYB[1][39] ), .CI(\SUMB[1][40] ), 
        .CO(\CARRYB[2][39] ), .S(\SUMB[2][39] ) );
  FA1A S2_14_51 ( .A(\ab[14][51] ), .B(\CARRYB[13][51] ), .CI(\SUMB[13][52] ), 
        .CO(\CARRYB[14][51] ), .S(\SUMB[14][51] ) );
  FA1A S2_14_50 ( .A(\ab[14][50] ), .B(\CARRYB[13][50] ), .CI(\SUMB[13][51] ), 
        .CO(\CARRYB[14][50] ), .S(\SUMB[14][50] ) );
  FA1A S2_14_49 ( .A(\ab[14][49] ), .B(\CARRYB[13][49] ), .CI(\SUMB[13][50] ), 
        .CO(\CARRYB[14][49] ), .S(\SUMB[14][49] ) );
  FA1A S2_14_48 ( .A(\ab[14][48] ), .B(\CARRYB[13][48] ), .CI(\SUMB[13][49] ), 
        .CO(\CARRYB[14][48] ), .S(\SUMB[14][48] ) );
  FA1A S2_14_47 ( .A(\ab[14][47] ), .B(\CARRYB[13][47] ), .CI(\SUMB[13][48] ), 
        .CO(\CARRYB[14][47] ), .S(\SUMB[14][47] ) );
  FA1A S2_14_46 ( .A(\ab[14][46] ), .B(\CARRYB[13][46] ), .CI(\SUMB[13][47] ), 
        .CO(\CARRYB[14][46] ), .S(\SUMB[14][46] ) );
  FA1A S2_14_45 ( .A(\ab[14][45] ), .B(\CARRYB[13][45] ), .CI(\SUMB[13][46] ), 
        .CO(\CARRYB[14][45] ), .S(\SUMB[14][45] ) );
  FA1A S2_13_51 ( .A(\ab[13][51] ), .B(\CARRYB[12][51] ), .CI(\SUMB[12][52] ), 
        .CO(\CARRYB[13][51] ), .S(\SUMB[13][51] ) );
  FA1A S2_13_50 ( .A(\ab[13][50] ), .B(\CARRYB[12][50] ), .CI(\SUMB[12][51] ), 
        .CO(\CARRYB[13][50] ), .S(\SUMB[13][50] ) );
  FA1A S2_13_49 ( .A(\ab[13][49] ), .B(\CARRYB[12][49] ), .CI(\SUMB[12][50] ), 
        .CO(\CARRYB[13][49] ), .S(\SUMB[13][49] ) );
  FA1A S2_13_48 ( .A(\ab[13][48] ), .B(\CARRYB[12][48] ), .CI(\SUMB[12][49] ), 
        .CO(\CARRYB[13][48] ), .S(\SUMB[13][48] ) );
  FA1A S2_13_47 ( .A(\ab[13][47] ), .B(\CARRYB[12][47] ), .CI(\SUMB[12][48] ), 
        .CO(\CARRYB[13][47] ), .S(\SUMB[13][47] ) );
  FA1A S2_13_46 ( .A(\ab[13][46] ), .B(\CARRYB[12][46] ), .CI(\SUMB[12][47] ), 
        .CO(\CARRYB[13][46] ), .S(\SUMB[13][46] ) );
  FA1A S2_13_45 ( .A(\ab[13][45] ), .B(\CARRYB[12][45] ), .CI(\SUMB[12][46] ), 
        .CO(\CARRYB[13][45] ), .S(\SUMB[13][45] ) );
  FA1A S2_12_51 ( .A(\ab[12][51] ), .B(\CARRYB[11][51] ), .CI(\SUMB[11][52] ), 
        .CO(\CARRYB[12][51] ), .S(\SUMB[12][51] ) );
  FA1A S2_12_50 ( .A(\ab[12][50] ), .B(\CARRYB[11][50] ), .CI(\SUMB[11][51] ), 
        .CO(\CARRYB[12][50] ), .S(\SUMB[12][50] ) );
  FA1A S2_12_49 ( .A(\ab[12][49] ), .B(\CARRYB[11][49] ), .CI(\SUMB[11][50] ), 
        .CO(\CARRYB[12][49] ), .S(\SUMB[12][49] ) );
  FA1A S2_12_48 ( .A(\ab[12][48] ), .B(\CARRYB[11][48] ), .CI(\SUMB[11][49] ), 
        .CO(\CARRYB[12][48] ), .S(\SUMB[12][48] ) );
  FA1A S2_12_47 ( .A(\ab[12][47] ), .B(\CARRYB[11][47] ), .CI(\SUMB[11][48] ), 
        .CO(\CARRYB[12][47] ), .S(\SUMB[12][47] ) );
  FA1A S2_12_46 ( .A(\ab[12][46] ), .B(\CARRYB[11][46] ), .CI(\SUMB[11][47] ), 
        .CO(\CARRYB[12][46] ), .S(\SUMB[12][46] ) );
  FA1A S2_12_45 ( .A(\ab[12][45] ), .B(\CARRYB[11][45] ), .CI(\SUMB[11][46] ), 
        .CO(\CARRYB[12][45] ), .S(\SUMB[12][45] ) );
  FA1A S2_11_51 ( .A(\ab[11][51] ), .B(\CARRYB[10][51] ), .CI(\SUMB[10][52] ), 
        .CO(\CARRYB[11][51] ), .S(\SUMB[11][51] ) );
  FA1A S2_11_50 ( .A(\ab[11][50] ), .B(\CARRYB[10][50] ), .CI(\SUMB[10][51] ), 
        .CO(\CARRYB[11][50] ), .S(\SUMB[11][50] ) );
  FA1A S2_11_49 ( .A(\ab[11][49] ), .B(\CARRYB[10][49] ), .CI(\SUMB[10][50] ), 
        .CO(\CARRYB[11][49] ), .S(\SUMB[11][49] ) );
  FA1A S2_11_48 ( .A(\ab[11][48] ), .B(\CARRYB[10][48] ), .CI(\SUMB[10][49] ), 
        .CO(\CARRYB[11][48] ), .S(\SUMB[11][48] ) );
  FA1A S2_11_47 ( .A(\ab[11][47] ), .B(\CARRYB[10][47] ), .CI(\SUMB[10][48] ), 
        .CO(\CARRYB[11][47] ), .S(\SUMB[11][47] ) );
  FA1A S2_11_46 ( .A(\ab[11][46] ), .B(\CARRYB[10][46] ), .CI(\SUMB[10][47] ), 
        .CO(\CARRYB[11][46] ), .S(\SUMB[11][46] ) );
  FA1A S2_11_45 ( .A(\ab[11][45] ), .B(\CARRYB[10][45] ), .CI(\SUMB[10][46] ), 
        .CO(\CARRYB[11][45] ), .S(\SUMB[11][45] ) );
  FA1A S2_10_51 ( .A(\ab[10][51] ), .B(\CARRYB[9][51] ), .CI(\SUMB[9][52] ), 
        .CO(\CARRYB[10][51] ), .S(\SUMB[10][51] ) );
  FA1A S2_10_50 ( .A(\ab[10][50] ), .B(\CARRYB[9][50] ), .CI(\SUMB[9][51] ), 
        .CO(\CARRYB[10][50] ), .S(\SUMB[10][50] ) );
  FA1A S2_10_49 ( .A(\ab[10][49] ), .B(\CARRYB[9][49] ), .CI(\SUMB[9][50] ), 
        .CO(\CARRYB[10][49] ), .S(\SUMB[10][49] ) );
  FA1A S2_10_48 ( .A(\ab[10][48] ), .B(\CARRYB[9][48] ), .CI(\SUMB[9][49] ), 
        .CO(\CARRYB[10][48] ), .S(\SUMB[10][48] ) );
  FA1A S2_10_47 ( .A(\ab[10][47] ), .B(\CARRYB[9][47] ), .CI(\SUMB[9][48] ), 
        .CO(\CARRYB[10][47] ), .S(\SUMB[10][47] ) );
  FA1A S2_10_46 ( .A(\ab[10][46] ), .B(\CARRYB[9][46] ), .CI(\SUMB[9][47] ), 
        .CO(\CARRYB[10][46] ), .S(\SUMB[10][46] ) );
  FA1A S2_10_45 ( .A(\ab[10][45] ), .B(\CARRYB[9][45] ), .CI(\SUMB[9][46] ), 
        .CO(\CARRYB[10][45] ), .S(\SUMB[10][45] ) );
  FA1A S2_9_51 ( .A(\ab[9][51] ), .B(\CARRYB[8][51] ), .CI(\SUMB[8][52] ), 
        .CO(\CARRYB[9][51] ), .S(\SUMB[9][51] ) );
  FA1A S2_9_50 ( .A(\ab[9][50] ), .B(\CARRYB[8][50] ), .CI(\SUMB[8][51] ), 
        .CO(\CARRYB[9][50] ), .S(\SUMB[9][50] ) );
  FA1A S2_9_49 ( .A(\ab[9][49] ), .B(\CARRYB[8][49] ), .CI(\SUMB[8][50] ), 
        .CO(\CARRYB[9][49] ), .S(\SUMB[9][49] ) );
  FA1A S2_9_48 ( .A(\ab[9][48] ), .B(\CARRYB[8][48] ), .CI(\SUMB[8][49] ), 
        .CO(\CARRYB[9][48] ), .S(\SUMB[9][48] ) );
  FA1A S2_9_47 ( .A(\ab[9][47] ), .B(\CARRYB[8][47] ), .CI(\SUMB[8][48] ), 
        .CO(\CARRYB[9][47] ), .S(\SUMB[9][47] ) );
  FA1A S2_9_46 ( .A(\ab[9][46] ), .B(\CARRYB[8][46] ), .CI(\SUMB[8][47] ), 
        .CO(\CARRYB[9][46] ), .S(\SUMB[9][46] ) );
  FA1A S2_8_51 ( .A(\ab[8][51] ), .B(\CARRYB[7][51] ), .CI(\SUMB[7][52] ), 
        .CO(\CARRYB[8][51] ), .S(\SUMB[8][51] ) );
  FA1A S2_8_50 ( .A(\ab[8][50] ), .B(\CARRYB[7][50] ), .CI(\SUMB[7][51] ), 
        .CO(\CARRYB[8][50] ), .S(\SUMB[8][50] ) );
  FA1A S2_8_49 ( .A(\ab[8][49] ), .B(\CARRYB[7][49] ), .CI(\SUMB[7][50] ), 
        .CO(\CARRYB[8][49] ), .S(\SUMB[8][49] ) );
  FA1A S2_8_48 ( .A(\ab[8][48] ), .B(\CARRYB[7][48] ), .CI(\SUMB[7][49] ), 
        .CO(\CARRYB[8][48] ), .S(\SUMB[8][48] ) );
  FA1A S2_8_47 ( .A(\ab[8][47] ), .B(\CARRYB[7][47] ), .CI(\SUMB[7][48] ), 
        .CO(\CARRYB[8][47] ), .S(\SUMB[8][47] ) );
  FA1A S2_9_45 ( .A(\ab[9][45] ), .B(\CARRYB[8][45] ), .CI(\SUMB[8][46] ), 
        .CO(\CARRYB[9][45] ), .S(\SUMB[9][45] ) );
  FA1A S2_7_51 ( .A(\ab[7][51] ), .B(\CARRYB[6][51] ), .CI(\SUMB[6][52] ), 
        .CO(\CARRYB[7][51] ), .S(\SUMB[7][51] ) );
  FA1A S2_7_50 ( .A(\ab[7][50] ), .B(\CARRYB[6][50] ), .CI(\SUMB[6][51] ), 
        .CO(\CARRYB[7][50] ), .S(\SUMB[7][50] ) );
  FA1A S2_7_49 ( .A(\ab[7][49] ), .B(\CARRYB[6][49] ), .CI(\SUMB[6][50] ), 
        .CO(\CARRYB[7][49] ), .S(\SUMB[7][49] ) );
  FA1A S2_7_48 ( .A(\ab[7][48] ), .B(\CARRYB[6][48] ), .CI(\SUMB[6][49] ), 
        .CO(\CARRYB[7][48] ), .S(\SUMB[7][48] ) );
  FA1A S2_8_45 ( .A(\ab[8][45] ), .B(\CARRYB[7][45] ), .CI(\SUMB[7][46] ), 
        .CO(\CARRYB[8][45] ), .S(\SUMB[8][45] ) );
  FA1A S2_8_46 ( .A(\ab[8][46] ), .B(\CARRYB[7][46] ), .CI(\SUMB[7][47] ), 
        .CO(\CARRYB[8][46] ), .S(\SUMB[8][46] ) );
  FA1A S2_6_51 ( .A(\ab[6][51] ), .B(\CARRYB[5][51] ), .CI(\SUMB[5][52] ), 
        .CO(\CARRYB[6][51] ), .S(\SUMB[6][51] ) );
  FA1A S2_6_50 ( .A(\ab[6][50] ), .B(\CARRYB[5][50] ), .CI(\SUMB[5][51] ), 
        .CO(\CARRYB[6][50] ), .S(\SUMB[6][50] ) );
  FA1A S2_6_49 ( .A(\ab[6][49] ), .B(\CARRYB[5][49] ), .CI(\SUMB[5][50] ), 
        .CO(\CARRYB[6][49] ), .S(\SUMB[6][49] ) );
  FA1A S2_7_46 ( .A(\ab[7][46] ), .B(\CARRYB[6][46] ), .CI(\SUMB[6][47] ), 
        .CO(\CARRYB[7][46] ), .S(\SUMB[7][46] ) );
  FA1A S2_7_47 ( .A(\ab[7][47] ), .B(\CARRYB[6][47] ), .CI(\SUMB[6][48] ), 
        .CO(\CARRYB[7][47] ), .S(\SUMB[7][47] ) );
  FA1A S2_5_51 ( .A(\ab[5][51] ), .B(\CARRYB[4][51] ), .CI(\SUMB[4][52] ), 
        .CO(\CARRYB[5][51] ), .S(\SUMB[5][51] ) );
  FA1A S2_5_50 ( .A(\ab[5][50] ), .B(\CARRYB[4][50] ), .CI(\SUMB[4][51] ), 
        .CO(\CARRYB[5][50] ), .S(\SUMB[5][50] ) );
  FA1A S2_6_47 ( .A(\ab[6][47] ), .B(\CARRYB[5][47] ), .CI(\SUMB[5][48] ), 
        .CO(\CARRYB[6][47] ), .S(\SUMB[6][47] ) );
  FA1A S2_6_48 ( .A(\ab[6][48] ), .B(\CARRYB[5][48] ), .CI(\SUMB[5][49] ), 
        .CO(\CARRYB[6][48] ), .S(\SUMB[6][48] ) );
  FA1A S2_7_45 ( .A(\ab[7][45] ), .B(\CARRYB[6][45] ), .CI(\SUMB[6][46] ), 
        .CO(\CARRYB[7][45] ), .S(\SUMB[7][45] ) );
  FA1A S2_4_51 ( .A(\ab[4][51] ), .B(\CARRYB[3][51] ), .CI(\SUMB[3][52] ), 
        .CO(\CARRYB[4][51] ), .S(\SUMB[4][51] ) );
  FA1A S2_5_48 ( .A(\ab[5][48] ), .B(\CARRYB[4][48] ), .CI(\SUMB[4][49] ), 
        .CO(\CARRYB[5][48] ), .S(\SUMB[5][48] ) );
  FA1A S2_5_49 ( .A(\ab[5][49] ), .B(\CARRYB[4][49] ), .CI(\SUMB[4][50] ), 
        .CO(\CARRYB[5][49] ), .S(\SUMB[5][49] ) );
  FA1A S2_6_46 ( .A(\ab[6][46] ), .B(\CARRYB[5][46] ), .CI(\SUMB[5][47] ), 
        .CO(\CARRYB[6][46] ), .S(\SUMB[6][46] ) );
  FA1A S2_6_45 ( .A(\ab[6][45] ), .B(\CARRYB[5][45] ), .CI(\SUMB[5][46] ), 
        .CO(\CARRYB[6][45] ), .S(\SUMB[6][45] ) );
  FA1A S2_4_49 ( .A(\ab[4][49] ), .B(\CARRYB[3][49] ), .CI(\SUMB[3][50] ), 
        .CO(\CARRYB[4][49] ), .S(\SUMB[4][49] ) );
  FA1A S2_4_50 ( .A(\ab[4][50] ), .B(\CARRYB[3][50] ), .CI(\SUMB[3][51] ), 
        .CO(\CARRYB[4][50] ), .S(\SUMB[4][50] ) );
  FA1A S2_5_47 ( .A(\ab[5][47] ), .B(\CARRYB[4][47] ), .CI(\SUMB[4][48] ), 
        .CO(\CARRYB[5][47] ), .S(\SUMB[5][47] ) );
  FA1A S2_5_46 ( .A(\ab[5][46] ), .B(\CARRYB[4][46] ), .CI(\SUMB[4][47] ), 
        .CO(\CARRYB[5][46] ), .S(\SUMB[5][46] ) );
  FA1A S2_5_45 ( .A(\ab[5][45] ), .B(\CARRYB[4][45] ), .CI(\SUMB[4][46] ), 
        .CO(\CARRYB[5][45] ), .S(\SUMB[5][45] ) );
  FA1A S2_3_50 ( .A(\ab[3][50] ), .B(\CARRYB[2][50] ), .CI(\SUMB[2][51] ), 
        .CO(\CARRYB[3][50] ), .S(\SUMB[3][50] ) );
  FA1A S2_3_51 ( .A(\ab[3][51] ), .B(\CARRYB[2][51] ), .CI(\SUMB[2][52] ), 
        .CO(\CARRYB[3][51] ), .S(\SUMB[3][51] ) );
  FA1A S2_4_48 ( .A(\ab[4][48] ), .B(\CARRYB[3][48] ), .CI(\SUMB[3][49] ), 
        .CO(\CARRYB[4][48] ), .S(\SUMB[4][48] ) );
  FA1A S2_4_47 ( .A(\ab[4][47] ), .B(\CARRYB[3][47] ), .CI(\SUMB[3][48] ), 
        .CO(\CARRYB[4][47] ), .S(\SUMB[4][47] ) );
  FA1A S2_4_46 ( .A(\ab[4][46] ), .B(\CARRYB[3][46] ), .CI(\SUMB[3][47] ), 
        .CO(\CARRYB[4][46] ), .S(\SUMB[4][46] ) );
  FA1A S2_4_45 ( .A(\ab[4][45] ), .B(\CARRYB[3][45] ), .CI(\SUMB[3][46] ), 
        .CO(\CARRYB[4][45] ), .S(\SUMB[4][45] ) );
  FA1A S2_2_51 ( .A(\ab[2][51] ), .B(\CARRYB[1][51] ), .CI(\SUMB[1][52] ), 
        .CO(\CARRYB[2][51] ), .S(\SUMB[2][51] ) );
  FA1A S2_3_49 ( .A(\ab[3][49] ), .B(\CARRYB[2][49] ), .CI(\SUMB[2][50] ), 
        .CO(\CARRYB[3][49] ), .S(\SUMB[3][49] ) );
  FA1A S2_3_48 ( .A(\ab[3][48] ), .B(\CARRYB[2][48] ), .CI(\SUMB[2][49] ), 
        .CO(\CARRYB[3][48] ), .S(\SUMB[3][48] ) );
  FA1A S2_3_47 ( .A(\ab[3][47] ), .B(\CARRYB[2][47] ), .CI(\SUMB[2][48] ), 
        .CO(\CARRYB[3][47] ), .S(\SUMB[3][47] ) );
  FA1A S2_3_46 ( .A(\ab[3][46] ), .B(\CARRYB[2][46] ), .CI(\SUMB[2][47] ), 
        .CO(\CARRYB[3][46] ), .S(\SUMB[3][46] ) );
  FA1A S2_3_45 ( .A(\ab[3][45] ), .B(\CARRYB[2][45] ), .CI(\SUMB[2][46] ), 
        .CO(\CARRYB[3][45] ), .S(\SUMB[3][45] ) );
  FA1A S2_2_50 ( .A(\ab[2][50] ), .B(\CARRYB[1][50] ), .CI(\SUMB[1][51] ), 
        .CO(\CARRYB[2][50] ), .S(\SUMB[2][50] ) );
  FA1A S2_2_49 ( .A(\ab[2][49] ), .B(\CARRYB[1][49] ), .CI(\SUMB[1][50] ), 
        .CO(\CARRYB[2][49] ), .S(\SUMB[2][49] ) );
  FA1A S2_2_48 ( .A(\ab[2][48] ), .B(\CARRYB[1][48] ), .CI(\SUMB[1][49] ), 
        .CO(\CARRYB[2][48] ), .S(\SUMB[2][48] ) );
  FA1A S2_2_47 ( .A(\ab[2][47] ), .B(\CARRYB[1][47] ), .CI(\SUMB[1][48] ), 
        .CO(\CARRYB[2][47] ), .S(\SUMB[2][47] ) );
  FA1A S2_2_46 ( .A(\ab[2][46] ), .B(\CARRYB[1][46] ), .CI(\SUMB[1][47] ), 
        .CO(\CARRYB[2][46] ), .S(\SUMB[2][46] ) );
  FA1A S2_2_45 ( .A(\ab[2][45] ), .B(\CARRYB[1][45] ), .CI(\SUMB[1][46] ), 
        .CO(\CARRYB[2][45] ), .S(\SUMB[2][45] ) );
  FA1A S5_94 ( .A(\ab[29][94] ), .B(\CARRYB[28][94] ), .CI(\ab[28][95] ), .CO(
        \CARRYB[29][94] ), .S(\SUMB[29][94] ) );
  FA1A S4_93 ( .A(\ab[29][93] ), .B(\CARRYB[28][93] ), .CI(\SUMB[28][94] ), 
        .CO(\CARRYB[29][93] ), .S(\SUMB[29][93] ) );
  FA1A S4_92 ( .A(\ab[29][92] ), .B(\CARRYB[28][92] ), .CI(\SUMB[28][93] ), 
        .CO(\CARRYB[29][92] ), .S(\SUMB[29][92] ) );
  FA1A S4_91 ( .A(\ab[29][91] ), .B(\CARRYB[28][91] ), .CI(\SUMB[28][92] ), 
        .CO(\CARRYB[29][91] ), .S(\SUMB[29][91] ) );
  FA1A S4_90 ( .A(\ab[29][90] ), .B(\CARRYB[28][90] ), .CI(\SUMB[28][91] ), 
        .CO(\CARRYB[29][90] ), .S(\SUMB[29][90] ) );
  FA1A S3_28_94 ( .A(\ab[28][94] ), .B(\CARRYB[27][94] ), .CI(\ab[27][95] ), 
        .CO(\CARRYB[28][94] ), .S(\SUMB[28][94] ) );
  FA1A S2_28_93 ( .A(\ab[28][93] ), .B(\CARRYB[27][93] ), .CI(\SUMB[27][94] ), 
        .CO(\CARRYB[28][93] ), .S(\SUMB[28][93] ) );
  FA1A S2_28_92 ( .A(\ab[28][92] ), .B(\CARRYB[27][92] ), .CI(\SUMB[27][93] ), 
        .CO(\CARRYB[28][92] ), .S(\SUMB[28][92] ) );
  FA1A S2_28_91 ( .A(\ab[28][91] ), .B(\CARRYB[27][91] ), .CI(\SUMB[27][92] ), 
        .CO(\CARRYB[28][91] ), .S(\SUMB[28][91] ) );
  FA1A S3_27_94 ( .A(\ab[27][94] ), .B(\CARRYB[26][94] ), .CI(\ab[26][95] ), 
        .CO(\CARRYB[27][94] ), .S(\SUMB[27][94] ) );
  FA1A S2_27_93 ( .A(\ab[27][93] ), .B(\CARRYB[26][93] ), .CI(\SUMB[26][94] ), 
        .CO(\CARRYB[27][93] ), .S(\SUMB[27][93] ) );
  FA1A S2_27_92 ( .A(\ab[27][92] ), .B(\CARRYB[26][92] ), .CI(\SUMB[26][93] ), 
        .CO(\CARRYB[27][92] ), .S(\SUMB[27][92] ) );
  FA1A S3_26_94 ( .A(\ab[26][94] ), .B(\CARRYB[25][94] ), .CI(\ab[25][95] ), 
        .CO(\CARRYB[26][94] ), .S(\SUMB[26][94] ) );
  FA1A S2_26_93 ( .A(\ab[26][93] ), .B(\CARRYB[25][93] ), .CI(\SUMB[25][94] ), 
        .CO(\CARRYB[26][93] ), .S(\SUMB[26][93] ) );
  FA1A S3_25_94 ( .A(\ab[25][94] ), .B(\CARRYB[24][94] ), .CI(\ab[24][95] ), 
        .CO(\CARRYB[25][94] ), .S(\SUMB[25][94] ) );
  FA1A S3_24_94 ( .A(\ab[24][94] ), .B(\CARRYB[23][94] ), .CI(\ab[23][95] ), 
        .CO(\CARRYB[24][94] ), .S(\SUMB[24][94] ) );
  FA1A S3_23_94 ( .A(\ab[23][94] ), .B(\CARRYB[22][94] ), .CI(\ab[22][95] ), 
        .CO(\CARRYB[23][94] ), .S(\SUMB[23][94] ) );
  FA1A S3_22_94 ( .A(\ab[22][94] ), .B(\CARRYB[21][94] ), .CI(\ab[21][95] ), 
        .CO(\CARRYB[22][94] ), .S(\SUMB[22][94] ) );
  FA1A S3_21_94 ( .A(\ab[21][94] ), .B(\CARRYB[20][94] ), .CI(\ab[20][95] ), 
        .CO(\CARRYB[21][94] ), .S(\SUMB[21][94] ) );
  FA1A S3_20_94 ( .A(\ab[20][94] ), .B(\CARRYB[19][94] ), .CI(\ab[19][95] ), 
        .CO(\CARRYB[20][94] ), .S(\SUMB[20][94] ) );
  FA1A S2_25_93 ( .A(\ab[25][93] ), .B(\CARRYB[24][93] ), .CI(\SUMB[24][94] ), 
        .CO(\CARRYB[25][93] ), .S(\SUMB[25][93] ) );
  FA1A S2_24_93 ( .A(\ab[24][93] ), .B(\CARRYB[23][93] ), .CI(\SUMB[23][94] ), 
        .CO(\CARRYB[24][93] ), .S(\SUMB[24][93] ) );
  FA1A S2_23_93 ( .A(\ab[23][93] ), .B(\CARRYB[22][93] ), .CI(\SUMB[22][94] ), 
        .CO(\CARRYB[23][93] ), .S(\SUMB[23][93] ) );
  FA1A S2_22_93 ( .A(\ab[22][93] ), .B(\CARRYB[21][93] ), .CI(\SUMB[21][94] ), 
        .CO(\CARRYB[22][93] ), .S(\SUMB[22][93] ) );
  FA1A S2_21_93 ( .A(\ab[21][93] ), .B(\CARRYB[20][93] ), .CI(\SUMB[20][94] ), 
        .CO(\CARRYB[21][93] ), .S(\SUMB[21][93] ) );
  FA1A S3_19_94 ( .A(\ab[19][94] ), .B(\CARRYB[18][94] ), .CI(\ab[18][95] ), 
        .CO(\CARRYB[19][94] ), .S(\SUMB[19][94] ) );
  FA1A S3_18_94 ( .A(\ab[18][94] ), .B(\CARRYB[17][94] ), .CI(\ab[17][95] ), 
        .CO(\CARRYB[18][94] ), .S(\SUMB[18][94] ) );
  FA1A S3_17_94 ( .A(\ab[17][94] ), .B(\CARRYB[16][94] ), .CI(\ab[16][95] ), 
        .CO(\CARRYB[17][94] ), .S(\SUMB[17][94] ) );
  FA1A S3_16_94 ( .A(\ab[16][94] ), .B(\CARRYB[15][94] ), .CI(\ab[15][95] ), 
        .CO(\CARRYB[16][94] ), .S(\SUMB[16][94] ) );
  FA1A S3_15_94 ( .A(\ab[15][94] ), .B(\CARRYB[14][94] ), .CI(\ab[14][95] ), 
        .CO(\CARRYB[15][94] ), .S(\SUMB[15][94] ) );
  FA1A S2_20_93 ( .A(\ab[20][93] ), .B(\CARRYB[19][93] ), .CI(\SUMB[19][94] ), 
        .CO(\CARRYB[20][93] ), .S(\SUMB[20][93] ) );
  FA1A S2_19_93 ( .A(\ab[19][93] ), .B(\CARRYB[18][93] ), .CI(\SUMB[18][94] ), 
        .CO(\CARRYB[19][93] ), .S(\SUMB[19][93] ) );
  FA1A S2_18_93 ( .A(\ab[18][93] ), .B(\CARRYB[17][93] ), .CI(\SUMB[17][94] ), 
        .CO(\CARRYB[18][93] ), .S(\SUMB[18][93] ) );
  FA1A S2_17_93 ( .A(\ab[17][93] ), .B(\CARRYB[16][93] ), .CI(\SUMB[16][94] ), 
        .CO(\CARRYB[17][93] ), .S(\SUMB[17][93] ) );
  FA1A S2_16_93 ( .A(\ab[16][93] ), .B(\CARRYB[15][93] ), .CI(\SUMB[15][94] ), 
        .CO(\CARRYB[16][93] ), .S(\SUMB[16][93] ) );
  FA1A S2_15_93 ( .A(\ab[15][93] ), .B(\CARRYB[14][93] ), .CI(\SUMB[14][94] ), 
        .CO(\CARRYB[15][93] ), .S(\SUMB[15][93] ) );
  FA1A S2_26_92 ( .A(\ab[26][92] ), .B(\CARRYB[25][92] ), .CI(\SUMB[25][93] ), 
        .CO(\CARRYB[26][92] ), .S(\SUMB[26][92] ) );
  FA1A S2_25_92 ( .A(\ab[25][92] ), .B(\CARRYB[24][92] ), .CI(\SUMB[24][93] ), 
        .CO(\CARRYB[25][92] ), .S(\SUMB[25][92] ) );
  FA1A S2_24_92 ( .A(\ab[24][92] ), .B(\CARRYB[23][92] ), .CI(\SUMB[23][93] ), 
        .CO(\CARRYB[24][92] ), .S(\SUMB[24][92] ) );
  FA1A S2_23_92 ( .A(\ab[23][92] ), .B(\CARRYB[22][92] ), .CI(\SUMB[22][93] ), 
        .CO(\CARRYB[23][92] ), .S(\SUMB[23][92] ) );
  FA1A S2_22_92 ( .A(\ab[22][92] ), .B(\CARRYB[21][92] ), .CI(\SUMB[21][93] ), 
        .CO(\CARRYB[22][92] ), .S(\SUMB[22][92] ) );
  FA1A S2_27_91 ( .A(\ab[27][91] ), .B(\CARRYB[26][91] ), .CI(\SUMB[26][92] ), 
        .CO(\CARRYB[27][91] ), .S(\SUMB[27][91] ) );
  FA1A S2_26_91 ( .A(\ab[26][91] ), .B(\CARRYB[25][91] ), .CI(\SUMB[25][92] ), 
        .CO(\CARRYB[26][91] ), .S(\SUMB[26][91] ) );
  FA1A S2_25_91 ( .A(\ab[25][91] ), .B(\CARRYB[24][91] ), .CI(\SUMB[24][92] ), 
        .CO(\CARRYB[25][91] ), .S(\SUMB[25][91] ) );
  FA1A S2_24_91 ( .A(\ab[24][91] ), .B(\CARRYB[23][91] ), .CI(\SUMB[23][92] ), 
        .CO(\CARRYB[24][91] ), .S(\SUMB[24][91] ) );
  FA1A S2_23_91 ( .A(\ab[23][91] ), .B(\CARRYB[22][91] ), .CI(\SUMB[22][92] ), 
        .CO(\CARRYB[23][91] ), .S(\SUMB[23][91] ) );
  FA1A S2_21_92 ( .A(\ab[21][92] ), .B(\CARRYB[20][92] ), .CI(\SUMB[20][93] ), 
        .CO(\CARRYB[21][92] ), .S(\SUMB[21][92] ) );
  FA1A S2_20_92 ( .A(\ab[20][92] ), .B(\CARRYB[19][92] ), .CI(\SUMB[19][93] ), 
        .CO(\CARRYB[20][92] ), .S(\SUMB[20][92] ) );
  FA1A S2_19_92 ( .A(\ab[19][92] ), .B(\CARRYB[18][92] ), .CI(\SUMB[18][93] ), 
        .CO(\CARRYB[19][92] ), .S(\SUMB[19][92] ) );
  FA1A S2_18_92 ( .A(\ab[18][92] ), .B(\CARRYB[17][92] ), .CI(\SUMB[17][93] ), 
        .CO(\CARRYB[18][92] ), .S(\SUMB[18][92] ) );
  FA1A S2_17_92 ( .A(\ab[17][92] ), .B(\CARRYB[16][92] ), .CI(\SUMB[16][93] ), 
        .CO(\CARRYB[17][92] ), .S(\SUMB[17][92] ) );
  FA1A S2_16_92 ( .A(\ab[16][92] ), .B(\CARRYB[15][92] ), .CI(\SUMB[15][93] ), 
        .CO(\CARRYB[16][92] ), .S(\SUMB[16][92] ) );
  FA1A S2_15_92 ( .A(\ab[15][92] ), .B(\CARRYB[14][92] ), .CI(\SUMB[14][93] ), 
        .CO(\CARRYB[15][92] ), .S(\SUMB[15][92] ) );
  FA1A S2_28_90 ( .A(\ab[28][90] ), .B(\CARRYB[27][90] ), .CI(\SUMB[27][91] ), 
        .CO(\CARRYB[28][90] ), .S(\SUMB[28][90] ) );
  FA1A S2_27_90 ( .A(\ab[27][90] ), .B(\CARRYB[26][90] ), .CI(\SUMB[26][91] ), 
        .CO(\CARRYB[27][90] ), .S(\SUMB[27][90] ) );
  FA1A S2_26_90 ( .A(\ab[26][90] ), .B(\CARRYB[25][90] ), .CI(\SUMB[25][91] ), 
        .CO(\CARRYB[26][90] ), .S(\SUMB[26][90] ) );
  FA1A S2_25_90 ( .A(\ab[25][90] ), .B(\CARRYB[24][90] ), .CI(\SUMB[24][91] ), 
        .CO(\CARRYB[25][90] ), .S(\SUMB[25][90] ) );
  FA1A S2_24_90 ( .A(\ab[24][90] ), .B(\CARRYB[23][90] ), .CI(\SUMB[23][91] ), 
        .CO(\CARRYB[24][90] ), .S(\SUMB[24][90] ) );
  FA1A S2_22_91 ( .A(\ab[22][91] ), .B(\CARRYB[21][91] ), .CI(\SUMB[21][92] ), 
        .CO(\CARRYB[22][91] ), .S(\SUMB[22][91] ) );
  FA1A S2_21_91 ( .A(\ab[21][91] ), .B(\CARRYB[20][91] ), .CI(\SUMB[20][92] ), 
        .CO(\CARRYB[21][91] ), .S(\SUMB[21][91] ) );
  FA1A S2_20_91 ( .A(\ab[20][91] ), .B(\CARRYB[19][91] ), .CI(\SUMB[19][92] ), 
        .CO(\CARRYB[20][91] ), .S(\SUMB[20][91] ) );
  FA1A S2_19_91 ( .A(\ab[19][91] ), .B(\CARRYB[18][91] ), .CI(\SUMB[18][92] ), 
        .CO(\CARRYB[19][91] ), .S(\SUMB[19][91] ) );
  FA1A S2_18_91 ( .A(\ab[18][91] ), .B(\CARRYB[17][91] ), .CI(\SUMB[17][92] ), 
        .CO(\CARRYB[18][91] ), .S(\SUMB[18][91] ) );
  FA1A S2_17_91 ( .A(\ab[17][91] ), .B(\CARRYB[16][91] ), .CI(\SUMB[16][92] ), 
        .CO(\CARRYB[17][91] ), .S(\SUMB[17][91] ) );
  FA1A S2_16_91 ( .A(\ab[16][91] ), .B(\CARRYB[15][91] ), .CI(\SUMB[15][92] ), 
        .CO(\CARRYB[16][91] ), .S(\SUMB[16][91] ) );
  FA1A S2_15_91 ( .A(\ab[15][91] ), .B(\CARRYB[14][91] ), .CI(\SUMB[14][92] ), 
        .CO(\CARRYB[15][91] ), .S(\SUMB[15][91] ) );
  FA1A S2_28_89 ( .A(\ab[28][89] ), .B(\CARRYB[27][89] ), .CI(\SUMB[27][90] ), 
        .CO(\CARRYB[28][89] ), .S(\SUMB[28][89] ) );
  FA1A S2_27_89 ( .A(\ab[27][89] ), .B(\CARRYB[26][89] ), .CI(\SUMB[26][90] ), 
        .CO(\CARRYB[27][89] ), .S(\SUMB[27][89] ) );
  FA1A S2_26_89 ( .A(\ab[26][89] ), .B(\CARRYB[25][89] ), .CI(\SUMB[25][90] ), 
        .CO(\CARRYB[26][89] ), .S(\SUMB[26][89] ) );
  FA1A S2_25_89 ( .A(\ab[25][89] ), .B(\CARRYB[24][89] ), .CI(\SUMB[24][90] ), 
        .CO(\CARRYB[25][89] ), .S(\SUMB[25][89] ) );
  FA1A S2_23_90 ( .A(\ab[23][90] ), .B(\CARRYB[22][90] ), .CI(\SUMB[22][91] ), 
        .CO(\CARRYB[23][90] ), .S(\SUMB[23][90] ) );
  FA1A S2_22_90 ( .A(\ab[22][90] ), .B(\CARRYB[21][90] ), .CI(\SUMB[21][91] ), 
        .CO(\CARRYB[22][90] ), .S(\SUMB[22][90] ) );
  FA1A S2_21_90 ( .A(\ab[21][90] ), .B(\CARRYB[20][90] ), .CI(\SUMB[20][91] ), 
        .CO(\CARRYB[21][90] ), .S(\SUMB[21][90] ) );
  FA1A S2_20_90 ( .A(\ab[20][90] ), .B(\CARRYB[19][90] ), .CI(\SUMB[19][91] ), 
        .CO(\CARRYB[20][90] ), .S(\SUMB[20][90] ) );
  FA1A S2_19_90 ( .A(\ab[19][90] ), .B(\CARRYB[18][90] ), .CI(\SUMB[18][91] ), 
        .CO(\CARRYB[19][90] ), .S(\SUMB[19][90] ) );
  FA1A S2_18_90 ( .A(\ab[18][90] ), .B(\CARRYB[17][90] ), .CI(\SUMB[17][91] ), 
        .CO(\CARRYB[18][90] ), .S(\SUMB[18][90] ) );
  FA1A S2_17_90 ( .A(\ab[17][90] ), .B(\CARRYB[16][90] ), .CI(\SUMB[16][91] ), 
        .CO(\CARRYB[17][90] ), .S(\SUMB[17][90] ) );
  FA1A S2_16_90 ( .A(\ab[16][90] ), .B(\CARRYB[15][90] ), .CI(\SUMB[15][91] ), 
        .CO(\CARRYB[16][90] ), .S(\SUMB[16][90] ) );
  FA1A S2_15_90 ( .A(\ab[15][90] ), .B(\CARRYB[14][90] ), .CI(\SUMB[14][91] ), 
        .CO(\CARRYB[15][90] ), .S(\SUMB[15][90] ) );
  FA1A S4_89 ( .A(\ab[29][89] ), .B(\CARRYB[28][89] ), .CI(\SUMB[28][90] ), 
        .CO(\CARRYB[29][89] ), .S(\SUMB[29][89] ) );
  FA1A S2_28_88 ( .A(\ab[28][88] ), .B(\CARRYB[27][88] ), .CI(\SUMB[27][89] ), 
        .CO(\CARRYB[28][88] ), .S(\SUMB[28][88] ) );
  FA1A S2_27_88 ( .A(\ab[27][88] ), .B(\CARRYB[26][88] ), .CI(\SUMB[26][89] ), 
        .CO(\CARRYB[27][88] ), .S(\SUMB[27][88] ) );
  FA1A S2_26_88 ( .A(\ab[26][88] ), .B(\CARRYB[25][88] ), .CI(\SUMB[25][89] ), 
        .CO(\CARRYB[26][88] ), .S(\SUMB[26][88] ) );
  FA1A S2_24_89 ( .A(\ab[24][89] ), .B(\CARRYB[23][89] ), .CI(\SUMB[23][90] ), 
        .CO(\CARRYB[24][89] ), .S(\SUMB[24][89] ) );
  FA1A S2_23_89 ( .A(\ab[23][89] ), .B(\CARRYB[22][89] ), .CI(\SUMB[22][90] ), 
        .CO(\CARRYB[23][89] ), .S(\SUMB[23][89] ) );
  FA1A S2_22_89 ( .A(\ab[22][89] ), .B(\CARRYB[21][89] ), .CI(\SUMB[21][90] ), 
        .CO(\CARRYB[22][89] ), .S(\SUMB[22][89] ) );
  FA1A S2_21_89 ( .A(\ab[21][89] ), .B(\CARRYB[20][89] ), .CI(\SUMB[20][90] ), 
        .CO(\CARRYB[21][89] ), .S(\SUMB[21][89] ) );
  FA1A S2_20_89 ( .A(\ab[20][89] ), .B(\CARRYB[19][89] ), .CI(\SUMB[19][90] ), 
        .CO(\CARRYB[20][89] ), .S(\SUMB[20][89] ) );
  FA1A S2_19_89 ( .A(\ab[19][89] ), .B(\CARRYB[18][89] ), .CI(\SUMB[18][90] ), 
        .CO(\CARRYB[19][89] ), .S(\SUMB[19][89] ) );
  FA1A S2_18_89 ( .A(\ab[18][89] ), .B(\CARRYB[17][89] ), .CI(\SUMB[17][90] ), 
        .CO(\CARRYB[18][89] ), .S(\SUMB[18][89] ) );
  FA1A S2_17_89 ( .A(\ab[17][89] ), .B(\CARRYB[16][89] ), .CI(\SUMB[16][90] ), 
        .CO(\CARRYB[17][89] ), .S(\SUMB[17][89] ) );
  FA1A S2_16_89 ( .A(\ab[16][89] ), .B(\CARRYB[15][89] ), .CI(\SUMB[15][90] ), 
        .CO(\CARRYB[16][89] ), .S(\SUMB[16][89] ) );
  FA1A S2_15_89 ( .A(\ab[15][89] ), .B(\CARRYB[14][89] ), .CI(\SUMB[14][90] ), 
        .CO(\CARRYB[15][89] ), .S(\SUMB[15][89] ) );
  FA1A S4_88 ( .A(\ab[29][88] ), .B(\CARRYB[28][88] ), .CI(\SUMB[28][89] ), 
        .CO(\CARRYB[29][88] ), .S(\SUMB[29][88] ) );
  FA1A S2_28_87 ( .A(\ab[28][87] ), .B(\CARRYB[27][87] ), .CI(\SUMB[27][88] ), 
        .CO(\CARRYB[28][87] ), .S(\SUMB[28][87] ) );
  FA1A S2_27_87 ( .A(\ab[27][87] ), .B(\CARRYB[26][87] ), .CI(\SUMB[26][88] ), 
        .CO(\CARRYB[27][87] ), .S(\SUMB[27][87] ) );
  FA1A S4_87 ( .A(\ab[29][87] ), .B(\CARRYB[28][87] ), .CI(\SUMB[28][88] ), 
        .CO(\CARRYB[29][87] ), .S(\SUMB[29][87] ) );
  FA1A S2_28_86 ( .A(\ab[28][86] ), .B(\CARRYB[27][86] ), .CI(\SUMB[27][87] ), 
        .CO(\CARRYB[28][86] ), .S(\SUMB[28][86] ) );
  FA1A S2_25_88 ( .A(\ab[25][88] ), .B(\CARRYB[24][88] ), .CI(\SUMB[24][89] ), 
        .CO(\CARRYB[25][88] ), .S(\SUMB[25][88] ) );
  FA1A S2_24_88 ( .A(\ab[24][88] ), .B(\CARRYB[23][88] ), .CI(\SUMB[23][89] ), 
        .CO(\CARRYB[24][88] ), .S(\SUMB[24][88] ) );
  FA1A S2_23_88 ( .A(\ab[23][88] ), .B(\CARRYB[22][88] ), .CI(\SUMB[22][89] ), 
        .CO(\CARRYB[23][88] ), .S(\SUMB[23][88] ) );
  FA1A S2_22_88 ( .A(\ab[22][88] ), .B(\CARRYB[21][88] ), .CI(\SUMB[21][89] ), 
        .CO(\CARRYB[22][88] ), .S(\SUMB[22][88] ) );
  FA1A S2_21_88 ( .A(\ab[21][88] ), .B(\CARRYB[20][88] ), .CI(\SUMB[20][89] ), 
        .CO(\CARRYB[21][88] ), .S(\SUMB[21][88] ) );
  FA1A S2_20_88 ( .A(\ab[20][88] ), .B(\CARRYB[19][88] ), .CI(\SUMB[19][89] ), 
        .CO(\CARRYB[20][88] ), .S(\SUMB[20][88] ) );
  FA1A S2_19_88 ( .A(\ab[19][88] ), .B(\CARRYB[18][88] ), .CI(\SUMB[18][89] ), 
        .CO(\CARRYB[19][88] ), .S(\SUMB[19][88] ) );
  FA1A S2_18_88 ( .A(\ab[18][88] ), .B(\CARRYB[17][88] ), .CI(\SUMB[17][89] ), 
        .CO(\CARRYB[18][88] ), .S(\SUMB[18][88] ) );
  FA1A S2_17_88 ( .A(\ab[17][88] ), .B(\CARRYB[16][88] ), .CI(\SUMB[16][89] ), 
        .CO(\CARRYB[17][88] ), .S(\SUMB[17][88] ) );
  FA1A S2_16_88 ( .A(\ab[16][88] ), .B(\CARRYB[15][88] ), .CI(\SUMB[15][89] ), 
        .CO(\CARRYB[16][88] ), .S(\SUMB[16][88] ) );
  FA1A S2_15_88 ( .A(\ab[15][88] ), .B(\CARRYB[14][88] ), .CI(\SUMB[14][89] ), 
        .CO(\CARRYB[15][88] ), .S(\SUMB[15][88] ) );
  FA1A S4_86 ( .A(\ab[29][86] ), .B(\CARRYB[28][86] ), .CI(\SUMB[28][87] ), 
        .CO(\CARRYB[29][86] ), .S(\SUMB[29][86] ) );
  FA1A S2_26_87 ( .A(\ab[26][87] ), .B(\CARRYB[25][87] ), .CI(\SUMB[25][88] ), 
        .CO(\CARRYB[26][87] ), .S(\SUMB[26][87] ) );
  FA1A S2_25_87 ( .A(\ab[25][87] ), .B(\CARRYB[24][87] ), .CI(\SUMB[24][88] ), 
        .CO(\CARRYB[25][87] ), .S(\SUMB[25][87] ) );
  FA1A S2_24_87 ( .A(\ab[24][87] ), .B(\CARRYB[23][87] ), .CI(\SUMB[23][88] ), 
        .CO(\CARRYB[24][87] ), .S(\SUMB[24][87] ) );
  FA1A S2_23_87 ( .A(\ab[23][87] ), .B(\CARRYB[22][87] ), .CI(\SUMB[22][88] ), 
        .CO(\CARRYB[23][87] ), .S(\SUMB[23][87] ) );
  FA1A S2_22_87 ( .A(\ab[22][87] ), .B(\CARRYB[21][87] ), .CI(\SUMB[21][88] ), 
        .CO(\CARRYB[22][87] ), .S(\SUMB[22][87] ) );
  FA1A S2_21_87 ( .A(\ab[21][87] ), .B(\CARRYB[20][87] ), .CI(\SUMB[20][88] ), 
        .CO(\CARRYB[21][87] ), .S(\SUMB[21][87] ) );
  FA1A S2_20_87 ( .A(\ab[20][87] ), .B(\CARRYB[19][87] ), .CI(\SUMB[19][88] ), 
        .CO(\CARRYB[20][87] ), .S(\SUMB[20][87] ) );
  FA1A S2_19_87 ( .A(\ab[19][87] ), .B(\CARRYB[18][87] ), .CI(\SUMB[18][88] ), 
        .CO(\CARRYB[19][87] ), .S(\SUMB[19][87] ) );
  FA1A S2_18_87 ( .A(\ab[18][87] ), .B(\CARRYB[17][87] ), .CI(\SUMB[17][88] ), 
        .CO(\CARRYB[18][87] ), .S(\SUMB[18][87] ) );
  FA1A S2_17_87 ( .A(\ab[17][87] ), .B(\CARRYB[16][87] ), .CI(\SUMB[16][88] ), 
        .CO(\CARRYB[17][87] ), .S(\SUMB[17][87] ) );
  FA1A S2_16_87 ( .A(\ab[16][87] ), .B(\CARRYB[15][87] ), .CI(\SUMB[15][88] ), 
        .CO(\CARRYB[16][87] ), .S(\SUMB[16][87] ) );
  FA1A S2_15_87 ( .A(\ab[15][87] ), .B(\CARRYB[14][87] ), .CI(\SUMB[14][88] ), 
        .CO(\CARRYB[15][87] ), .S(\SUMB[15][87] ) );
  FA1A S4_85 ( .A(\ab[29][85] ), .B(\CARRYB[28][85] ), .CI(\SUMB[28][86] ), 
        .CO(\CARRYB[29][85] ), .S(\SUMB[29][85] ) );
  FA1A S2_27_86 ( .A(\ab[27][86] ), .B(\CARRYB[26][86] ), .CI(\SUMB[26][87] ), 
        .CO(\CARRYB[27][86] ), .S(\SUMB[27][86] ) );
  FA1A S2_26_86 ( .A(\ab[26][86] ), .B(\CARRYB[25][86] ), .CI(\SUMB[25][87] ), 
        .CO(\CARRYB[26][86] ), .S(\SUMB[26][86] ) );
  FA1A S2_25_86 ( .A(\ab[25][86] ), .B(\CARRYB[24][86] ), .CI(\SUMB[24][87] ), 
        .CO(\CARRYB[25][86] ), .S(\SUMB[25][86] ) );
  FA1A S2_24_86 ( .A(\ab[24][86] ), .B(\CARRYB[23][86] ), .CI(\SUMB[23][87] ), 
        .CO(\CARRYB[24][86] ), .S(\SUMB[24][86] ) );
  FA1A S2_23_86 ( .A(\ab[23][86] ), .B(\CARRYB[22][86] ), .CI(\SUMB[22][87] ), 
        .CO(\CARRYB[23][86] ), .S(\SUMB[23][86] ) );
  FA1A S2_22_86 ( .A(\ab[22][86] ), .B(\CARRYB[21][86] ), .CI(\SUMB[21][87] ), 
        .CO(\CARRYB[22][86] ), .S(\SUMB[22][86] ) );
  FA1A S2_21_86 ( .A(\ab[21][86] ), .B(\CARRYB[20][86] ), .CI(\SUMB[20][87] ), 
        .CO(\CARRYB[21][86] ), .S(\SUMB[21][86] ) );
  FA1A S2_20_86 ( .A(\ab[20][86] ), .B(\CARRYB[19][86] ), .CI(\SUMB[19][87] ), 
        .CO(\CARRYB[20][86] ), .S(\SUMB[20][86] ) );
  FA1A S2_19_86 ( .A(\ab[19][86] ), .B(\CARRYB[18][86] ), .CI(\SUMB[18][87] ), 
        .CO(\CARRYB[19][86] ), .S(\SUMB[19][86] ) );
  FA1A S2_18_86 ( .A(\ab[18][86] ), .B(\CARRYB[17][86] ), .CI(\SUMB[17][87] ), 
        .CO(\CARRYB[18][86] ), .S(\SUMB[18][86] ) );
  FA1A S2_17_86 ( .A(\ab[17][86] ), .B(\CARRYB[16][86] ), .CI(\SUMB[16][87] ), 
        .CO(\CARRYB[17][86] ), .S(\SUMB[17][86] ) );
  FA1A S2_16_86 ( .A(\ab[16][86] ), .B(\CARRYB[15][86] ), .CI(\SUMB[15][87] ), 
        .CO(\CARRYB[16][86] ), .S(\SUMB[16][86] ) );
  FA1A S2_15_86 ( .A(\ab[15][86] ), .B(\CARRYB[14][86] ), .CI(\SUMB[14][87] ), 
        .CO(\CARRYB[15][86] ), .S(\SUMB[15][86] ) );
  FA1A S2_28_85 ( .A(\ab[28][85] ), .B(\CARRYB[27][85] ), .CI(\SUMB[27][86] ), 
        .CO(\CARRYB[28][85] ), .S(\SUMB[28][85] ) );
  FA1A S2_27_85 ( .A(\ab[27][85] ), .B(\CARRYB[26][85] ), .CI(\SUMB[26][86] ), 
        .CO(\CARRYB[27][85] ), .S(\SUMB[27][85] ) );
  FA1A S2_26_85 ( .A(\ab[26][85] ), .B(\CARRYB[25][85] ), .CI(\SUMB[25][86] ), 
        .CO(\CARRYB[26][85] ), .S(\SUMB[26][85] ) );
  FA1A S2_25_85 ( .A(\ab[25][85] ), .B(\CARRYB[24][85] ), .CI(\SUMB[24][86] ), 
        .CO(\CARRYB[25][85] ), .S(\SUMB[25][85] ) );
  FA1A S2_24_85 ( .A(\ab[24][85] ), .B(\CARRYB[23][85] ), .CI(\SUMB[23][86] ), 
        .CO(\CARRYB[24][85] ), .S(\SUMB[24][85] ) );
  FA1A S2_23_85 ( .A(\ab[23][85] ), .B(\CARRYB[22][85] ), .CI(\SUMB[22][86] ), 
        .CO(\CARRYB[23][85] ), .S(\SUMB[23][85] ) );
  FA1A S2_22_85 ( .A(\ab[22][85] ), .B(\CARRYB[21][85] ), .CI(\SUMB[21][86] ), 
        .CO(\CARRYB[22][85] ), .S(\SUMB[22][85] ) );
  FA1A S2_21_85 ( .A(\ab[21][85] ), .B(\CARRYB[20][85] ), .CI(\SUMB[20][86] ), 
        .CO(\CARRYB[21][85] ), .S(\SUMB[21][85] ) );
  FA1A S2_20_85 ( .A(\ab[20][85] ), .B(\CARRYB[19][85] ), .CI(\SUMB[19][86] ), 
        .CO(\CARRYB[20][85] ), .S(\SUMB[20][85] ) );
  FA1A S2_19_85 ( .A(\ab[19][85] ), .B(\CARRYB[18][85] ), .CI(\SUMB[18][86] ), 
        .CO(\CARRYB[19][85] ), .S(\SUMB[19][85] ) );
  FA1A S2_18_85 ( .A(\ab[18][85] ), .B(\CARRYB[17][85] ), .CI(\SUMB[17][86] ), 
        .CO(\CARRYB[18][85] ), .S(\SUMB[18][85] ) );
  FA1A S2_17_85 ( .A(\ab[17][85] ), .B(\CARRYB[16][85] ), .CI(\SUMB[16][86] ), 
        .CO(\CARRYB[17][85] ), .S(\SUMB[17][85] ) );
  FA1A S2_16_85 ( .A(\ab[16][85] ), .B(\CARRYB[15][85] ), .CI(\SUMB[15][86] ), 
        .CO(\CARRYB[16][85] ), .S(\SUMB[16][85] ) );
  FA1A S2_15_85 ( .A(\ab[15][85] ), .B(\CARRYB[14][85] ), .CI(\SUMB[14][86] ), 
        .CO(\CARRYB[15][85] ), .S(\SUMB[15][85] ) );
  FA1A S4_80 ( .A(\ab[29][80] ), .B(\CARRYB[28][80] ), .CI(\SUMB[28][81] ), 
        .CO(\CARRYB[29][80] ), .S(\SUMB[29][80] ) );
  FA1A S4_81 ( .A(\ab[29][81] ), .B(\CARRYB[28][81] ), .CI(\SUMB[28][82] ), 
        .CO(\CARRYB[29][81] ), .S(\SUMB[29][81] ) );
  FA1A S2_28_81 ( .A(\ab[28][81] ), .B(\CARRYB[27][81] ), .CI(\SUMB[27][82] ), 
        .CO(\CARRYB[28][81] ), .S(\SUMB[28][81] ) );
  FA1A S2_27_81 ( .A(\ab[27][81] ), .B(\CARRYB[26][81] ), .CI(\SUMB[26][82] ), 
        .CO(\CARRYB[27][81] ), .S(\SUMB[27][81] ) );
  FA1A S2_26_81 ( .A(\ab[26][81] ), .B(\CARRYB[25][81] ), .CI(\SUMB[25][82] ), 
        .CO(\CARRYB[26][81] ), .S(\SUMB[26][81] ) );
  FA1A S2_25_81 ( .A(\ab[25][81] ), .B(\CARRYB[24][81] ), .CI(\SUMB[24][82] ), 
        .CO(\CARRYB[25][81] ), .S(\SUMB[25][81] ) );
  FA1A S2_24_81 ( .A(\ab[24][81] ), .B(\CARRYB[23][81] ), .CI(\SUMB[23][82] ), 
        .CO(\CARRYB[24][81] ), .S(\SUMB[24][81] ) );
  FA1A S2_23_81 ( .A(\ab[23][81] ), .B(\CARRYB[22][81] ), .CI(\SUMB[22][82] ), 
        .CO(\CARRYB[23][81] ), .S(\SUMB[23][81] ) );
  FA1A S2_22_81 ( .A(\ab[22][81] ), .B(\CARRYB[21][81] ), .CI(\SUMB[21][82] ), 
        .CO(\CARRYB[22][81] ), .S(\SUMB[22][81] ) );
  FA1A S2_21_81 ( .A(\ab[21][81] ), .B(\CARRYB[20][81] ), .CI(\SUMB[20][82] ), 
        .CO(\CARRYB[21][81] ), .S(\SUMB[21][81] ) );
  FA1A S2_20_81 ( .A(\ab[20][81] ), .B(\CARRYB[19][81] ), .CI(\SUMB[19][82] ), 
        .CO(\CARRYB[20][81] ), .S(\SUMB[20][81] ) );
  FA1A S2_19_81 ( .A(\ab[19][81] ), .B(\CARRYB[18][81] ), .CI(\SUMB[18][82] ), 
        .CO(\CARRYB[19][81] ), .S(\SUMB[19][81] ) );
  FA1A S2_18_81 ( .A(\ab[18][81] ), .B(\CARRYB[17][81] ), .CI(\SUMB[17][82] ), 
        .CO(\CARRYB[18][81] ), .S(\SUMB[18][81] ) );
  FA1A S2_17_81 ( .A(\ab[17][81] ), .B(\CARRYB[16][81] ), .CI(\SUMB[16][82] ), 
        .CO(\CARRYB[17][81] ), .S(\SUMB[17][81] ) );
  FA1A S2_16_81 ( .A(\ab[16][81] ), .B(\CARRYB[15][81] ), .CI(\SUMB[15][82] ), 
        .CO(\CARRYB[16][81] ), .S(\SUMB[16][81] ) );
  FA1A S2_15_81 ( .A(\ab[15][81] ), .B(\CARRYB[14][81] ), .CI(\SUMB[14][82] ), 
        .CO(\CARRYB[15][81] ), .S(\SUMB[15][81] ) );
  FA1A S2_28_80 ( .A(\ab[28][80] ), .B(\CARRYB[27][80] ), .CI(\SUMB[27][81] ), 
        .CO(\CARRYB[28][80] ), .S(\SUMB[28][80] ) );
  FA1A S4_82 ( .A(\ab[29][82] ), .B(\CARRYB[28][82] ), .CI(\SUMB[28][83] ), 
        .CO(\CARRYB[29][82] ), .S(\SUMB[29][82] ) );
  FA1A S2_27_80 ( .A(\ab[27][80] ), .B(\CARRYB[26][80] ), .CI(\SUMB[26][81] ), 
        .CO(\CARRYB[27][80] ), .S(\SUMB[27][80] ) );
  FA1A S2_28_82 ( .A(\ab[28][82] ), .B(\CARRYB[27][82] ), .CI(\SUMB[27][83] ), 
        .CO(\CARRYB[28][82] ), .S(\SUMB[28][82] ) );
  FA1A S4_83 ( .A(\ab[29][83] ), .B(\CARRYB[28][83] ), .CI(\SUMB[28][84] ), 
        .CO(\CARRYB[29][83] ), .S(\SUMB[29][83] ) );
  FA1A S2_26_80 ( .A(\ab[26][80] ), .B(\CARRYB[25][80] ), .CI(\SUMB[25][81] ), 
        .CO(\CARRYB[26][80] ), .S(\SUMB[26][80] ) );
  FA1A S2_27_82 ( .A(\ab[27][82] ), .B(\CARRYB[26][82] ), .CI(\SUMB[26][83] ), 
        .CO(\CARRYB[27][82] ), .S(\SUMB[27][82] ) );
  FA1A S2_28_84 ( .A(\ab[28][84] ), .B(\CARRYB[27][84] ), .CI(\SUMB[27][85] ), 
        .CO(\CARRYB[28][84] ), .S(\SUMB[28][84] ) );
  FA1A S2_28_83 ( .A(\ab[28][83] ), .B(\CARRYB[27][83] ), .CI(\SUMB[27][84] ), 
        .CO(\CARRYB[28][83] ), .S(\SUMB[28][83] ) );
  FA1A S2_25_80 ( .A(\ab[25][80] ), .B(\CARRYB[24][80] ), .CI(\SUMB[24][81] ), 
        .CO(\CARRYB[25][80] ), .S(\SUMB[25][80] ) );
  FA1A S2_26_82 ( .A(\ab[26][82] ), .B(\CARRYB[25][82] ), .CI(\SUMB[25][83] ), 
        .CO(\CARRYB[26][82] ), .S(\SUMB[26][82] ) );
  FA1A S2_27_84 ( .A(\ab[27][84] ), .B(\CARRYB[26][84] ), .CI(\SUMB[26][85] ), 
        .CO(\CARRYB[27][84] ), .S(\SUMB[27][84] ) );
  FA1A S2_27_83 ( .A(\ab[27][83] ), .B(\CARRYB[26][83] ), .CI(\SUMB[26][84] ), 
        .CO(\CARRYB[27][83] ), .S(\SUMB[27][83] ) );
  FA1A S2_25_82 ( .A(\ab[25][82] ), .B(\CARRYB[24][82] ), .CI(\SUMB[24][83] ), 
        .CO(\CARRYB[25][82] ), .S(\SUMB[25][82] ) );
  FA1A S2_26_84 ( .A(\ab[26][84] ), .B(\CARRYB[25][84] ), .CI(\SUMB[25][85] ), 
        .CO(\CARRYB[26][84] ), .S(\SUMB[26][84] ) );
  FA1A S2_26_83 ( .A(\ab[26][83] ), .B(\CARRYB[25][83] ), .CI(\SUMB[25][84] ), 
        .CO(\CARRYB[26][83] ), .S(\SUMB[26][83] ) );
  FA1A S2_24_80 ( .A(\ab[24][80] ), .B(\CARRYB[23][80] ), .CI(\SUMB[23][81] ), 
        .CO(\CARRYB[24][80] ), .S(\SUMB[24][80] ) );
  FA1A S2_24_82 ( .A(\ab[24][82] ), .B(\CARRYB[23][82] ), .CI(\SUMB[23][83] ), 
        .CO(\CARRYB[24][82] ), .S(\SUMB[24][82] ) );
  FA1A S2_25_84 ( .A(\ab[25][84] ), .B(\CARRYB[24][84] ), .CI(\SUMB[24][85] ), 
        .CO(\CARRYB[25][84] ), .S(\SUMB[25][84] ) );
  FA1A S2_25_83 ( .A(\ab[25][83] ), .B(\CARRYB[24][83] ), .CI(\SUMB[24][84] ), 
        .CO(\CARRYB[25][83] ), .S(\SUMB[25][83] ) );
  FA1A S2_23_80 ( .A(\ab[23][80] ), .B(\CARRYB[22][80] ), .CI(\SUMB[22][81] ), 
        .CO(\CARRYB[23][80] ), .S(\SUMB[23][80] ) );
  FA1A S2_23_82 ( .A(\ab[23][82] ), .B(\CARRYB[22][82] ), .CI(\SUMB[22][83] ), 
        .CO(\CARRYB[23][82] ), .S(\SUMB[23][82] ) );
  FA1A S2_24_84 ( .A(\ab[24][84] ), .B(\CARRYB[23][84] ), .CI(\SUMB[23][85] ), 
        .CO(\CARRYB[24][84] ), .S(\SUMB[24][84] ) );
  FA1A S2_24_83 ( .A(\ab[24][83] ), .B(\CARRYB[23][83] ), .CI(\SUMB[23][84] ), 
        .CO(\CARRYB[24][83] ), .S(\SUMB[24][83] ) );
  FA1A S2_22_82 ( .A(\ab[22][82] ), .B(\CARRYB[21][82] ), .CI(\SUMB[21][83] ), 
        .CO(\CARRYB[22][82] ), .S(\SUMB[22][82] ) );
  FA1A S2_22_80 ( .A(\ab[22][80] ), .B(\CARRYB[21][80] ), .CI(\SUMB[21][81] ), 
        .CO(\CARRYB[22][80] ), .S(\SUMB[22][80] ) );
  FA1A S2_23_84 ( .A(\ab[23][84] ), .B(\CARRYB[22][84] ), .CI(\SUMB[22][85] ), 
        .CO(\CARRYB[23][84] ), .S(\SUMB[23][84] ) );
  FA1A S2_23_83 ( .A(\ab[23][83] ), .B(\CARRYB[22][83] ), .CI(\SUMB[22][84] ), 
        .CO(\CARRYB[23][83] ), .S(\SUMB[23][83] ) );
  FA1A S2_21_82 ( .A(\ab[21][82] ), .B(\CARRYB[20][82] ), .CI(\SUMB[20][83] ), 
        .CO(\CARRYB[21][82] ), .S(\SUMB[21][82] ) );
  FA1A S2_21_80 ( .A(\ab[21][80] ), .B(\CARRYB[20][80] ), .CI(\SUMB[20][81] ), 
        .CO(\CARRYB[21][80] ), .S(\SUMB[21][80] ) );
  FA1A S2_22_84 ( .A(\ab[22][84] ), .B(\CARRYB[21][84] ), .CI(\SUMB[21][85] ), 
        .CO(\CARRYB[22][84] ), .S(\SUMB[22][84] ) );
  FA1A S2_22_83 ( .A(\ab[22][83] ), .B(\CARRYB[21][83] ), .CI(\SUMB[21][84] ), 
        .CO(\CARRYB[22][83] ), .S(\SUMB[22][83] ) );
  FA1A S2_20_82 ( .A(\ab[20][82] ), .B(\CARRYB[19][82] ), .CI(\SUMB[19][83] ), 
        .CO(\CARRYB[20][82] ), .S(\SUMB[20][82] ) );
  FA1A S2_20_80 ( .A(\ab[20][80] ), .B(\CARRYB[19][80] ), .CI(\SUMB[19][81] ), 
        .CO(\CARRYB[20][80] ), .S(\SUMB[20][80] ) );
  FA1A S2_21_84 ( .A(\ab[21][84] ), .B(\CARRYB[20][84] ), .CI(\SUMB[20][85] ), 
        .CO(\CARRYB[21][84] ), .S(\SUMB[21][84] ) );
  FA1A S2_21_83 ( .A(\ab[21][83] ), .B(\CARRYB[20][83] ), .CI(\SUMB[20][84] ), 
        .CO(\CARRYB[21][83] ), .S(\SUMB[21][83] ) );
  FA1A S2_19_82 ( .A(\ab[19][82] ), .B(\CARRYB[18][82] ), .CI(\SUMB[18][83] ), 
        .CO(\CARRYB[19][82] ), .S(\SUMB[19][82] ) );
  FA1A S2_20_84 ( .A(\ab[20][84] ), .B(\CARRYB[19][84] ), .CI(\SUMB[19][85] ), 
        .CO(\CARRYB[20][84] ), .S(\SUMB[20][84] ) );
  FA1A S2_20_83 ( .A(\ab[20][83] ), .B(\CARRYB[19][83] ), .CI(\SUMB[19][84] ), 
        .CO(\CARRYB[20][83] ), .S(\SUMB[20][83] ) );
  FA1A S2_18_82 ( .A(\ab[18][82] ), .B(\CARRYB[17][82] ), .CI(\SUMB[17][83] ), 
        .CO(\CARRYB[18][82] ), .S(\SUMB[18][82] ) );
  FA1A S2_19_84 ( .A(\ab[19][84] ), .B(\CARRYB[18][84] ), .CI(\SUMB[18][85] ), 
        .CO(\CARRYB[19][84] ), .S(\SUMB[19][84] ) );
  FA1A S2_19_83 ( .A(\ab[19][83] ), .B(\CARRYB[18][83] ), .CI(\SUMB[18][84] ), 
        .CO(\CARRYB[19][83] ), .S(\SUMB[19][83] ) );
  FA1A S2_18_84 ( .A(\ab[18][84] ), .B(\CARRYB[17][84] ), .CI(\SUMB[17][85] ), 
        .CO(\CARRYB[18][84] ), .S(\SUMB[18][84] ) );
  FA1A S2_18_83 ( .A(\ab[18][83] ), .B(\CARRYB[17][83] ), .CI(\SUMB[17][84] ), 
        .CO(\CARRYB[18][83] ), .S(\SUMB[18][83] ) );
  FA1A S2_17_84 ( .A(\ab[17][84] ), .B(\CARRYB[16][84] ), .CI(\SUMB[16][85] ), 
        .CO(\CARRYB[17][84] ), .S(\SUMB[17][84] ) );
  FA1A S2_17_83 ( .A(\ab[17][83] ), .B(\CARRYB[16][83] ), .CI(\SUMB[16][84] ), 
        .CO(\CARRYB[17][83] ), .S(\SUMB[17][83] ) );
  FA1A S2_16_84 ( .A(\ab[16][84] ), .B(\CARRYB[15][84] ), .CI(\SUMB[15][85] ), 
        .CO(\CARRYB[16][84] ), .S(\SUMB[16][84] ) );
  FA1A S2_19_80 ( .A(\ab[19][80] ), .B(\CARRYB[18][80] ), .CI(\SUMB[18][81] ), 
        .CO(\CARRYB[19][80] ), .S(\SUMB[19][80] ) );
  FA1A S2_18_80 ( .A(\ab[18][80] ), .B(\CARRYB[17][80] ), .CI(\SUMB[17][81] ), 
        .CO(\CARRYB[18][80] ), .S(\SUMB[18][80] ) );
  FA1A S2_17_82 ( .A(\ab[17][82] ), .B(\CARRYB[16][82] ), .CI(\SUMB[16][83] ), 
        .CO(\CARRYB[17][82] ), .S(\SUMB[17][82] ) );
  FA1A S2_17_80 ( .A(\ab[17][80] ), .B(\CARRYB[16][80] ), .CI(\SUMB[16][81] ), 
        .CO(\CARRYB[17][80] ), .S(\SUMB[17][80] ) );
  FA1A S2_16_83 ( .A(\ab[16][83] ), .B(\CARRYB[15][83] ), .CI(\SUMB[15][84] ), 
        .CO(\CARRYB[16][83] ), .S(\SUMB[16][83] ) );
  FA1A S2_16_82 ( .A(\ab[16][82] ), .B(\CARRYB[15][82] ), .CI(\SUMB[15][83] ), 
        .CO(\CARRYB[16][82] ), .S(\SUMB[16][82] ) );
  FA1A S2_15_84 ( .A(\ab[15][84] ), .B(\CARRYB[14][84] ), .CI(\SUMB[14][85] ), 
        .CO(\CARRYB[15][84] ), .S(\SUMB[15][84] ) );
  FA1A S2_15_83 ( .A(\ab[15][83] ), .B(\CARRYB[14][83] ), .CI(\SUMB[14][84] ), 
        .CO(\CARRYB[15][83] ), .S(\SUMB[15][83] ) );
  FA1A S2_15_82 ( .A(\ab[15][82] ), .B(\CARRYB[14][82] ), .CI(\SUMB[14][83] ), 
        .CO(\CARRYB[15][82] ), .S(\SUMB[15][82] ) );
  FA1A S2_16_80 ( .A(\ab[16][80] ), .B(\CARRYB[15][80] ), .CI(\SUMB[15][81] ), 
        .CO(\CARRYB[16][80] ), .S(\SUMB[16][80] ) );
  FA1A S2_15_80 ( .A(\ab[15][80] ), .B(\CARRYB[14][80] ), .CI(\SUMB[14][81] ), 
        .CO(\CARRYB[15][80] ), .S(\SUMB[15][80] ) );
  FA1A S4_84 ( .A(\ab[29][84] ), .B(\CARRYB[28][84] ), .CI(\SUMB[28][85] ), 
        .CO(\CARRYB[29][84] ), .S(\SUMB[29][84] ) );
  FA1A S4_73 ( .A(\ab[29][73] ), .B(\CARRYB[28][73] ), .CI(\SUMB[28][74] ), 
        .CO(\CARRYB[29][73] ), .S(\SUMB[29][73] ) );
  FA1A S4_78 ( .A(\ab[29][78] ), .B(\CARRYB[28][78] ), .CI(\SUMB[28][79] ), 
        .CO(\CARRYB[29][78] ), .S(\SUMB[29][78] ) );
  FA1A S4_77 ( .A(\ab[29][77] ), .B(\CARRYB[28][77] ), .CI(\SUMB[28][78] ), 
        .CO(\CARRYB[29][77] ), .S(\SUMB[29][77] ) );
  FA1A S2_28_73 ( .A(\ab[28][73] ), .B(\CARRYB[27][73] ), .CI(\SUMB[27][74] ), 
        .CO(\CARRYB[28][73] ), .S(\SUMB[28][73] ) );
  FA1A S2_28_79 ( .A(\ab[28][79] ), .B(\CARRYB[27][79] ), .CI(\SUMB[27][80] ), 
        .CO(\CARRYB[28][79] ), .S(\SUMB[28][79] ) );
  FA1A S2_28_78 ( .A(\ab[28][78] ), .B(\CARRYB[27][78] ), .CI(\SUMB[27][79] ), 
        .CO(\CARRYB[28][78] ), .S(\SUMB[28][78] ) );
  FA1A S2_28_77 ( .A(\ab[28][77] ), .B(\CARRYB[27][77] ), .CI(\SUMB[27][78] ), 
        .CO(\CARRYB[28][77] ), .S(\SUMB[28][77] ) );
  FA1A S4_75 ( .A(\ab[29][75] ), .B(\CARRYB[28][75] ), .CI(\SUMB[28][76] ), 
        .CO(\CARRYB[29][75] ), .S(\SUMB[29][75] ) );
  FA1A S4_71 ( .A(\ab[29][71] ), .B(\CARRYB[28][71] ), .CI(\SUMB[28][72] ), 
        .CO(\CARRYB[29][71] ), .S(\SUMB[29][71] ) );
  FA1A S2_27_79 ( .A(\ab[27][79] ), .B(\CARRYB[26][79] ), .CI(\SUMB[26][80] ), 
        .CO(\CARRYB[27][79] ), .S(\SUMB[27][79] ) );
  FA1A S2_27_78 ( .A(\ab[27][78] ), .B(\CARRYB[26][78] ), .CI(\SUMB[26][79] ), 
        .CO(\CARRYB[27][78] ), .S(\SUMB[27][78] ) );
  FA1A S2_28_76 ( .A(\ab[28][76] ), .B(\CARRYB[27][76] ), .CI(\SUMB[27][77] ), 
        .CO(\CARRYB[28][76] ), .S(\SUMB[28][76] ) );
  FA1A S2_28_75 ( .A(\ab[28][75] ), .B(\CARRYB[27][75] ), .CI(\SUMB[27][76] ), 
        .CO(\CARRYB[28][75] ), .S(\SUMB[28][75] ) );
  FA1A S2_28_74 ( .A(\ab[28][74] ), .B(\CARRYB[27][74] ), .CI(\SUMB[27][75] ), 
        .CO(\CARRYB[28][74] ), .S(\SUMB[28][74] ) );
  FA1A S2_28_72 ( .A(\ab[28][72] ), .B(\CARRYB[27][72] ), .CI(\SUMB[27][73] ), 
        .CO(\CARRYB[28][72] ), .S(\SUMB[28][72] ) );
  FA1A S4_69 ( .A(\ab[29][69] ), .B(\CARRYB[28][69] ), .CI(\SUMB[28][70] ), 
        .CO(\CARRYB[29][69] ), .S(\SUMB[29][69] ) );
  FA1A S2_26_79 ( .A(\ab[26][79] ), .B(\CARRYB[25][79] ), .CI(\SUMB[25][80] ), 
        .CO(\CARRYB[26][79] ), .S(\SUMB[26][79] ) );
  FA1A S2_27_77 ( .A(\ab[27][77] ), .B(\CARRYB[26][77] ), .CI(\SUMB[26][78] ), 
        .CO(\CARRYB[27][77] ), .S(\SUMB[27][77] ) );
  FA1A S2_27_76 ( .A(\ab[27][76] ), .B(\CARRYB[26][76] ), .CI(\SUMB[26][77] ), 
        .CO(\CARRYB[27][76] ), .S(\SUMB[27][76] ) );
  FA1A S2_27_75 ( .A(\ab[27][75] ), .B(\CARRYB[26][75] ), .CI(\SUMB[26][76] ), 
        .CO(\CARRYB[27][75] ), .S(\SUMB[27][75] ) );
  FA1A S2_27_74 ( .A(\ab[27][74] ), .B(\CARRYB[26][74] ), .CI(\SUMB[26][75] ), 
        .CO(\CARRYB[27][74] ), .S(\SUMB[27][74] ) );
  FA1A S2_27_73 ( .A(\ab[27][73] ), .B(\CARRYB[26][73] ), .CI(\SUMB[26][74] ), 
        .CO(\CARRYB[27][73] ), .S(\SUMB[27][73] ) );
  FA1A S2_28_69 ( .A(\ab[28][69] ), .B(\CARRYB[27][69] ), .CI(\SUMB[27][70] ), 
        .CO(\CARRYB[28][69] ), .S(\SUMB[28][69] ) );
  FA1A S2_26_78 ( .A(\ab[26][78] ), .B(\CARRYB[25][78] ), .CI(\SUMB[25][79] ), 
        .CO(\CARRYB[26][78] ), .S(\SUMB[26][78] ) );
  FA1A S2_26_77 ( .A(\ab[26][77] ), .B(\CARRYB[25][77] ), .CI(\SUMB[25][78] ), 
        .CO(\CARRYB[26][77] ), .S(\SUMB[26][77] ) );
  FA1A S2_26_76 ( .A(\ab[26][76] ), .B(\CARRYB[25][76] ), .CI(\SUMB[25][77] ), 
        .CO(\CARRYB[26][76] ), .S(\SUMB[26][76] ) );
  FA1A S2_26_75 ( .A(\ab[26][75] ), .B(\CARRYB[25][75] ), .CI(\SUMB[25][76] ), 
        .CO(\CARRYB[26][75] ), .S(\SUMB[26][75] ) );
  FA1A S2_26_74 ( .A(\ab[26][74] ), .B(\CARRYB[25][74] ), .CI(\SUMB[25][75] ), 
        .CO(\CARRYB[26][74] ), .S(\SUMB[26][74] ) );
  FA1A S2_25_79 ( .A(\ab[25][79] ), .B(\CARRYB[24][79] ), .CI(\SUMB[24][80] ), 
        .CO(\CARRYB[25][79] ), .S(\SUMB[25][79] ) );
  FA1A S2_25_78 ( .A(\ab[25][78] ), .B(\CARRYB[24][78] ), .CI(\SUMB[24][79] ), 
        .CO(\CARRYB[25][78] ), .S(\SUMB[25][78] ) );
  FA1A S2_25_77 ( .A(\ab[25][77] ), .B(\CARRYB[24][77] ), .CI(\SUMB[24][78] ), 
        .CO(\CARRYB[25][77] ), .S(\SUMB[25][77] ) );
  FA1A S2_25_76 ( .A(\ab[25][76] ), .B(\CARRYB[24][76] ), .CI(\SUMB[24][77] ), 
        .CO(\CARRYB[25][76] ), .S(\SUMB[25][76] ) );
  FA1A S2_25_75 ( .A(\ab[25][75] ), .B(\CARRYB[24][75] ), .CI(\SUMB[24][76] ), 
        .CO(\CARRYB[25][75] ), .S(\SUMB[25][75] ) );
  FA1A S2_24_79 ( .A(\ab[24][79] ), .B(\CARRYB[23][79] ), .CI(\SUMB[23][80] ), 
        .CO(\CARRYB[24][79] ), .S(\SUMB[24][79] ) );
  FA1A S2_24_78 ( .A(\ab[24][78] ), .B(\CARRYB[23][78] ), .CI(\SUMB[23][79] ), 
        .CO(\CARRYB[24][78] ), .S(\SUMB[24][78] ) );
  FA1A S2_24_77 ( .A(\ab[24][77] ), .B(\CARRYB[23][77] ), .CI(\SUMB[23][78] ), 
        .CO(\CARRYB[24][77] ), .S(\SUMB[24][77] ) );
  FA1A S2_24_76 ( .A(\ab[24][76] ), .B(\CARRYB[23][76] ), .CI(\SUMB[23][77] ), 
        .CO(\CARRYB[24][76] ), .S(\SUMB[24][76] ) );
  FA1A S4_57 ( .A(\ab[29][57] ), .B(\CARRYB[28][57] ), .CI(\SUMB[28][58] ), 
        .CO(\CARRYB[29][57] ), .S(\SUMB[29][57] ) );
  FA1A S2_23_79 ( .A(\ab[23][79] ), .B(\CARRYB[22][79] ), .CI(\SUMB[22][80] ), 
        .CO(\CARRYB[23][79] ), .S(\SUMB[23][79] ) );
  FA1A S2_23_78 ( .A(\ab[23][78] ), .B(\CARRYB[22][78] ), .CI(\SUMB[22][79] ), 
        .CO(\CARRYB[23][78] ), .S(\SUMB[23][78] ) );
  FA1A S2_23_77 ( .A(\ab[23][77] ), .B(\CARRYB[22][77] ), .CI(\SUMB[22][78] ), 
        .CO(\CARRYB[23][77] ), .S(\SUMB[23][77] ) );
  FA1A S2_28_57 ( .A(\ab[28][57] ), .B(\CARRYB[27][57] ), .CI(\SUMB[27][58] ), 
        .CO(\CARRYB[28][57] ), .S(\SUMB[28][57] ) );
  FA1A S2_22_79 ( .A(\ab[22][79] ), .B(\CARRYB[21][79] ), .CI(\SUMB[21][80] ), 
        .CO(\CARRYB[22][79] ), .S(\SUMB[22][79] ) );
  FA1A S2_22_78 ( .A(\ab[22][78] ), .B(\CARRYB[21][78] ), .CI(\SUMB[21][79] ), 
        .CO(\CARRYB[22][78] ), .S(\SUMB[22][78] ) );
  FA1A S2_28_71 ( .A(\ab[28][71] ), .B(\CARRYB[27][71] ), .CI(\SUMB[27][72] ), 
        .CO(\CARRYB[28][71] ), .S(\SUMB[28][71] ) );
  FA1A S2_28_70 ( .A(\ab[28][70] ), .B(\CARRYB[27][70] ), .CI(\SUMB[27][71] ), 
        .CO(\CARRYB[28][70] ), .S(\SUMB[28][70] ) );
  FA1A S2_21_79 ( .A(\ab[21][79] ), .B(\CARRYB[20][79] ), .CI(\SUMB[20][80] ), 
        .CO(\CARRYB[21][79] ), .S(\SUMB[21][79] ) );
  FA1A S2_27_72 ( .A(\ab[27][72] ), .B(\CARRYB[26][72] ), .CI(\SUMB[26][73] ), 
        .CO(\CARRYB[27][72] ), .S(\SUMB[27][72] ) );
  FA1A S2_27_71 ( .A(\ab[27][71] ), .B(\CARRYB[26][71] ), .CI(\SUMB[26][72] ), 
        .CO(\CARRYB[27][71] ), .S(\SUMB[27][71] ) );
  FA1A S2_27_70 ( .A(\ab[27][70] ), .B(\CARRYB[26][70] ), .CI(\SUMB[26][71] ), 
        .CO(\CARRYB[27][70] ), .S(\SUMB[27][70] ) );
  FA1A S2_27_57 ( .A(\ab[27][57] ), .B(\CARRYB[26][57] ), .CI(\SUMB[26][58] ), 
        .CO(\CARRYB[27][57] ), .S(\SUMB[27][57] ) );
  FA1A S2_26_73 ( .A(\ab[26][73] ), .B(\CARRYB[25][73] ), .CI(\SUMB[25][74] ), 
        .CO(\CARRYB[26][73] ), .S(\SUMB[26][73] ) );
  FA1A S2_26_72 ( .A(\ab[26][72] ), .B(\CARRYB[25][72] ), .CI(\SUMB[25][73] ), 
        .CO(\CARRYB[26][72] ), .S(\SUMB[26][72] ) );
  FA1A S2_26_71 ( .A(\ab[26][71] ), .B(\CARRYB[25][71] ), .CI(\SUMB[25][72] ), 
        .CO(\CARRYB[26][71] ), .S(\SUMB[26][71] ) );
  FA1A S2_25_74 ( .A(\ab[25][74] ), .B(\CARRYB[24][74] ), .CI(\SUMB[24][75] ), 
        .CO(\CARRYB[25][74] ), .S(\SUMB[25][74] ) );
  FA1A S2_25_73 ( .A(\ab[25][73] ), .B(\CARRYB[24][73] ), .CI(\SUMB[24][74] ), 
        .CO(\CARRYB[25][73] ), .S(\SUMB[25][73] ) );
  FA1A S2_25_72 ( .A(\ab[25][72] ), .B(\CARRYB[24][72] ), .CI(\SUMB[24][73] ), 
        .CO(\CARRYB[25][72] ), .S(\SUMB[25][72] ) );
  FA1A S2_27_69 ( .A(\ab[27][69] ), .B(\CARRYB[26][69] ), .CI(\SUMB[26][70] ), 
        .CO(\CARRYB[27][69] ), .S(\SUMB[27][69] ) );
  FA1A S2_26_57 ( .A(\ab[26][57] ), .B(\CARRYB[25][57] ), .CI(\SUMB[25][58] ), 
        .CO(\CARRYB[26][57] ), .S(\SUMB[26][57] ) );
  FA1A S2_24_75 ( .A(\ab[24][75] ), .B(\CARRYB[23][75] ), .CI(\SUMB[23][76] ), 
        .CO(\CARRYB[24][75] ), .S(\SUMB[24][75] ) );
  FA1A S2_24_74 ( .A(\ab[24][74] ), .B(\CARRYB[23][74] ), .CI(\SUMB[23][75] ), 
        .CO(\CARRYB[24][74] ), .S(\SUMB[24][74] ) );
  FA1A S2_24_73 ( .A(\ab[24][73] ), .B(\CARRYB[23][73] ), .CI(\SUMB[23][74] ), 
        .CO(\CARRYB[24][73] ), .S(\SUMB[24][73] ) );
  FA1A S2_26_69 ( .A(\ab[26][69] ), .B(\CARRYB[25][69] ), .CI(\SUMB[25][70] ), 
        .CO(\CARRYB[26][69] ), .S(\SUMB[26][69] ) );
  FA1A S2_26_70 ( .A(\ab[26][70] ), .B(\CARRYB[25][70] ), .CI(\SUMB[25][71] ), 
        .CO(\CARRYB[26][70] ), .S(\SUMB[26][70] ) );
  FA1A S2_25_57 ( .A(\ab[25][57] ), .B(\CARRYB[24][57] ), .CI(\SUMB[24][58] ), 
        .CO(\CARRYB[25][57] ), .S(\SUMB[25][57] ) );
  FA1A S2_23_76 ( .A(\ab[23][76] ), .B(\CARRYB[22][76] ), .CI(\SUMB[22][77] ), 
        .CO(\CARRYB[23][76] ), .S(\SUMB[23][76] ) );
  FA1A S2_23_75 ( .A(\ab[23][75] ), .B(\CARRYB[22][75] ), .CI(\SUMB[22][76] ), 
        .CO(\CARRYB[23][75] ), .S(\SUMB[23][75] ) );
  FA1A S2_23_74 ( .A(\ab[23][74] ), .B(\CARRYB[22][74] ), .CI(\SUMB[22][75] ), 
        .CO(\CARRYB[23][74] ), .S(\SUMB[23][74] ) );
  FA1A S2_25_69 ( .A(\ab[25][69] ), .B(\CARRYB[24][69] ), .CI(\SUMB[24][70] ), 
        .CO(\CARRYB[25][69] ), .S(\SUMB[25][69] ) );
  FA1A S2_25_70 ( .A(\ab[25][70] ), .B(\CARRYB[24][70] ), .CI(\SUMB[24][71] ), 
        .CO(\CARRYB[25][70] ), .S(\SUMB[25][70] ) );
  FA1A S2_25_71 ( .A(\ab[25][71] ), .B(\CARRYB[24][71] ), .CI(\SUMB[24][72] ), 
        .CO(\CARRYB[25][71] ), .S(\SUMB[25][71] ) );
  FA1A S2_24_57 ( .A(\ab[24][57] ), .B(\CARRYB[23][57] ), .CI(\SUMB[23][58] ), 
        .CO(\CARRYB[24][57] ), .S(\SUMB[24][57] ) );
  FA1A S2_22_77 ( .A(\ab[22][77] ), .B(\CARRYB[21][77] ), .CI(\SUMB[21][78] ), 
        .CO(\CARRYB[22][77] ), .S(\SUMB[22][77] ) );
  FA1A S2_22_76 ( .A(\ab[22][76] ), .B(\CARRYB[21][76] ), .CI(\SUMB[21][77] ), 
        .CO(\CARRYB[22][76] ), .S(\SUMB[22][76] ) );
  FA1A S2_22_75 ( .A(\ab[22][75] ), .B(\CARRYB[21][75] ), .CI(\SUMB[21][76] ), 
        .CO(\CARRYB[22][75] ), .S(\SUMB[22][75] ) );
  FA1A S2_24_69 ( .A(\ab[24][69] ), .B(\CARRYB[23][69] ), .CI(\SUMB[23][70] ), 
        .CO(\CARRYB[24][69] ), .S(\SUMB[24][69] ) );
  FA1A S2_24_70 ( .A(\ab[24][70] ), .B(\CARRYB[23][70] ), .CI(\SUMB[23][71] ), 
        .CO(\CARRYB[24][70] ), .S(\SUMB[24][70] ) );
  FA1A S2_24_71 ( .A(\ab[24][71] ), .B(\CARRYB[23][71] ), .CI(\SUMB[23][72] ), 
        .CO(\CARRYB[24][71] ), .S(\SUMB[24][71] ) );
  FA1A S2_24_72 ( .A(\ab[24][72] ), .B(\CARRYB[23][72] ), .CI(\SUMB[23][73] ), 
        .CO(\CARRYB[24][72] ), .S(\SUMB[24][72] ) );
  FA1A S2_21_78 ( .A(\ab[21][78] ), .B(\CARRYB[20][78] ), .CI(\SUMB[20][79] ), 
        .CO(\CARRYB[21][78] ), .S(\SUMB[21][78] ) );
  FA1A S2_21_77 ( .A(\ab[21][77] ), .B(\CARRYB[20][77] ), .CI(\SUMB[20][78] ), 
        .CO(\CARRYB[21][77] ), .S(\SUMB[21][77] ) );
  FA1A S2_21_76 ( .A(\ab[21][76] ), .B(\CARRYB[20][76] ), .CI(\SUMB[20][77] ), 
        .CO(\CARRYB[21][76] ), .S(\SUMB[21][76] ) );
  FA1A S2_23_69 ( .A(\ab[23][69] ), .B(\CARRYB[22][69] ), .CI(\SUMB[22][70] ), 
        .CO(\CARRYB[23][69] ), .S(\SUMB[23][69] ) );
  FA1A S2_23_70 ( .A(\ab[23][70] ), .B(\CARRYB[22][70] ), .CI(\SUMB[22][71] ), 
        .CO(\CARRYB[23][70] ), .S(\SUMB[23][70] ) );
  FA1A S2_23_71 ( .A(\ab[23][71] ), .B(\CARRYB[22][71] ), .CI(\SUMB[22][72] ), 
        .CO(\CARRYB[23][71] ), .S(\SUMB[23][71] ) );
  FA1A S2_23_72 ( .A(\ab[23][72] ), .B(\CARRYB[22][72] ), .CI(\SUMB[22][73] ), 
        .CO(\CARRYB[23][72] ), .S(\SUMB[23][72] ) );
  FA1A S2_23_73 ( .A(\ab[23][73] ), .B(\CARRYB[22][73] ), .CI(\SUMB[22][74] ), 
        .CO(\CARRYB[23][73] ), .S(\SUMB[23][73] ) );
  FA1A S2_23_57 ( .A(\ab[23][57] ), .B(\CARRYB[22][57] ), .CI(\SUMB[22][58] ), 
        .CO(\CARRYB[23][57] ), .S(\SUMB[23][57] ) );
  FA1A S2_20_79 ( .A(\ab[20][79] ), .B(\CARRYB[19][79] ), .CI(\SUMB[19][80] ), 
        .CO(\CARRYB[20][79] ), .S(\SUMB[20][79] ) );
  FA1A S2_20_78 ( .A(\ab[20][78] ), .B(\CARRYB[19][78] ), .CI(\SUMB[19][79] ), 
        .CO(\CARRYB[20][78] ), .S(\SUMB[20][78] ) );
  FA1A S2_20_77 ( .A(\ab[20][77] ), .B(\CARRYB[19][77] ), .CI(\SUMB[19][78] ), 
        .CO(\CARRYB[20][77] ), .S(\SUMB[20][77] ) );
  FA1A S2_22_70 ( .A(\ab[22][70] ), .B(\CARRYB[21][70] ), .CI(\SUMB[21][71] ), 
        .CO(\CARRYB[22][70] ), .S(\SUMB[22][70] ) );
  FA1A S2_22_71 ( .A(\ab[22][71] ), .B(\CARRYB[21][71] ), .CI(\SUMB[21][72] ), 
        .CO(\CARRYB[22][71] ), .S(\SUMB[22][71] ) );
  FA1A S2_22_72 ( .A(\ab[22][72] ), .B(\CARRYB[21][72] ), .CI(\SUMB[21][73] ), 
        .CO(\CARRYB[22][72] ), .S(\SUMB[22][72] ) );
  FA1A S2_22_73 ( .A(\ab[22][73] ), .B(\CARRYB[21][73] ), .CI(\SUMB[21][74] ), 
        .CO(\CARRYB[22][73] ), .S(\SUMB[22][73] ) );
  FA1A S2_22_74 ( .A(\ab[22][74] ), .B(\CARRYB[21][74] ), .CI(\SUMB[21][75] ), 
        .CO(\CARRYB[22][74] ), .S(\SUMB[22][74] ) );
  FA1A S2_19_79 ( .A(\ab[19][79] ), .B(\CARRYB[18][79] ), .CI(\SUMB[18][80] ), 
        .CO(\CARRYB[19][79] ), .S(\SUMB[19][79] ) );
  FA1A S2_19_78 ( .A(\ab[19][78] ), .B(\CARRYB[18][78] ), .CI(\SUMB[18][79] ), 
        .CO(\CARRYB[19][78] ), .S(\SUMB[19][78] ) );
  FA1A S2_21_71 ( .A(\ab[21][71] ), .B(\CARRYB[20][71] ), .CI(\SUMB[20][72] ), 
        .CO(\CARRYB[21][71] ), .S(\SUMB[21][71] ) );
  FA1A S2_21_72 ( .A(\ab[21][72] ), .B(\CARRYB[20][72] ), .CI(\SUMB[20][73] ), 
        .CO(\CARRYB[21][72] ), .S(\SUMB[21][72] ) );
  FA1A S2_21_73 ( .A(\ab[21][73] ), .B(\CARRYB[20][73] ), .CI(\SUMB[20][74] ), 
        .CO(\CARRYB[21][73] ), .S(\SUMB[21][73] ) );
  FA1A S2_21_74 ( .A(\ab[21][74] ), .B(\CARRYB[20][74] ), .CI(\SUMB[20][75] ), 
        .CO(\CARRYB[21][74] ), .S(\SUMB[21][74] ) );
  FA1A S2_21_75 ( .A(\ab[21][75] ), .B(\CARRYB[20][75] ), .CI(\SUMB[20][76] ), 
        .CO(\CARRYB[21][75] ), .S(\SUMB[21][75] ) );
  FA1A S2_18_79 ( .A(\ab[18][79] ), .B(\CARRYB[17][79] ), .CI(\SUMB[17][80] ), 
        .CO(\CARRYB[18][79] ), .S(\SUMB[18][79] ) );
  FA1A S2_20_72 ( .A(\ab[20][72] ), .B(\CARRYB[19][72] ), .CI(\SUMB[19][73] ), 
        .CO(\CARRYB[20][72] ), .S(\SUMB[20][72] ) );
  FA1A S2_20_73 ( .A(\ab[20][73] ), .B(\CARRYB[19][73] ), .CI(\SUMB[19][74] ), 
        .CO(\CARRYB[20][73] ), .S(\SUMB[20][73] ) );
  FA1A S2_20_74 ( .A(\ab[20][74] ), .B(\CARRYB[19][74] ), .CI(\SUMB[19][75] ), 
        .CO(\CARRYB[20][74] ), .S(\SUMB[20][74] ) );
  FA1A S2_20_75 ( .A(\ab[20][75] ), .B(\CARRYB[19][75] ), .CI(\SUMB[19][76] ), 
        .CO(\CARRYB[20][75] ), .S(\SUMB[20][75] ) );
  FA1A S2_20_76 ( .A(\ab[20][76] ), .B(\CARRYB[19][76] ), .CI(\SUMB[19][77] ), 
        .CO(\CARRYB[20][76] ), .S(\SUMB[20][76] ) );
  FA1A S2_22_69 ( .A(\ab[22][69] ), .B(\CARRYB[21][69] ), .CI(\SUMB[21][70] ), 
        .CO(\CARRYB[22][69] ), .S(\SUMB[22][69] ) );
  FA1A S2_22_57 ( .A(\ab[22][57] ), .B(\CARRYB[21][57] ), .CI(\SUMB[21][58] ), 
        .CO(\CARRYB[22][57] ), .S(\SUMB[22][57] ) );
  FA1A S2_19_73 ( .A(\ab[19][73] ), .B(\CARRYB[18][73] ), .CI(\SUMB[18][74] ), 
        .CO(\CARRYB[19][73] ), .S(\SUMB[19][73] ) );
  FA1A S2_19_74 ( .A(\ab[19][74] ), .B(\CARRYB[18][74] ), .CI(\SUMB[18][75] ), 
        .CO(\CARRYB[19][74] ), .S(\SUMB[19][74] ) );
  FA1A S2_19_75 ( .A(\ab[19][75] ), .B(\CARRYB[18][75] ), .CI(\SUMB[18][76] ), 
        .CO(\CARRYB[19][75] ), .S(\SUMB[19][75] ) );
  FA1A S2_19_76 ( .A(\ab[19][76] ), .B(\CARRYB[18][76] ), .CI(\SUMB[18][77] ), 
        .CO(\CARRYB[19][76] ), .S(\SUMB[19][76] ) );
  FA1A S2_19_77 ( .A(\ab[19][77] ), .B(\CARRYB[18][77] ), .CI(\SUMB[18][78] ), 
        .CO(\CARRYB[19][77] ), .S(\SUMB[19][77] ) );
  FA1A S2_21_69 ( .A(\ab[21][69] ), .B(\CARRYB[20][69] ), .CI(\SUMB[20][70] ), 
        .CO(\CARRYB[21][69] ), .S(\SUMB[21][69] ) );
  FA1A S2_21_70 ( .A(\ab[21][70] ), .B(\CARRYB[20][70] ), .CI(\SUMB[20][71] ), 
        .CO(\CARRYB[21][70] ), .S(\SUMB[21][70] ) );
  FA1A S2_21_57 ( .A(\ab[21][57] ), .B(\CARRYB[20][57] ), .CI(\SUMB[20][58] ), 
        .CO(\CARRYB[21][57] ), .S(\SUMB[21][57] ) );
  FA1A S2_18_74 ( .A(\ab[18][74] ), .B(\CARRYB[17][74] ), .CI(\SUMB[17][75] ), 
        .CO(\CARRYB[18][74] ), .S(\SUMB[18][74] ) );
  FA1A S2_18_75 ( .A(\ab[18][75] ), .B(\CARRYB[17][75] ), .CI(\SUMB[17][76] ), 
        .CO(\CARRYB[18][75] ), .S(\SUMB[18][75] ) );
  FA1A S2_18_76 ( .A(\ab[18][76] ), .B(\CARRYB[17][76] ), .CI(\SUMB[17][77] ), 
        .CO(\CARRYB[18][76] ), .S(\SUMB[18][76] ) );
  FA1A S2_18_77 ( .A(\ab[18][77] ), .B(\CARRYB[17][77] ), .CI(\SUMB[17][78] ), 
        .CO(\CARRYB[18][77] ), .S(\SUMB[18][77] ) );
  FA1A S2_18_78 ( .A(\ab[18][78] ), .B(\CARRYB[17][78] ), .CI(\SUMB[17][79] ), 
        .CO(\CARRYB[18][78] ), .S(\SUMB[18][78] ) );
  FA1A S2_20_69 ( .A(\ab[20][69] ), .B(\CARRYB[19][69] ), .CI(\SUMB[19][70] ), 
        .CO(\CARRYB[20][69] ), .S(\SUMB[20][69] ) );
  FA1A S2_20_70 ( .A(\ab[20][70] ), .B(\CARRYB[19][70] ), .CI(\SUMB[19][71] ), 
        .CO(\CARRYB[20][70] ), .S(\SUMB[20][70] ) );
  FA1A S2_20_71 ( .A(\ab[20][71] ), .B(\CARRYB[19][71] ), .CI(\SUMB[19][72] ), 
        .CO(\CARRYB[20][71] ), .S(\SUMB[20][71] ) );
  FA1A S2_20_57 ( .A(\ab[20][57] ), .B(\CARRYB[19][57] ), .CI(\SUMB[19][58] ), 
        .CO(\CARRYB[20][57] ), .S(\SUMB[20][57] ) );
  FA1A S2_17_75 ( .A(\ab[17][75] ), .B(\CARRYB[16][75] ), .CI(\SUMB[16][76] ), 
        .CO(\CARRYB[17][75] ), .S(\SUMB[17][75] ) );
  FA1A S2_17_76 ( .A(\ab[17][76] ), .B(\CARRYB[16][76] ), .CI(\SUMB[16][77] ), 
        .CO(\CARRYB[17][76] ), .S(\SUMB[17][76] ) );
  FA1A S2_17_77 ( .A(\ab[17][77] ), .B(\CARRYB[16][77] ), .CI(\SUMB[16][78] ), 
        .CO(\CARRYB[17][77] ), .S(\SUMB[17][77] ) );
  FA1A S2_17_78 ( .A(\ab[17][78] ), .B(\CARRYB[16][78] ), .CI(\SUMB[16][79] ), 
        .CO(\CARRYB[17][78] ), .S(\SUMB[17][78] ) );
  FA1A S2_17_79 ( .A(\ab[17][79] ), .B(\CARRYB[16][79] ), .CI(\SUMB[16][80] ), 
        .CO(\CARRYB[17][79] ), .S(\SUMB[17][79] ) );
  FA1A S2_19_70 ( .A(\ab[19][70] ), .B(\CARRYB[18][70] ), .CI(\SUMB[18][71] ), 
        .CO(\CARRYB[19][70] ), .S(\SUMB[19][70] ) );
  FA1A S2_19_69 ( .A(\ab[19][69] ), .B(\CARRYB[18][69] ), .CI(\SUMB[18][70] ), 
        .CO(\CARRYB[19][69] ), .S(\SUMB[19][69] ) );
  FA1A S2_19_71 ( .A(\ab[19][71] ), .B(\CARRYB[18][71] ), .CI(\SUMB[18][72] ), 
        .CO(\CARRYB[19][71] ), .S(\SUMB[19][71] ) );
  FA1A S2_19_72 ( .A(\ab[19][72] ), .B(\CARRYB[18][72] ), .CI(\SUMB[18][73] ), 
        .CO(\CARRYB[19][72] ), .S(\SUMB[19][72] ) );
  FA1A S2_19_57 ( .A(\ab[19][57] ), .B(\CARRYB[18][57] ), .CI(\SUMB[18][58] ), 
        .CO(\CARRYB[19][57] ), .S(\SUMB[19][57] ) );
  FA1A S2_16_76 ( .A(\ab[16][76] ), .B(\CARRYB[15][76] ), .CI(\SUMB[15][77] ), 
        .CO(\CARRYB[16][76] ), .S(\SUMB[16][76] ) );
  FA1A S2_16_77 ( .A(\ab[16][77] ), .B(\CARRYB[15][77] ), .CI(\SUMB[15][78] ), 
        .CO(\CARRYB[16][77] ), .S(\SUMB[16][77] ) );
  FA1A S2_16_78 ( .A(\ab[16][78] ), .B(\CARRYB[15][78] ), .CI(\SUMB[15][79] ), 
        .CO(\CARRYB[16][78] ), .S(\SUMB[16][78] ) );
  FA1A S2_16_79 ( .A(\ab[16][79] ), .B(\CARRYB[15][79] ), .CI(\SUMB[15][80] ), 
        .CO(\CARRYB[16][79] ), .S(\SUMB[16][79] ) );
  FA1A S2_18_71 ( .A(\ab[18][71] ), .B(\CARRYB[17][71] ), .CI(\SUMB[17][72] ), 
        .CO(\CARRYB[18][71] ), .S(\SUMB[18][71] ) );
  FA1A S2_18_70 ( .A(\ab[18][70] ), .B(\CARRYB[17][70] ), .CI(\SUMB[17][71] ), 
        .CO(\CARRYB[18][70] ), .S(\SUMB[18][70] ) );
  FA1A S2_18_69 ( .A(\ab[18][69] ), .B(\CARRYB[17][69] ), .CI(\SUMB[17][70] ), 
        .CO(\CARRYB[18][69] ), .S(\SUMB[18][69] ) );
  FA1A S2_18_72 ( .A(\ab[18][72] ), .B(\CARRYB[17][72] ), .CI(\SUMB[17][73] ), 
        .CO(\CARRYB[18][72] ), .S(\SUMB[18][72] ) );
  FA1A S2_18_73 ( .A(\ab[18][73] ), .B(\CARRYB[17][73] ), .CI(\SUMB[17][74] ), 
        .CO(\CARRYB[18][73] ), .S(\SUMB[18][73] ) );
  FA1A S2_18_57 ( .A(\ab[18][57] ), .B(\CARRYB[17][57] ), .CI(\SUMB[17][58] ), 
        .CO(\CARRYB[18][57] ), .S(\SUMB[18][57] ) );
  FA1A S2_15_77 ( .A(\ab[15][77] ), .B(\CARRYB[14][77] ), .CI(\SUMB[14][78] ), 
        .CO(\CARRYB[15][77] ), .S(\SUMB[15][77] ) );
  FA1A S2_15_78 ( .A(\ab[15][78] ), .B(\CARRYB[14][78] ), .CI(\SUMB[14][79] ), 
        .CO(\CARRYB[15][78] ), .S(\SUMB[15][78] ) );
  FA1A S2_15_79 ( .A(\ab[15][79] ), .B(\CARRYB[14][79] ), .CI(\SUMB[14][80] ), 
        .CO(\CARRYB[15][79] ), .S(\SUMB[15][79] ) );
  FA1A S2_17_72 ( .A(\ab[17][72] ), .B(\CARRYB[16][72] ), .CI(\SUMB[16][73] ), 
        .CO(\CARRYB[17][72] ), .S(\SUMB[17][72] ) );
  FA1A S2_17_71 ( .A(\ab[17][71] ), .B(\CARRYB[16][71] ), .CI(\SUMB[16][72] ), 
        .CO(\CARRYB[17][71] ), .S(\SUMB[17][71] ) );
  FA1A S2_17_70 ( .A(\ab[17][70] ), .B(\CARRYB[16][70] ), .CI(\SUMB[16][71] ), 
        .CO(\CARRYB[17][70] ), .S(\SUMB[17][70] ) );
  FA1A S2_17_69 ( .A(\ab[17][69] ), .B(\CARRYB[16][69] ), .CI(\SUMB[16][70] ), 
        .CO(\CARRYB[17][69] ), .S(\SUMB[17][69] ) );
  FA1A S2_17_73 ( .A(\ab[17][73] ), .B(\CARRYB[16][73] ), .CI(\SUMB[16][74] ), 
        .CO(\CARRYB[17][73] ), .S(\SUMB[17][73] ) );
  FA1A S2_17_74 ( .A(\ab[17][74] ), .B(\CARRYB[16][74] ), .CI(\SUMB[16][75] ), 
        .CO(\CARRYB[17][74] ), .S(\SUMB[17][74] ) );
  FA1A S2_17_57 ( .A(\ab[17][57] ), .B(\CARRYB[16][57] ), .CI(\SUMB[16][58] ), 
        .CO(\CARRYB[17][57] ), .S(\SUMB[17][57] ) );
  FA1A S2_16_73 ( .A(\ab[16][73] ), .B(\CARRYB[15][73] ), .CI(\SUMB[15][74] ), 
        .CO(\CARRYB[16][73] ), .S(\SUMB[16][73] ) );
  FA1A S2_16_72 ( .A(\ab[16][72] ), .B(\CARRYB[15][72] ), .CI(\SUMB[15][73] ), 
        .CO(\CARRYB[16][72] ), .S(\SUMB[16][72] ) );
  FA1A S2_16_71 ( .A(\ab[16][71] ), .B(\CARRYB[15][71] ), .CI(\SUMB[15][72] ), 
        .CO(\CARRYB[16][71] ), .S(\SUMB[16][71] ) );
  FA1A S2_16_70 ( .A(\ab[16][70] ), .B(\CARRYB[15][70] ), .CI(\SUMB[15][71] ), 
        .CO(\CARRYB[16][70] ), .S(\SUMB[16][70] ) );
  FA1A S2_16_69 ( .A(\ab[16][69] ), .B(\CARRYB[15][69] ), .CI(\SUMB[15][70] ), 
        .CO(\CARRYB[16][69] ), .S(\SUMB[16][69] ) );
  FA1A S2_16_74 ( .A(\ab[16][74] ), .B(\CARRYB[15][74] ), .CI(\SUMB[15][75] ), 
        .CO(\CARRYB[16][74] ), .S(\SUMB[16][74] ) );
  FA1A S2_16_75 ( .A(\ab[16][75] ), .B(\CARRYB[15][75] ), .CI(\SUMB[15][76] ), 
        .CO(\CARRYB[16][75] ), .S(\SUMB[16][75] ) );
  FA1A S2_16_57 ( .A(\ab[16][57] ), .B(\CARRYB[15][57] ), .CI(\SUMB[15][58] ), 
        .CO(\CARRYB[16][57] ), .S(\SUMB[16][57] ) );
  FA1A S2_15_74 ( .A(\ab[15][74] ), .B(\CARRYB[14][74] ), .CI(\SUMB[14][75] ), 
        .CO(\CARRYB[15][74] ), .S(\SUMB[15][74] ) );
  FA1A S2_15_73 ( .A(\ab[15][73] ), .B(\CARRYB[14][73] ), .CI(\SUMB[14][74] ), 
        .CO(\CARRYB[15][73] ), .S(\SUMB[15][73] ) );
  FA1A S2_15_72 ( .A(\ab[15][72] ), .B(\CARRYB[14][72] ), .CI(\SUMB[14][73] ), 
        .CO(\CARRYB[15][72] ), .S(\SUMB[15][72] ) );
  FA1A S2_15_71 ( .A(\ab[15][71] ), .B(\CARRYB[14][71] ), .CI(\SUMB[14][72] ), 
        .CO(\CARRYB[15][71] ), .S(\SUMB[15][71] ) );
  FA1A S2_15_70 ( .A(\ab[15][70] ), .B(\CARRYB[14][70] ), .CI(\SUMB[14][71] ), 
        .CO(\CARRYB[15][70] ), .S(\SUMB[15][70] ) );
  FA1A S2_15_69 ( .A(\ab[15][69] ), .B(\CARRYB[14][69] ), .CI(\SUMB[14][70] ), 
        .CO(\CARRYB[15][69] ), .S(\SUMB[15][69] ) );
  FA1A S2_15_75 ( .A(\ab[15][75] ), .B(\CARRYB[14][75] ), .CI(\SUMB[14][76] ), 
        .CO(\CARRYB[15][75] ), .S(\SUMB[15][75] ) );
  FA1A S2_15_76 ( .A(\ab[15][76] ), .B(\CARRYB[14][76] ), .CI(\SUMB[14][77] ), 
        .CO(\CARRYB[15][76] ), .S(\SUMB[15][76] ) );
  FA1A S2_15_57 ( .A(\ab[15][57] ), .B(\CARRYB[14][57] ), .CI(\SUMB[14][58] ), 
        .CO(\CARRYB[15][57] ), .S(\SUMB[15][57] ) );
  FA1A S4_79 ( .A(\ab[29][79] ), .B(\CARRYB[28][79] ), .CI(\SUMB[28][80] ), 
        .CO(\CARRYB[29][79] ), .S(\SUMB[29][79] ) );
  FA1A S4_72 ( .A(\ab[29][72] ), .B(\CARRYB[28][72] ), .CI(\SUMB[28][73] ), 
        .CO(\CARRYB[29][72] ), .S(\SUMB[29][72] ) );
  FA1A S4_76 ( .A(\ab[29][76] ), .B(\CARRYB[28][76] ), .CI(\SUMB[28][77] ), 
        .CO(\CARRYB[29][76] ), .S(\SUMB[29][76] ) );
  FA1A S4_74 ( .A(\ab[29][74] ), .B(\CARRYB[28][74] ), .CI(\SUMB[28][75] ), 
        .CO(\CARRYB[29][74] ), .S(\SUMB[29][74] ) );
  FA1A S4_70 ( .A(\ab[29][70] ), .B(\CARRYB[28][70] ), .CI(\SUMB[28][71] ), 
        .CO(\CARRYB[29][70] ), .S(\SUMB[29][70] ) );
  FA1A S2_28_56 ( .A(\ab[28][56] ), .B(\CARRYB[27][56] ), .CI(\SUMB[27][57] ), 
        .CO(\CARRYB[28][56] ), .S(\SUMB[28][56] ) );
  FA1A S4_54 ( .A(\ab[29][54] ), .B(\CARRYB[28][54] ), .CI(\SUMB[28][55] ), 
        .CO(\CARRYB[29][54] ), .S(\SUMB[29][54] ) );
  FA1A S4_53 ( .A(\ab[29][53] ), .B(\CARRYB[28][53] ), .CI(\SUMB[28][54] ), 
        .CO(\CARRYB[29][53] ), .S(\SUMB[29][53] ) );
  FA1A S4_64 ( .A(\ab[29][64] ), .B(\CARRYB[28][64] ), .CI(\SUMB[28][65] ), 
        .CO(\CARRYB[29][64] ), .S(\SUMB[29][64] ) );
  FA1A S4_65 ( .A(\ab[29][65] ), .B(\CARRYB[28][65] ), .CI(\SUMB[28][66] ), 
        .CO(\CARRYB[29][65] ), .S(\SUMB[29][65] ) );
  FA1A S4_66 ( .A(\ab[29][66] ), .B(\CARRYB[28][66] ), .CI(\SUMB[28][67] ), 
        .CO(\CARRYB[29][66] ), .S(\SUMB[29][66] ) );
  FA1A S4_67 ( .A(\ab[29][67] ), .B(\CARRYB[28][67] ), .CI(\SUMB[28][68] ), 
        .CO(\CARRYB[29][67] ), .S(\SUMB[29][67] ) );
  FA1A S4_58 ( .A(\ab[29][58] ), .B(\CARRYB[28][58] ), .CI(\SUMB[28][59] ), 
        .CO(\CARRYB[29][58] ), .S(\SUMB[29][58] ) );
  FA1A S2_28_55 ( .A(\ab[28][55] ), .B(\CARRYB[27][55] ), .CI(\SUMB[27][56] ), 
        .CO(\CARRYB[28][55] ), .S(\SUMB[28][55] ) );
  FA1A S2_28_54 ( .A(\ab[28][54] ), .B(\CARRYB[27][54] ), .CI(\SUMB[27][55] ), 
        .CO(\CARRYB[28][54] ), .S(\SUMB[28][54] ) );
  FA1A S2_28_53 ( .A(\ab[28][53] ), .B(\CARRYB[27][53] ), .CI(\SUMB[27][54] ), 
        .CO(\CARRYB[28][53] ), .S(\SUMB[28][53] ) );
  FA1A S2_28_59 ( .A(\ab[28][59] ), .B(\CARRYB[27][59] ), .CI(\SUMB[27][60] ), 
        .CO(\CARRYB[28][59] ), .S(\SUMB[28][59] ) );
  FA1A S2_28_64 ( .A(\ab[28][64] ), .B(\CARRYB[27][64] ), .CI(\SUMB[27][65] ), 
        .CO(\CARRYB[28][64] ), .S(\SUMB[28][64] ) );
  FA1A S2_28_65 ( .A(\ab[28][65] ), .B(\CARRYB[27][65] ), .CI(\SUMB[27][66] ), 
        .CO(\CARRYB[28][65] ), .S(\SUMB[28][65] ) );
  FA1A S2_28_66 ( .A(\ab[28][66] ), .B(\CARRYB[27][66] ), .CI(\SUMB[27][67] ), 
        .CO(\CARRYB[28][66] ), .S(\SUMB[28][66] ) );
  FA1A S2_28_67 ( .A(\ab[28][67] ), .B(\CARRYB[27][67] ), .CI(\SUMB[27][68] ), 
        .CO(\CARRYB[28][67] ), .S(\SUMB[28][67] ) );
  FA1A S2_28_68 ( .A(\ab[28][68] ), .B(\CARRYB[27][68] ), .CI(\SUMB[27][69] ), 
        .CO(\CARRYB[28][68] ), .S(\SUMB[28][68] ) );
  FA1A S2_28_58 ( .A(\ab[28][58] ), .B(\CARRYB[27][58] ), .CI(\SUMB[27][59] ), 
        .CO(\CARRYB[28][58] ), .S(\SUMB[28][58] ) );
  FA1A S2_27_56 ( .A(\ab[27][56] ), .B(\CARRYB[26][56] ), .CI(\SUMB[26][57] ), 
        .CO(\CARRYB[27][56] ), .S(\SUMB[27][56] ) );
  FA1A S2_27_55 ( .A(\ab[27][55] ), .B(\CARRYB[26][55] ), .CI(\SUMB[26][56] ), 
        .CO(\CARRYB[27][55] ), .S(\SUMB[27][55] ) );
  FA1A S2_27_54 ( .A(\ab[27][54] ), .B(\CARRYB[26][54] ), .CI(\SUMB[26][55] ), 
        .CO(\CARRYB[27][54] ), .S(\SUMB[27][54] ) );
  FA1A S2_27_59 ( .A(\ab[27][59] ), .B(\CARRYB[26][59] ), .CI(\SUMB[26][60] ), 
        .CO(\CARRYB[27][59] ), .S(\SUMB[27][59] ) );
  FA1A S2_27_65 ( .A(\ab[27][65] ), .B(\CARRYB[26][65] ), .CI(\SUMB[26][66] ), 
        .CO(\CARRYB[27][65] ), .S(\SUMB[27][65] ) );
  FA1A S2_27_66 ( .A(\ab[27][66] ), .B(\CARRYB[26][66] ), .CI(\SUMB[26][67] ), 
        .CO(\CARRYB[27][66] ), .S(\SUMB[27][66] ) );
  FA1A S2_27_67 ( .A(\ab[27][67] ), .B(\CARRYB[26][67] ), .CI(\SUMB[26][68] ), 
        .CO(\CARRYB[27][67] ), .S(\SUMB[27][67] ) );
  FA1A S2_27_68 ( .A(\ab[27][68] ), .B(\CARRYB[26][68] ), .CI(\SUMB[26][69] ), 
        .CO(\CARRYB[27][68] ), .S(\SUMB[27][68] ) );
  FA1A S2_27_58 ( .A(\ab[27][58] ), .B(\CARRYB[26][58] ), .CI(\SUMB[26][59] ), 
        .CO(\CARRYB[27][58] ), .S(\SUMB[27][58] ) );
  FA1A S4_60 ( .A(\ab[29][60] ), .B(\CARRYB[28][60] ), .CI(\SUMB[28][61] ), 
        .CO(\CARRYB[29][60] ), .S(\SUMB[29][60] ) );
  FA1A S2_27_53 ( .A(\ab[27][53] ), .B(\CARRYB[26][53] ), .CI(\SUMB[26][54] ), 
        .CO(\CARRYB[27][53] ), .S(\SUMB[27][53] ) );
  FA1A S2_26_56 ( .A(\ab[26][56] ), .B(\CARRYB[25][56] ), .CI(\SUMB[25][57] ), 
        .CO(\CARRYB[26][56] ), .S(\SUMB[26][56] ) );
  FA1A S2_26_55 ( .A(\ab[26][55] ), .B(\CARRYB[25][55] ), .CI(\SUMB[25][56] ), 
        .CO(\CARRYB[26][55] ), .S(\SUMB[26][55] ) );
  FA1A S2_26_59 ( .A(\ab[26][59] ), .B(\CARRYB[25][59] ), .CI(\SUMB[25][60] ), 
        .CO(\CARRYB[26][59] ), .S(\SUMB[26][59] ) );
  FA1A S2_26_66 ( .A(\ab[26][66] ), .B(\CARRYB[25][66] ), .CI(\SUMB[25][67] ), 
        .CO(\CARRYB[26][66] ), .S(\SUMB[26][66] ) );
  FA1A S2_26_67 ( .A(\ab[26][67] ), .B(\CARRYB[25][67] ), .CI(\SUMB[25][68] ), 
        .CO(\CARRYB[26][67] ), .S(\SUMB[26][67] ) );
  FA1A S2_26_68 ( .A(\ab[26][68] ), .B(\CARRYB[25][68] ), .CI(\SUMB[25][69] ), 
        .CO(\CARRYB[26][68] ), .S(\SUMB[26][68] ) );
  FA1A S2_26_58 ( .A(\ab[26][58] ), .B(\CARRYB[25][58] ), .CI(\SUMB[25][59] ), 
        .CO(\CARRYB[26][58] ), .S(\SUMB[26][58] ) );
  FA1A S2_28_60 ( .A(\ab[28][60] ), .B(\CARRYB[27][60] ), .CI(\SUMB[27][61] ), 
        .CO(\CARRYB[28][60] ), .S(\SUMB[28][60] ) );
  FA1A S2_26_54 ( .A(\ab[26][54] ), .B(\CARRYB[25][54] ), .CI(\SUMB[25][55] ), 
        .CO(\CARRYB[26][54] ), .S(\SUMB[26][54] ) );
  FA1A S2_25_56 ( .A(\ab[25][56] ), .B(\CARRYB[24][56] ), .CI(\SUMB[24][57] ), 
        .CO(\CARRYB[25][56] ), .S(\SUMB[25][56] ) );
  FA1A S2_25_59 ( .A(\ab[25][59] ), .B(\CARRYB[24][59] ), .CI(\SUMB[24][60] ), 
        .CO(\CARRYB[25][59] ), .S(\SUMB[25][59] ) );
  FA1A S2_25_67 ( .A(\ab[25][67] ), .B(\CARRYB[24][67] ), .CI(\SUMB[24][68] ), 
        .CO(\CARRYB[25][67] ), .S(\SUMB[25][67] ) );
  FA1A S2_25_68 ( .A(\ab[25][68] ), .B(\CARRYB[24][68] ), .CI(\SUMB[24][69] ), 
        .CO(\CARRYB[25][68] ), .S(\SUMB[25][68] ) );
  FA1A S2_25_58 ( .A(\ab[25][58] ), .B(\CARRYB[24][58] ), .CI(\SUMB[24][59] ), 
        .CO(\CARRYB[25][58] ), .S(\SUMB[25][58] ) );
  FA1A S2_27_60 ( .A(\ab[27][60] ), .B(\CARRYB[26][60] ), .CI(\SUMB[26][61] ), 
        .CO(\CARRYB[27][60] ), .S(\SUMB[27][60] ) );
  FA1A S2_27_64 ( .A(\ab[27][64] ), .B(\CARRYB[26][64] ), .CI(\SUMB[26][65] ), 
        .CO(\CARRYB[27][64] ), .S(\SUMB[27][64] ) );
  FA1A S2_25_55 ( .A(\ab[25][55] ), .B(\CARRYB[24][55] ), .CI(\SUMB[24][56] ), 
        .CO(\CARRYB[25][55] ), .S(\SUMB[25][55] ) );
  FA1A S2_24_59 ( .A(\ab[24][59] ), .B(\CARRYB[23][59] ), .CI(\SUMB[23][60] ), 
        .CO(\CARRYB[24][59] ), .S(\SUMB[24][59] ) );
  FA1A S2_24_68 ( .A(\ab[24][68] ), .B(\CARRYB[23][68] ), .CI(\SUMB[23][69] ), 
        .CO(\CARRYB[24][68] ), .S(\SUMB[24][68] ) );
  FA1A S2_24_58 ( .A(\ab[24][58] ), .B(\CARRYB[23][58] ), .CI(\SUMB[23][59] ), 
        .CO(\CARRYB[24][58] ), .S(\SUMB[24][58] ) );
  FA1A S2_26_60 ( .A(\ab[26][60] ), .B(\CARRYB[25][60] ), .CI(\SUMB[25][61] ), 
        .CO(\CARRYB[26][60] ), .S(\SUMB[26][60] ) );
  FA1A S2_26_64 ( .A(\ab[26][64] ), .B(\CARRYB[25][64] ), .CI(\SUMB[25][65] ), 
        .CO(\CARRYB[26][64] ), .S(\SUMB[26][64] ) );
  FA1A S2_26_65 ( .A(\ab[26][65] ), .B(\CARRYB[25][65] ), .CI(\SUMB[25][66] ), 
        .CO(\CARRYB[26][65] ), .S(\SUMB[26][65] ) );
  FA1A S2_24_56 ( .A(\ab[24][56] ), .B(\CARRYB[23][56] ), .CI(\SUMB[23][57] ), 
        .CO(\CARRYB[24][56] ), .S(\SUMB[24][56] ) );
  FA1A S2_26_53 ( .A(\ab[26][53] ), .B(\CARRYB[25][53] ), .CI(\SUMB[25][54] ), 
        .CO(\CARRYB[26][53] ), .S(\SUMB[26][53] ) );
  FA1A S2_23_59 ( .A(\ab[23][59] ), .B(\CARRYB[22][59] ), .CI(\SUMB[22][60] ), 
        .CO(\CARRYB[23][59] ), .S(\SUMB[23][59] ) );
  FA1A S2_23_58 ( .A(\ab[23][58] ), .B(\CARRYB[22][58] ), .CI(\SUMB[22][59] ), 
        .CO(\CARRYB[23][58] ), .S(\SUMB[23][58] ) );
  FA1A S2_25_64 ( .A(\ab[25][64] ), .B(\CARRYB[24][64] ), .CI(\SUMB[24][65] ), 
        .CO(\CARRYB[25][64] ), .S(\SUMB[25][64] ) );
  FA1A S2_25_60 ( .A(\ab[25][60] ), .B(\CARRYB[24][60] ), .CI(\SUMB[24][61] ), 
        .CO(\CARRYB[25][60] ), .S(\SUMB[25][60] ) );
  FA1A S2_25_65 ( .A(\ab[25][65] ), .B(\CARRYB[24][65] ), .CI(\SUMB[24][66] ), 
        .CO(\CARRYB[25][65] ), .S(\SUMB[25][65] ) );
  FA1A S2_25_66 ( .A(\ab[25][66] ), .B(\CARRYB[24][66] ), .CI(\SUMB[24][67] ), 
        .CO(\CARRYB[25][66] ), .S(\SUMB[25][66] ) );
  FA1A S2_25_53 ( .A(\ab[25][53] ), .B(\CARRYB[24][53] ), .CI(\SUMB[24][54] ), 
        .CO(\CARRYB[25][53] ), .S(\SUMB[25][53] ) );
  FA1A S2_25_54 ( .A(\ab[25][54] ), .B(\CARRYB[24][54] ), .CI(\SUMB[24][55] ), 
        .CO(\CARRYB[25][54] ), .S(\SUMB[25][54] ) );
  FA1A S2_22_59 ( .A(\ab[22][59] ), .B(\CARRYB[21][59] ), .CI(\SUMB[21][60] ), 
        .CO(\CARRYB[22][59] ), .S(\SUMB[22][59] ) );
  FA1A S2_22_58 ( .A(\ab[22][58] ), .B(\CARRYB[21][58] ), .CI(\SUMB[21][59] ), 
        .CO(\CARRYB[22][58] ), .S(\SUMB[22][58] ) );
  FA1A S2_24_65 ( .A(\ab[24][65] ), .B(\CARRYB[23][65] ), .CI(\SUMB[23][66] ), 
        .CO(\CARRYB[24][65] ), .S(\SUMB[24][65] ) );
  FA1A S2_24_64 ( .A(\ab[24][64] ), .B(\CARRYB[23][64] ), .CI(\SUMB[23][65] ), 
        .CO(\CARRYB[24][64] ), .S(\SUMB[24][64] ) );
  FA1A S2_24_60 ( .A(\ab[24][60] ), .B(\CARRYB[23][60] ), .CI(\SUMB[23][61] ), 
        .CO(\CARRYB[24][60] ), .S(\SUMB[24][60] ) );
  FA1A S2_24_66 ( .A(\ab[24][66] ), .B(\CARRYB[23][66] ), .CI(\SUMB[23][67] ), 
        .CO(\CARRYB[24][66] ), .S(\SUMB[24][66] ) );
  FA1A S2_24_67 ( .A(\ab[24][67] ), .B(\CARRYB[23][67] ), .CI(\SUMB[23][68] ), 
        .CO(\CARRYB[24][67] ), .S(\SUMB[24][67] ) );
  FA1A S2_24_53 ( .A(\ab[24][53] ), .B(\CARRYB[23][53] ), .CI(\SUMB[23][54] ), 
        .CO(\CARRYB[24][53] ), .S(\SUMB[24][53] ) );
  FA1A S2_24_54 ( .A(\ab[24][54] ), .B(\CARRYB[23][54] ), .CI(\SUMB[23][55] ), 
        .CO(\CARRYB[24][54] ), .S(\SUMB[24][54] ) );
  FA1A S2_24_55 ( .A(\ab[24][55] ), .B(\CARRYB[23][55] ), .CI(\SUMB[23][56] ), 
        .CO(\CARRYB[24][55] ), .S(\SUMB[24][55] ) );
  FA1A S2_21_59 ( .A(\ab[21][59] ), .B(\CARRYB[20][59] ), .CI(\SUMB[20][60] ), 
        .CO(\CARRYB[21][59] ), .S(\SUMB[21][59] ) );
  FA1A S2_23_66 ( .A(\ab[23][66] ), .B(\CARRYB[22][66] ), .CI(\SUMB[22][67] ), 
        .CO(\CARRYB[23][66] ), .S(\SUMB[23][66] ) );
  FA1A S2_23_65 ( .A(\ab[23][65] ), .B(\CARRYB[22][65] ), .CI(\SUMB[22][66] ), 
        .CO(\CARRYB[23][65] ), .S(\SUMB[23][65] ) );
  FA1A S2_23_64 ( .A(\ab[23][64] ), .B(\CARRYB[22][64] ), .CI(\SUMB[22][65] ), 
        .CO(\CARRYB[23][64] ), .S(\SUMB[23][64] ) );
  FA1A S2_23_60 ( .A(\ab[23][60] ), .B(\CARRYB[22][60] ), .CI(\SUMB[22][61] ), 
        .CO(\CARRYB[23][60] ), .S(\SUMB[23][60] ) );
  FA1A S2_23_67 ( .A(\ab[23][67] ), .B(\CARRYB[22][67] ), .CI(\SUMB[22][68] ), 
        .CO(\CARRYB[23][67] ), .S(\SUMB[23][67] ) );
  FA1A S2_23_68 ( .A(\ab[23][68] ), .B(\CARRYB[22][68] ), .CI(\SUMB[22][69] ), 
        .CO(\CARRYB[23][68] ), .S(\SUMB[23][68] ) );
  FA1A S2_23_54 ( .A(\ab[23][54] ), .B(\CARRYB[22][54] ), .CI(\SUMB[22][55] ), 
        .CO(\CARRYB[23][54] ), .S(\SUMB[23][54] ) );
  FA1A S2_23_53 ( .A(\ab[23][53] ), .B(\CARRYB[22][53] ), .CI(\SUMB[22][54] ), 
        .CO(\CARRYB[23][53] ), .S(\SUMB[23][53] ) );
  FA1A S2_23_55 ( .A(\ab[23][55] ), .B(\CARRYB[22][55] ), .CI(\SUMB[22][56] ), 
        .CO(\CARRYB[23][55] ), .S(\SUMB[23][55] ) );
  FA1A S2_23_56 ( .A(\ab[23][56] ), .B(\CARRYB[22][56] ), .CI(\SUMB[22][57] ), 
        .CO(\CARRYB[23][56] ), .S(\SUMB[23][56] ) );
  FA1A S2_22_67 ( .A(\ab[22][67] ), .B(\CARRYB[21][67] ), .CI(\SUMB[21][68] ), 
        .CO(\CARRYB[22][67] ), .S(\SUMB[22][67] ) );
  FA1A S2_22_66 ( .A(\ab[22][66] ), .B(\CARRYB[21][66] ), .CI(\SUMB[21][67] ), 
        .CO(\CARRYB[22][66] ), .S(\SUMB[22][66] ) );
  FA1A S2_22_65 ( .A(\ab[22][65] ), .B(\CARRYB[21][65] ), .CI(\SUMB[21][66] ), 
        .CO(\CARRYB[22][65] ), .S(\SUMB[22][65] ) );
  FA1A S2_22_64 ( .A(\ab[22][64] ), .B(\CARRYB[21][64] ), .CI(\SUMB[21][65] ), 
        .CO(\CARRYB[22][64] ), .S(\SUMB[22][64] ) );
  FA1A S2_22_60 ( .A(\ab[22][60] ), .B(\CARRYB[21][60] ), .CI(\SUMB[21][61] ), 
        .CO(\CARRYB[22][60] ), .S(\SUMB[22][60] ) );
  FA1A S2_22_68 ( .A(\ab[22][68] ), .B(\CARRYB[21][68] ), .CI(\SUMB[21][69] ), 
        .CO(\CARRYB[22][68] ), .S(\SUMB[22][68] ) );
  FA1A S2_22_55 ( .A(\ab[22][55] ), .B(\CARRYB[21][55] ), .CI(\SUMB[21][56] ), 
        .CO(\CARRYB[22][55] ), .S(\SUMB[22][55] ) );
  FA1A S2_22_54 ( .A(\ab[22][54] ), .B(\CARRYB[21][54] ), .CI(\SUMB[21][55] ), 
        .CO(\CARRYB[22][54] ), .S(\SUMB[22][54] ) );
  FA1A S2_22_53 ( .A(\ab[22][53] ), .B(\CARRYB[21][53] ), .CI(\SUMB[21][54] ), 
        .CO(\CARRYB[22][53] ), .S(\SUMB[22][53] ) );
  FA1A S2_22_56 ( .A(\ab[22][56] ), .B(\CARRYB[21][56] ), .CI(\SUMB[21][57] ), 
        .CO(\CARRYB[22][56] ), .S(\SUMB[22][56] ) );
  FA1A S2_21_68 ( .A(\ab[21][68] ), .B(\CARRYB[20][68] ), .CI(\SUMB[20][69] ), 
        .CO(\CARRYB[21][68] ), .S(\SUMB[21][68] ) );
  FA1A S2_21_67 ( .A(\ab[21][67] ), .B(\CARRYB[20][67] ), .CI(\SUMB[20][68] ), 
        .CO(\CARRYB[21][67] ), .S(\SUMB[21][67] ) );
  FA1A S2_21_66 ( .A(\ab[21][66] ), .B(\CARRYB[20][66] ), .CI(\SUMB[20][67] ), 
        .CO(\CARRYB[21][66] ), .S(\SUMB[21][66] ) );
  FA1A S2_21_65 ( .A(\ab[21][65] ), .B(\CARRYB[20][65] ), .CI(\SUMB[20][66] ), 
        .CO(\CARRYB[21][65] ), .S(\SUMB[21][65] ) );
  FA1A S2_21_64 ( .A(\ab[21][64] ), .B(\CARRYB[20][64] ), .CI(\SUMB[20][65] ), 
        .CO(\CARRYB[21][64] ), .S(\SUMB[21][64] ) );
  FA1A S2_21_60 ( .A(\ab[21][60] ), .B(\CARRYB[20][60] ), .CI(\SUMB[20][61] ), 
        .CO(\CARRYB[21][60] ), .S(\SUMB[21][60] ) );
  FA1A S2_21_56 ( .A(\ab[21][56] ), .B(\CARRYB[20][56] ), .CI(\SUMB[20][57] ), 
        .CO(\CARRYB[21][56] ), .S(\SUMB[21][56] ) );
  FA1A S2_21_55 ( .A(\ab[21][55] ), .B(\CARRYB[20][55] ), .CI(\SUMB[20][56] ), 
        .CO(\CARRYB[21][55] ), .S(\SUMB[21][55] ) );
  FA1A S2_21_54 ( .A(\ab[21][54] ), .B(\CARRYB[20][54] ), .CI(\SUMB[20][55] ), 
        .CO(\CARRYB[21][54] ), .S(\SUMB[21][54] ) );
  FA1A S2_21_53 ( .A(\ab[21][53] ), .B(\CARRYB[20][53] ), .CI(\SUMB[20][54] ), 
        .CO(\CARRYB[21][53] ), .S(\SUMB[21][53] ) );
  FA1A S2_21_58 ( .A(\ab[21][58] ), .B(\CARRYB[20][58] ), .CI(\SUMB[20][59] ), 
        .CO(\CARRYB[21][58] ), .S(\SUMB[21][58] ) );
  FA1A S2_20_68 ( .A(\ab[20][68] ), .B(\CARRYB[19][68] ), .CI(\SUMB[19][69] ), 
        .CO(\CARRYB[20][68] ), .S(\SUMB[20][68] ) );
  FA1A S2_20_67 ( .A(\ab[20][67] ), .B(\CARRYB[19][67] ), .CI(\SUMB[19][68] ), 
        .CO(\CARRYB[20][67] ), .S(\SUMB[20][67] ) );
  FA1A S2_20_66 ( .A(\ab[20][66] ), .B(\CARRYB[19][66] ), .CI(\SUMB[19][67] ), 
        .CO(\CARRYB[20][66] ), .S(\SUMB[20][66] ) );
  FA1A S2_20_65 ( .A(\ab[20][65] ), .B(\CARRYB[19][65] ), .CI(\SUMB[19][66] ), 
        .CO(\CARRYB[20][65] ), .S(\SUMB[20][65] ) );
  FA1A S2_20_64 ( .A(\ab[20][64] ), .B(\CARRYB[19][64] ), .CI(\SUMB[19][65] ), 
        .CO(\CARRYB[20][64] ), .S(\SUMB[20][64] ) );
  FA1A S2_20_60 ( .A(\ab[20][60] ), .B(\CARRYB[19][60] ), .CI(\SUMB[19][61] ), 
        .CO(\CARRYB[20][60] ), .S(\SUMB[20][60] ) );
  FA1A S2_20_56 ( .A(\ab[20][56] ), .B(\CARRYB[19][56] ), .CI(\SUMB[19][57] ), 
        .CO(\CARRYB[20][56] ), .S(\SUMB[20][56] ) );
  FA1A S2_20_55 ( .A(\ab[20][55] ), .B(\CARRYB[19][55] ), .CI(\SUMB[19][56] ), 
        .CO(\CARRYB[20][55] ), .S(\SUMB[20][55] ) );
  FA1A S2_20_54 ( .A(\ab[20][54] ), .B(\CARRYB[19][54] ), .CI(\SUMB[19][55] ), 
        .CO(\CARRYB[20][54] ), .S(\SUMB[20][54] ) );
  FA1A S2_20_53 ( .A(\ab[20][53] ), .B(\CARRYB[19][53] ), .CI(\SUMB[19][54] ), 
        .CO(\CARRYB[20][53] ), .S(\SUMB[20][53] ) );
  FA1A S2_20_58 ( .A(\ab[20][58] ), .B(\CARRYB[19][58] ), .CI(\SUMB[19][59] ), 
        .CO(\CARRYB[20][58] ), .S(\SUMB[20][58] ) );
  FA1A S2_20_59 ( .A(\ab[20][59] ), .B(\CARRYB[19][59] ), .CI(\SUMB[19][60] ), 
        .CO(\CARRYB[20][59] ), .S(\SUMB[20][59] ) );
  FA1A S2_19_68 ( .A(\ab[19][68] ), .B(\CARRYB[18][68] ), .CI(\SUMB[18][69] ), 
        .CO(\CARRYB[19][68] ), .S(\SUMB[19][68] ) );
  FA1A S2_19_67 ( .A(\ab[19][67] ), .B(\CARRYB[18][67] ), .CI(\SUMB[18][68] ), 
        .CO(\CARRYB[19][67] ), .S(\SUMB[19][67] ) );
  FA1A S2_19_66 ( .A(\ab[19][66] ), .B(\CARRYB[18][66] ), .CI(\SUMB[18][67] ), 
        .CO(\CARRYB[19][66] ), .S(\SUMB[19][66] ) );
  FA1A S2_19_65 ( .A(\ab[19][65] ), .B(\CARRYB[18][65] ), .CI(\SUMB[18][66] ), 
        .CO(\CARRYB[19][65] ), .S(\SUMB[19][65] ) );
  FA1A S2_19_64 ( .A(\ab[19][64] ), .B(\CARRYB[18][64] ), .CI(\SUMB[18][65] ), 
        .CO(\CARRYB[19][64] ), .S(\SUMB[19][64] ) );
  FA1A S2_19_60 ( .A(\ab[19][60] ), .B(\CARRYB[18][60] ), .CI(\SUMB[18][61] ), 
        .CO(\CARRYB[19][60] ), .S(\SUMB[19][60] ) );
  FA1A S2_19_58 ( .A(\ab[19][58] ), .B(\CARRYB[18][58] ), .CI(\SUMB[18][59] ), 
        .CO(\CARRYB[19][58] ), .S(\SUMB[19][58] ) );
  FA1A S2_19_56 ( .A(\ab[19][56] ), .B(\CARRYB[18][56] ), .CI(\SUMB[18][57] ), 
        .CO(\CARRYB[19][56] ), .S(\SUMB[19][56] ) );
  FA1A S2_19_55 ( .A(\ab[19][55] ), .B(\CARRYB[18][55] ), .CI(\SUMB[18][56] ), 
        .CO(\CARRYB[19][55] ), .S(\SUMB[19][55] ) );
  FA1A S2_19_54 ( .A(\ab[19][54] ), .B(\CARRYB[18][54] ), .CI(\SUMB[18][55] ), 
        .CO(\CARRYB[19][54] ), .S(\SUMB[19][54] ) );
  FA1A S2_19_53 ( .A(\ab[19][53] ), .B(\CARRYB[18][53] ), .CI(\SUMB[18][54] ), 
        .CO(\CARRYB[19][53] ), .S(\SUMB[19][53] ) );
  FA1A S2_19_59 ( .A(\ab[19][59] ), .B(\CARRYB[18][59] ), .CI(\SUMB[18][60] ), 
        .CO(\CARRYB[19][59] ), .S(\SUMB[19][59] ) );
  FA1A S2_18_68 ( .A(\ab[18][68] ), .B(\CARRYB[17][68] ), .CI(\SUMB[17][69] ), 
        .CO(\CARRYB[18][68] ), .S(\SUMB[18][68] ) );
  FA1A S2_18_67 ( .A(\ab[18][67] ), .B(\CARRYB[17][67] ), .CI(\SUMB[17][68] ), 
        .CO(\CARRYB[18][67] ), .S(\SUMB[18][67] ) );
  FA1A S2_18_66 ( .A(\ab[18][66] ), .B(\CARRYB[17][66] ), .CI(\SUMB[17][67] ), 
        .CO(\CARRYB[18][66] ), .S(\SUMB[18][66] ) );
  FA1A S2_18_65 ( .A(\ab[18][65] ), .B(\CARRYB[17][65] ), .CI(\SUMB[17][66] ), 
        .CO(\CARRYB[18][65] ), .S(\SUMB[18][65] ) );
  FA1A S2_18_64 ( .A(\ab[18][64] ), .B(\CARRYB[17][64] ), .CI(\SUMB[17][65] ), 
        .CO(\CARRYB[18][64] ), .S(\SUMB[18][64] ) );
  FA1A S2_18_60 ( .A(\ab[18][60] ), .B(\CARRYB[17][60] ), .CI(\SUMB[17][61] ), 
        .CO(\CARRYB[18][60] ), .S(\SUMB[18][60] ) );
  FA1A S2_18_53 ( .A(\ab[18][53] ), .B(\CARRYB[17][53] ), .CI(\SUMB[17][54] ), 
        .CO(\CARRYB[18][53] ), .S(\SUMB[18][53] ) );
  FA1A S2_18_59 ( .A(\ab[18][59] ), .B(\CARRYB[17][59] ), .CI(\SUMB[17][60] ), 
        .CO(\CARRYB[18][59] ), .S(\SUMB[18][59] ) );
  FA1A S2_18_58 ( .A(\ab[18][58] ), .B(\CARRYB[17][58] ), .CI(\SUMB[17][59] ), 
        .CO(\CARRYB[18][58] ), .S(\SUMB[18][58] ) );
  FA1A S2_18_56 ( .A(\ab[18][56] ), .B(\CARRYB[17][56] ), .CI(\SUMB[17][57] ), 
        .CO(\CARRYB[18][56] ), .S(\SUMB[18][56] ) );
  FA1A S2_18_55 ( .A(\ab[18][55] ), .B(\CARRYB[17][55] ), .CI(\SUMB[17][56] ), 
        .CO(\CARRYB[18][55] ), .S(\SUMB[18][55] ) );
  FA1A S2_18_54 ( .A(\ab[18][54] ), .B(\CARRYB[17][54] ), .CI(\SUMB[17][55] ), 
        .CO(\CARRYB[18][54] ), .S(\SUMB[18][54] ) );
  FA1A S2_17_68 ( .A(\ab[17][68] ), .B(\CARRYB[16][68] ), .CI(\SUMB[16][69] ), 
        .CO(\CARRYB[17][68] ), .S(\SUMB[17][68] ) );
  FA1A S2_17_67 ( .A(\ab[17][67] ), .B(\CARRYB[16][67] ), .CI(\SUMB[16][68] ), 
        .CO(\CARRYB[17][67] ), .S(\SUMB[17][67] ) );
  FA1A S2_17_66 ( .A(\ab[17][66] ), .B(\CARRYB[16][66] ), .CI(\SUMB[16][67] ), 
        .CO(\CARRYB[17][66] ), .S(\SUMB[17][66] ) );
  FA1A S2_17_65 ( .A(\ab[17][65] ), .B(\CARRYB[16][65] ), .CI(\SUMB[16][66] ), 
        .CO(\CARRYB[17][65] ), .S(\SUMB[17][65] ) );
  FA1A S2_17_64 ( .A(\ab[17][64] ), .B(\CARRYB[16][64] ), .CI(\SUMB[16][65] ), 
        .CO(\CARRYB[17][64] ), .S(\SUMB[17][64] ) );
  FA1A S2_17_60 ( .A(\ab[17][60] ), .B(\CARRYB[16][60] ), .CI(\SUMB[16][61] ), 
        .CO(\CARRYB[17][60] ), .S(\SUMB[17][60] ) );
  FA1A S2_17_54 ( .A(\ab[17][54] ), .B(\CARRYB[16][54] ), .CI(\SUMB[16][55] ), 
        .CO(\CARRYB[17][54] ), .S(\SUMB[17][54] ) );
  FA1A S2_17_53 ( .A(\ab[17][53] ), .B(\CARRYB[16][53] ), .CI(\SUMB[16][54] ), 
        .CO(\CARRYB[17][53] ), .S(\SUMB[17][53] ) );
  FA1A S2_17_59 ( .A(\ab[17][59] ), .B(\CARRYB[16][59] ), .CI(\SUMB[16][60] ), 
        .CO(\CARRYB[17][59] ), .S(\SUMB[17][59] ) );
  FA1A S2_17_58 ( .A(\ab[17][58] ), .B(\CARRYB[16][58] ), .CI(\SUMB[16][59] ), 
        .CO(\CARRYB[17][58] ), .S(\SUMB[17][58] ) );
  FA1A S2_17_56 ( .A(\ab[17][56] ), .B(\CARRYB[16][56] ), .CI(\SUMB[16][57] ), 
        .CO(\CARRYB[17][56] ), .S(\SUMB[17][56] ) );
  FA1A S2_17_55 ( .A(\ab[17][55] ), .B(\CARRYB[16][55] ), .CI(\SUMB[16][56] ), 
        .CO(\CARRYB[17][55] ), .S(\SUMB[17][55] ) );
  FA1A S2_16_68 ( .A(\ab[16][68] ), .B(\CARRYB[15][68] ), .CI(\SUMB[15][69] ), 
        .CO(\CARRYB[16][68] ), .S(\SUMB[16][68] ) );
  FA1A S2_16_67 ( .A(\ab[16][67] ), .B(\CARRYB[15][67] ), .CI(\SUMB[15][68] ), 
        .CO(\CARRYB[16][67] ), .S(\SUMB[16][67] ) );
  FA1A S2_16_66 ( .A(\ab[16][66] ), .B(\CARRYB[15][66] ), .CI(\SUMB[15][67] ), 
        .CO(\CARRYB[16][66] ), .S(\SUMB[16][66] ) );
  FA1A S2_16_65 ( .A(\ab[16][65] ), .B(\CARRYB[15][65] ), .CI(\SUMB[15][66] ), 
        .CO(\CARRYB[16][65] ), .S(\SUMB[16][65] ) );
  FA1A S2_16_64 ( .A(\ab[16][64] ), .B(\CARRYB[15][64] ), .CI(\SUMB[15][65] ), 
        .CO(\CARRYB[16][64] ), .S(\SUMB[16][64] ) );
  FA1A S2_16_60 ( .A(\ab[16][60] ), .B(\CARRYB[15][60] ), .CI(\SUMB[15][61] ), 
        .CO(\CARRYB[16][60] ), .S(\SUMB[16][60] ) );
  FA1A S2_16_55 ( .A(\ab[16][55] ), .B(\CARRYB[15][55] ), .CI(\SUMB[15][56] ), 
        .CO(\CARRYB[16][55] ), .S(\SUMB[16][55] ) );
  FA1A S2_16_54 ( .A(\ab[16][54] ), .B(\CARRYB[15][54] ), .CI(\SUMB[15][55] ), 
        .CO(\CARRYB[16][54] ), .S(\SUMB[16][54] ) );
  FA1A S2_16_53 ( .A(\ab[16][53] ), .B(\CARRYB[15][53] ), .CI(\SUMB[15][54] ), 
        .CO(\CARRYB[16][53] ), .S(\SUMB[16][53] ) );
  FA1A S2_16_59 ( .A(\ab[16][59] ), .B(\CARRYB[15][59] ), .CI(\SUMB[15][60] ), 
        .CO(\CARRYB[16][59] ), .S(\SUMB[16][59] ) );
  FA1A S2_16_58 ( .A(\ab[16][58] ), .B(\CARRYB[15][58] ), .CI(\SUMB[15][59] ), 
        .CO(\CARRYB[16][58] ), .S(\SUMB[16][58] ) );
  FA1A S2_16_56 ( .A(\ab[16][56] ), .B(\CARRYB[15][56] ), .CI(\SUMB[15][57] ), 
        .CO(\CARRYB[16][56] ), .S(\SUMB[16][56] ) );
  FA1A S2_15_68 ( .A(\ab[15][68] ), .B(\CARRYB[14][68] ), .CI(\SUMB[14][69] ), 
        .CO(\CARRYB[15][68] ), .S(\SUMB[15][68] ) );
  FA1A S2_15_67 ( .A(\ab[15][67] ), .B(\CARRYB[14][67] ), .CI(\SUMB[14][68] ), 
        .CO(\CARRYB[15][67] ), .S(\SUMB[15][67] ) );
  FA1A S2_15_66 ( .A(\ab[15][66] ), .B(\CARRYB[14][66] ), .CI(\SUMB[14][67] ), 
        .CO(\CARRYB[15][66] ), .S(\SUMB[15][66] ) );
  FA1A S2_15_65 ( .A(\ab[15][65] ), .B(\CARRYB[14][65] ), .CI(\SUMB[14][66] ), 
        .CO(\CARRYB[15][65] ), .S(\SUMB[15][65] ) );
  FA1A S2_15_64 ( .A(\ab[15][64] ), .B(\CARRYB[14][64] ), .CI(\SUMB[14][65] ), 
        .CO(\CARRYB[15][64] ), .S(\SUMB[15][64] ) );
  FA1A S2_15_60 ( .A(\ab[15][60] ), .B(\CARRYB[14][60] ), .CI(\SUMB[14][61] ), 
        .CO(\CARRYB[15][60] ), .S(\SUMB[15][60] ) );
  FA1A S2_15_56 ( .A(\ab[15][56] ), .B(\CARRYB[14][56] ), .CI(\SUMB[14][57] ), 
        .CO(\CARRYB[15][56] ), .S(\SUMB[15][56] ) );
  FA1A S2_15_55 ( .A(\ab[15][55] ), .B(\CARRYB[14][55] ), .CI(\SUMB[14][56] ), 
        .CO(\CARRYB[15][55] ), .S(\SUMB[15][55] ) );
  FA1A S2_15_54 ( .A(\ab[15][54] ), .B(\CARRYB[14][54] ), .CI(\SUMB[14][55] ), 
        .CO(\CARRYB[15][54] ), .S(\SUMB[15][54] ) );
  FA1A S2_15_53 ( .A(\ab[15][53] ), .B(\CARRYB[14][53] ), .CI(\SUMB[14][54] ), 
        .CO(\CARRYB[15][53] ), .S(\SUMB[15][53] ) );
  FA1A S2_15_59 ( .A(\ab[15][59] ), .B(\CARRYB[14][59] ), .CI(\SUMB[14][60] ), 
        .CO(\CARRYB[15][59] ), .S(\SUMB[15][59] ) );
  FA1A S2_15_58 ( .A(\ab[15][58] ), .B(\CARRYB[14][58] ), .CI(\SUMB[14][59] ), 
        .CO(\CARRYB[15][58] ), .S(\SUMB[15][58] ) );
  FA1A S2_14_55 ( .A(\ab[14][55] ), .B(\CARRYB[13][55] ), .CI(\SUMB[13][56] ), 
        .CO(\CARRYB[14][55] ), .S(\SUMB[14][55] ) );
  FA1A S2_13_55 ( .A(\ab[13][55] ), .B(\CARRYB[12][55] ), .CI(\SUMB[12][56] ), 
        .CO(\CARRYB[13][55] ), .S(\SUMB[13][55] ) );
  FA1A S2_12_55 ( .A(\ab[12][55] ), .B(\CARRYB[11][55] ), .CI(\SUMB[11][56] ), 
        .CO(\CARRYB[12][55] ), .S(\SUMB[12][55] ) );
  FA1A S2_11_55 ( .A(\ab[11][55] ), .B(\CARRYB[10][55] ), .CI(\SUMB[10][56] ), 
        .CO(\CARRYB[11][55] ), .S(\SUMB[11][55] ) );
  FA1A S2_10_55 ( .A(\ab[10][55] ), .B(\CARRYB[9][55] ), .CI(\SUMB[9][56] ), 
        .CO(\CARRYB[10][55] ), .S(\SUMB[10][55] ) );
  FA1A S2_9_55 ( .A(\ab[9][55] ), .B(\CARRYB[8][55] ), .CI(\SUMB[8][56] ), 
        .CO(\CARRYB[9][55] ), .S(\SUMB[9][55] ) );
  FA1A S2_8_55 ( .A(\ab[8][55] ), .B(\CARRYB[7][55] ), .CI(\SUMB[7][56] ), 
        .CO(\CARRYB[8][55] ), .S(\SUMB[8][55] ) );
  FA1A S2_7_55 ( .A(\ab[7][55] ), .B(\CARRYB[6][55] ), .CI(\SUMB[6][56] ), 
        .CO(\CARRYB[7][55] ), .S(\SUMB[7][55] ) );
  FA1A S2_6_55 ( .A(\ab[6][55] ), .B(\CARRYB[5][55] ), .CI(\SUMB[5][56] ), 
        .CO(\CARRYB[6][55] ), .S(\SUMB[6][55] ) );
  FA1A S2_5_55 ( .A(\ab[5][55] ), .B(\CARRYB[4][55] ), .CI(\SUMB[4][56] ), 
        .CO(\CARRYB[5][55] ), .S(\SUMB[5][55] ) );
  FA1A S2_4_55 ( .A(\ab[4][55] ), .B(\CARRYB[3][55] ), .CI(\SUMB[3][56] ), 
        .CO(\CARRYB[4][55] ), .S(\SUMB[4][55] ) );
  FA1A S2_3_55 ( .A(\ab[3][55] ), .B(\CARRYB[2][55] ), .CI(\SUMB[2][56] ), 
        .CO(\CARRYB[3][55] ), .S(\SUMB[3][55] ) );
  FA1A S2_2_55 ( .A(\ab[2][55] ), .B(\CARRYB[1][55] ), .CI(\SUMB[1][56] ), 
        .CO(\CARRYB[2][55] ), .S(\SUMB[2][55] ) );
  FA1A S4_68 ( .A(\ab[29][68] ), .B(\CARRYB[28][68] ), .CI(\SUMB[28][69] ), 
        .CO(\CARRYB[29][68] ), .S(\SUMB[29][68] ) );
  FA1A S4_56 ( .A(\ab[29][56] ), .B(\CARRYB[28][56] ), .CI(\SUMB[28][57] ), 
        .CO(\CARRYB[29][56] ), .S(\SUMB[29][56] ) );
  FA1A S4_55 ( .A(\ab[29][55] ), .B(\CARRYB[28][55] ), .CI(\SUMB[28][56] ), 
        .CO(\CARRYB[29][55] ), .S(\SUMB[29][55] ) );
  FA1A S4_59 ( .A(\ab[29][59] ), .B(\CARRYB[28][59] ), .CI(\SUMB[28][60] ), 
        .CO(\CARRYB[29][59] ), .S(\SUMB[29][59] ) );
  FA1A S4_39 ( .A(\ab[29][39] ), .B(\CARRYB[28][39] ), .CI(\SUMB[28][40] ), 
        .CO(\CARRYB[29][39] ), .S(\SUMB[29][39] ) );
  FA1A S4_44 ( .A(\ab[29][44] ), .B(\CARRYB[28][44] ), .CI(\SUMB[28][45] ), 
        .CO(\CARRYB[29][44] ), .S(\SUMB[29][44] ) );
  FA1A S4_43 ( .A(\ab[29][43] ), .B(\CARRYB[28][43] ), .CI(\SUMB[28][44] ), 
        .CO(\CARRYB[29][43] ), .S(\SUMB[29][43] ) );
  FA1A S2_28_52 ( .A(\ab[28][52] ), .B(\CARRYB[27][52] ), .CI(\SUMB[27][53] ), 
        .CO(\CARRYB[28][52] ), .S(\SUMB[28][52] ) );
  FA1A S2_28_44 ( .A(\ab[28][44] ), .B(\CARRYB[27][44] ), .CI(\SUMB[27][45] ), 
        .CO(\CARRYB[28][44] ), .S(\SUMB[28][44] ) );
  FA1A S4_61 ( .A(\ab[29][61] ), .B(\CARRYB[28][61] ), .CI(\SUMB[28][62] ), 
        .CO(\CARRYB[29][61] ), .S(\SUMB[29][61] ) );
  FA1A S4_62 ( .A(\ab[29][62] ), .B(\CARRYB[28][62] ), .CI(\SUMB[28][63] ), 
        .CO(\CARRYB[29][62] ), .S(\SUMB[29][62] ) );
  FA1A S4_42 ( .A(\ab[29][42] ), .B(\CARRYB[28][42] ), .CI(\SUMB[28][43] ), 
        .CO(\CARRYB[29][42] ), .S(\SUMB[29][42] ) );
  FA1A S4_41 ( .A(\ab[29][41] ), .B(\CARRYB[28][41] ), .CI(\SUMB[28][42] ), 
        .CO(\CARRYB[29][41] ), .S(\SUMB[29][41] ) );
  FA1A S4_40 ( .A(\ab[29][40] ), .B(\CARRYB[28][40] ), .CI(\SUMB[28][41] ), 
        .CO(\CARRYB[29][40] ), .S(\SUMB[29][40] ) );
  FA1A S2_28_61 ( .A(\ab[28][61] ), .B(\CARRYB[27][61] ), .CI(\SUMB[27][62] ), 
        .CO(\CARRYB[28][61] ), .S(\SUMB[28][61] ) );
  FA1A S2_28_62 ( .A(\ab[28][62] ), .B(\CARRYB[27][62] ), .CI(\SUMB[27][63] ), 
        .CO(\CARRYB[28][62] ), .S(\SUMB[28][62] ) );
  FA1A S2_28_63 ( .A(\ab[28][63] ), .B(\CARRYB[27][63] ), .CI(\SUMB[27][64] ), 
        .CO(\CARRYB[28][63] ), .S(\SUMB[28][63] ) );
  FA1A S2_28_43 ( .A(\ab[28][43] ), .B(\CARRYB[27][43] ), .CI(\SUMB[27][44] ), 
        .CO(\CARRYB[28][43] ), .S(\SUMB[28][43] ) );
  FA1A S2_28_42 ( .A(\ab[28][42] ), .B(\CARRYB[27][42] ), .CI(\SUMB[27][43] ), 
        .CO(\CARRYB[28][42] ), .S(\SUMB[28][42] ) );
  FA1A S2_28_41 ( .A(\ab[28][41] ), .B(\CARRYB[27][41] ), .CI(\SUMB[27][42] ), 
        .CO(\CARRYB[28][41] ), .S(\SUMB[28][41] ) );
  FA1A S2_28_40 ( .A(\ab[28][40] ), .B(\CARRYB[27][40] ), .CI(\SUMB[27][41] ), 
        .CO(\CARRYB[28][40] ), .S(\SUMB[28][40] ) );
  FA1A S2_28_39 ( .A(\ab[28][39] ), .B(\CARRYB[27][39] ), .CI(\SUMB[27][40] ), 
        .CO(\CARRYB[28][39] ), .S(\SUMB[28][39] ) );
  FA1A S2_27_62 ( .A(\ab[27][62] ), .B(\CARRYB[26][62] ), .CI(\SUMB[26][63] ), 
        .CO(\CARRYB[27][62] ), .S(\SUMB[27][62] ) );
  FA1A S2_27_61 ( .A(\ab[27][61] ), .B(\CARRYB[26][61] ), .CI(\SUMB[26][62] ), 
        .CO(\CARRYB[27][61] ), .S(\SUMB[27][61] ) );
  FA1A S2_27_63 ( .A(\ab[27][63] ), .B(\CARRYB[26][63] ), .CI(\SUMB[26][64] ), 
        .CO(\CARRYB[27][63] ), .S(\SUMB[27][63] ) );
  FA1A S2_27_44 ( .A(\ab[27][44] ), .B(\CARRYB[26][44] ), .CI(\SUMB[26][45] ), 
        .CO(\CARRYB[27][44] ), .S(\SUMB[27][44] ) );
  FA1A S2_27_43 ( .A(\ab[27][43] ), .B(\CARRYB[26][43] ), .CI(\SUMB[26][44] ), 
        .CO(\CARRYB[27][43] ), .S(\SUMB[27][43] ) );
  FA1A S2_27_42 ( .A(\ab[27][42] ), .B(\CARRYB[26][42] ), .CI(\SUMB[26][43] ), 
        .CO(\CARRYB[27][42] ), .S(\SUMB[27][42] ) );
  FA1A S2_27_41 ( .A(\ab[27][41] ), .B(\CARRYB[26][41] ), .CI(\SUMB[26][42] ), 
        .CO(\CARRYB[27][41] ), .S(\SUMB[27][41] ) );
  FA1A S2_27_40 ( .A(\ab[27][40] ), .B(\CARRYB[26][40] ), .CI(\SUMB[26][41] ), 
        .CO(\CARRYB[27][40] ), .S(\SUMB[27][40] ) );
  FA1A S2_27_39 ( .A(\ab[27][39] ), .B(\CARRYB[26][39] ), .CI(\SUMB[26][40] ), 
        .CO(\CARRYB[27][39] ), .S(\SUMB[27][39] ) );
  FA1A S2_27_52 ( .A(\ab[27][52] ), .B(\CARRYB[26][52] ), .CI(\SUMB[26][53] ), 
        .CO(\CARRYB[27][52] ), .S(\SUMB[27][52] ) );
  FA1A S2_26_63 ( .A(\ab[26][63] ), .B(\CARRYB[25][63] ), .CI(\SUMB[25][64] ), 
        .CO(\CARRYB[26][63] ), .S(\SUMB[26][63] ) );
  FA1A S2_26_62 ( .A(\ab[26][62] ), .B(\CARRYB[25][62] ), .CI(\SUMB[25][63] ), 
        .CO(\CARRYB[26][62] ), .S(\SUMB[26][62] ) );
  FA1A S2_26_61 ( .A(\ab[26][61] ), .B(\CARRYB[25][61] ), .CI(\SUMB[25][62] ), 
        .CO(\CARRYB[26][61] ), .S(\SUMB[26][61] ) );
  FA1A S2_26_44 ( .A(\ab[26][44] ), .B(\CARRYB[25][44] ), .CI(\SUMB[25][45] ), 
        .CO(\CARRYB[26][44] ), .S(\SUMB[26][44] ) );
  FA1A S2_26_43 ( .A(\ab[26][43] ), .B(\CARRYB[25][43] ), .CI(\SUMB[25][44] ), 
        .CO(\CARRYB[26][43] ), .S(\SUMB[26][43] ) );
  FA1A S2_26_42 ( .A(\ab[26][42] ), .B(\CARRYB[25][42] ), .CI(\SUMB[25][43] ), 
        .CO(\CARRYB[26][42] ), .S(\SUMB[26][42] ) );
  FA1A S2_26_41 ( .A(\ab[26][41] ), .B(\CARRYB[25][41] ), .CI(\SUMB[25][42] ), 
        .CO(\CARRYB[26][41] ), .S(\SUMB[26][41] ) );
  FA1A S2_26_40 ( .A(\ab[26][40] ), .B(\CARRYB[25][40] ), .CI(\SUMB[25][41] ), 
        .CO(\CARRYB[26][40] ), .S(\SUMB[26][40] ) );
  FA1A S2_26_39 ( .A(\ab[26][39] ), .B(\CARRYB[25][39] ), .CI(\SUMB[25][40] ), 
        .CO(\CARRYB[26][39] ), .S(\SUMB[26][39] ) );
  FA1A S2_26_52 ( .A(\ab[26][52] ), .B(\CARRYB[25][52] ), .CI(\SUMB[25][53] ), 
        .CO(\CARRYB[26][52] ), .S(\SUMB[26][52] ) );
  FA1A S2_25_63 ( .A(\ab[25][63] ), .B(\CARRYB[24][63] ), .CI(\SUMB[24][64] ), 
        .CO(\CARRYB[25][63] ), .S(\SUMB[25][63] ) );
  FA1A S2_25_62 ( .A(\ab[25][62] ), .B(\CARRYB[24][62] ), .CI(\SUMB[24][63] ), 
        .CO(\CARRYB[25][62] ), .S(\SUMB[25][62] ) );
  FA1A S2_25_61 ( .A(\ab[25][61] ), .B(\CARRYB[24][61] ), .CI(\SUMB[24][62] ), 
        .CO(\CARRYB[25][61] ), .S(\SUMB[25][61] ) );
  FA1A S2_25_44 ( .A(\ab[25][44] ), .B(\CARRYB[24][44] ), .CI(\SUMB[24][45] ), 
        .CO(\CARRYB[25][44] ), .S(\SUMB[25][44] ) );
  FA1A S2_25_43 ( .A(\ab[25][43] ), .B(\CARRYB[24][43] ), .CI(\SUMB[24][44] ), 
        .CO(\CARRYB[25][43] ), .S(\SUMB[25][43] ) );
  FA1A S2_25_42 ( .A(\ab[25][42] ), .B(\CARRYB[24][42] ), .CI(\SUMB[24][43] ), 
        .CO(\CARRYB[25][42] ), .S(\SUMB[25][42] ) );
  FA1A S2_25_41 ( .A(\ab[25][41] ), .B(\CARRYB[24][41] ), .CI(\SUMB[24][42] ), 
        .CO(\CARRYB[25][41] ), .S(\SUMB[25][41] ) );
  FA1A S2_25_40 ( .A(\ab[25][40] ), .B(\CARRYB[24][40] ), .CI(\SUMB[24][41] ), 
        .CO(\CARRYB[25][40] ), .S(\SUMB[25][40] ) );
  FA1A S2_25_39 ( .A(\ab[25][39] ), .B(\CARRYB[24][39] ), .CI(\SUMB[24][40] ), 
        .CO(\CARRYB[25][39] ), .S(\SUMB[25][39] ) );
  FA1A S2_25_52 ( .A(\ab[25][52] ), .B(\CARRYB[24][52] ), .CI(\SUMB[24][53] ), 
        .CO(\CARRYB[25][52] ), .S(\SUMB[25][52] ) );
  FA1A S2_24_63 ( .A(\ab[24][63] ), .B(\CARRYB[23][63] ), .CI(\SUMB[23][64] ), 
        .CO(\CARRYB[24][63] ), .S(\SUMB[24][63] ) );
  FA1A S2_24_62 ( .A(\ab[24][62] ), .B(\CARRYB[23][62] ), .CI(\SUMB[23][63] ), 
        .CO(\CARRYB[24][62] ), .S(\SUMB[24][62] ) );
  FA1A S2_24_61 ( .A(\ab[24][61] ), .B(\CARRYB[23][61] ), .CI(\SUMB[23][62] ), 
        .CO(\CARRYB[24][61] ), .S(\SUMB[24][61] ) );
  FA1A S2_24_44 ( .A(\ab[24][44] ), .B(\CARRYB[23][44] ), .CI(\SUMB[23][45] ), 
        .CO(\CARRYB[24][44] ), .S(\SUMB[24][44] ) );
  FA1A S2_24_43 ( .A(\ab[24][43] ), .B(\CARRYB[23][43] ), .CI(\SUMB[23][44] ), 
        .CO(\CARRYB[24][43] ), .S(\SUMB[24][43] ) );
  FA1A S2_24_42 ( .A(\ab[24][42] ), .B(\CARRYB[23][42] ), .CI(\SUMB[23][43] ), 
        .CO(\CARRYB[24][42] ), .S(\SUMB[24][42] ) );
  FA1A S2_24_41 ( .A(\ab[24][41] ), .B(\CARRYB[23][41] ), .CI(\SUMB[23][42] ), 
        .CO(\CARRYB[24][41] ), .S(\SUMB[24][41] ) );
  FA1A S2_24_40 ( .A(\ab[24][40] ), .B(\CARRYB[23][40] ), .CI(\SUMB[23][41] ), 
        .CO(\CARRYB[24][40] ), .S(\SUMB[24][40] ) );
  FA1A S2_24_39 ( .A(\ab[24][39] ), .B(\CARRYB[23][39] ), .CI(\SUMB[23][40] ), 
        .CO(\CARRYB[24][39] ), .S(\SUMB[24][39] ) );
  FA1A S2_24_52 ( .A(\ab[24][52] ), .B(\CARRYB[23][52] ), .CI(\SUMB[23][53] ), 
        .CO(\CARRYB[24][52] ), .S(\SUMB[24][52] ) );
  FA1A S2_23_63 ( .A(\ab[23][63] ), .B(\CARRYB[22][63] ), .CI(\SUMB[22][64] ), 
        .CO(\CARRYB[23][63] ), .S(\SUMB[23][63] ) );
  FA1A S2_23_62 ( .A(\ab[23][62] ), .B(\CARRYB[22][62] ), .CI(\SUMB[22][63] ), 
        .CO(\CARRYB[23][62] ), .S(\SUMB[23][62] ) );
  FA1A S2_23_61 ( .A(\ab[23][61] ), .B(\CARRYB[22][61] ), .CI(\SUMB[22][62] ), 
        .CO(\CARRYB[23][61] ), .S(\SUMB[23][61] ) );
  FA1A S2_23_44 ( .A(\ab[23][44] ), .B(\CARRYB[22][44] ), .CI(\SUMB[22][45] ), 
        .CO(\CARRYB[23][44] ), .S(\SUMB[23][44] ) );
  FA1A S2_23_43 ( .A(\ab[23][43] ), .B(\CARRYB[22][43] ), .CI(\SUMB[22][44] ), 
        .CO(\CARRYB[23][43] ), .S(\SUMB[23][43] ) );
  FA1A S2_23_42 ( .A(\ab[23][42] ), .B(\CARRYB[22][42] ), .CI(\SUMB[22][43] ), 
        .CO(\CARRYB[23][42] ), .S(\SUMB[23][42] ) );
  FA1A S2_23_41 ( .A(\ab[23][41] ), .B(\CARRYB[22][41] ), .CI(\SUMB[22][42] ), 
        .CO(\CARRYB[23][41] ), .S(\SUMB[23][41] ) );
  FA1A S2_23_40 ( .A(\ab[23][40] ), .B(\CARRYB[22][40] ), .CI(\SUMB[22][41] ), 
        .CO(\CARRYB[23][40] ), .S(\SUMB[23][40] ) );
  FA1A S2_23_39 ( .A(\ab[23][39] ), .B(\CARRYB[22][39] ), .CI(\SUMB[22][40] ), 
        .CO(\CARRYB[23][39] ), .S(\SUMB[23][39] ) );
  FA1A S2_23_52 ( .A(\ab[23][52] ), .B(\CARRYB[22][52] ), .CI(\SUMB[22][53] ), 
        .CO(\CARRYB[23][52] ), .S(\SUMB[23][52] ) );
  FA1A S2_22_63 ( .A(\ab[22][63] ), .B(\CARRYB[21][63] ), .CI(\SUMB[21][64] ), 
        .CO(\CARRYB[22][63] ), .S(\SUMB[22][63] ) );
  FA1A S2_22_62 ( .A(\ab[22][62] ), .B(\CARRYB[21][62] ), .CI(\SUMB[21][63] ), 
        .CO(\CARRYB[22][62] ), .S(\SUMB[22][62] ) );
  FA1A S2_22_61 ( .A(\ab[22][61] ), .B(\CARRYB[21][61] ), .CI(\SUMB[21][62] ), 
        .CO(\CARRYB[22][61] ), .S(\SUMB[22][61] ) );
  FA1A S2_22_44 ( .A(\ab[22][44] ), .B(\CARRYB[21][44] ), .CI(\SUMB[21][45] ), 
        .CO(\CARRYB[22][44] ), .S(\SUMB[22][44] ) );
  FA1A S2_22_43 ( .A(\ab[22][43] ), .B(\CARRYB[21][43] ), .CI(\SUMB[21][44] ), 
        .CO(\CARRYB[22][43] ), .S(\SUMB[22][43] ) );
  FA1A S2_22_42 ( .A(\ab[22][42] ), .B(\CARRYB[21][42] ), .CI(\SUMB[21][43] ), 
        .CO(\CARRYB[22][42] ), .S(\SUMB[22][42] ) );
  FA1A S2_22_41 ( .A(\ab[22][41] ), .B(\CARRYB[21][41] ), .CI(\SUMB[21][42] ), 
        .CO(\CARRYB[22][41] ), .S(\SUMB[22][41] ) );
  FA1A S2_22_40 ( .A(\ab[22][40] ), .B(\CARRYB[21][40] ), .CI(\SUMB[21][41] ), 
        .CO(\CARRYB[22][40] ), .S(\SUMB[22][40] ) );
  FA1A S2_22_39 ( .A(\ab[22][39] ), .B(\CARRYB[21][39] ), .CI(\SUMB[21][40] ), 
        .CO(\CARRYB[22][39] ), .S(\SUMB[22][39] ) );
  FA1A S2_22_52 ( .A(\ab[22][52] ), .B(\CARRYB[21][52] ), .CI(\SUMB[21][53] ), 
        .CO(\CARRYB[22][52] ), .S(\SUMB[22][52] ) );
  FA1A S2_21_63 ( .A(\ab[21][63] ), .B(\CARRYB[20][63] ), .CI(\SUMB[20][64] ), 
        .CO(\CARRYB[21][63] ), .S(\SUMB[21][63] ) );
  FA1A S2_21_62 ( .A(\ab[21][62] ), .B(\CARRYB[20][62] ), .CI(\SUMB[20][63] ), 
        .CO(\CARRYB[21][62] ), .S(\SUMB[21][62] ) );
  FA1A S2_21_61 ( .A(\ab[21][61] ), .B(\CARRYB[20][61] ), .CI(\SUMB[20][62] ), 
        .CO(\CARRYB[21][61] ), .S(\SUMB[21][61] ) );
  FA1A S2_21_44 ( .A(\ab[21][44] ), .B(\CARRYB[20][44] ), .CI(\SUMB[20][45] ), 
        .CO(\CARRYB[21][44] ), .S(\SUMB[21][44] ) );
  FA1A S2_21_43 ( .A(\ab[21][43] ), .B(\CARRYB[20][43] ), .CI(\SUMB[20][44] ), 
        .CO(\CARRYB[21][43] ), .S(\SUMB[21][43] ) );
  FA1A S2_21_42 ( .A(\ab[21][42] ), .B(\CARRYB[20][42] ), .CI(\SUMB[20][43] ), 
        .CO(\CARRYB[21][42] ), .S(\SUMB[21][42] ) );
  FA1A S2_21_41 ( .A(\ab[21][41] ), .B(\CARRYB[20][41] ), .CI(\SUMB[20][42] ), 
        .CO(\CARRYB[21][41] ), .S(\SUMB[21][41] ) );
  FA1A S2_21_40 ( .A(\ab[21][40] ), .B(\CARRYB[20][40] ), .CI(\SUMB[20][41] ), 
        .CO(\CARRYB[21][40] ), .S(\SUMB[21][40] ) );
  FA1A S2_21_39 ( .A(\ab[21][39] ), .B(\CARRYB[20][39] ), .CI(\SUMB[20][40] ), 
        .CO(\CARRYB[21][39] ), .S(\SUMB[21][39] ) );
  FA1A S2_21_52 ( .A(\ab[21][52] ), .B(\CARRYB[20][52] ), .CI(\SUMB[20][53] ), 
        .CO(\CARRYB[21][52] ), .S(\SUMB[21][52] ) );
  FA1A S2_20_63 ( .A(\ab[20][63] ), .B(\CARRYB[19][63] ), .CI(\SUMB[19][64] ), 
        .CO(\CARRYB[20][63] ), .S(\SUMB[20][63] ) );
  FA1A S2_20_62 ( .A(\ab[20][62] ), .B(\CARRYB[19][62] ), .CI(\SUMB[19][63] ), 
        .CO(\CARRYB[20][62] ), .S(\SUMB[20][62] ) );
  FA1A S2_20_61 ( .A(\ab[20][61] ), .B(\CARRYB[19][61] ), .CI(\SUMB[19][62] ), 
        .CO(\CARRYB[20][61] ), .S(\SUMB[20][61] ) );
  FA1A S2_20_44 ( .A(\ab[20][44] ), .B(\CARRYB[19][44] ), .CI(\SUMB[19][45] ), 
        .CO(\CARRYB[20][44] ), .S(\SUMB[20][44] ) );
  FA1A S2_20_43 ( .A(\ab[20][43] ), .B(\CARRYB[19][43] ), .CI(\SUMB[19][44] ), 
        .CO(\CARRYB[20][43] ), .S(\SUMB[20][43] ) );
  FA1A S2_20_42 ( .A(\ab[20][42] ), .B(\CARRYB[19][42] ), .CI(\SUMB[19][43] ), 
        .CO(\CARRYB[20][42] ), .S(\SUMB[20][42] ) );
  FA1A S2_20_41 ( .A(\ab[20][41] ), .B(\CARRYB[19][41] ), .CI(\SUMB[19][42] ), 
        .CO(\CARRYB[20][41] ), .S(\SUMB[20][41] ) );
  FA1A S2_20_40 ( .A(\ab[20][40] ), .B(\CARRYB[19][40] ), .CI(\SUMB[19][41] ), 
        .CO(\CARRYB[20][40] ), .S(\SUMB[20][40] ) );
  FA1A S2_20_39 ( .A(\ab[20][39] ), .B(\CARRYB[19][39] ), .CI(\SUMB[19][40] ), 
        .CO(\CARRYB[20][39] ), .S(\SUMB[20][39] ) );
  FA1A S2_20_52 ( .A(\ab[20][52] ), .B(\CARRYB[19][52] ), .CI(\SUMB[19][53] ), 
        .CO(\CARRYB[20][52] ), .S(\SUMB[20][52] ) );
  FA1A S2_19_63 ( .A(\ab[19][63] ), .B(\CARRYB[18][63] ), .CI(\SUMB[18][64] ), 
        .CO(\CARRYB[19][63] ), .S(\SUMB[19][63] ) );
  FA1A S2_19_62 ( .A(\ab[19][62] ), .B(\CARRYB[18][62] ), .CI(\SUMB[18][63] ), 
        .CO(\CARRYB[19][62] ), .S(\SUMB[19][62] ) );
  FA1A S2_19_61 ( .A(\ab[19][61] ), .B(\CARRYB[18][61] ), .CI(\SUMB[18][62] ), 
        .CO(\CARRYB[19][61] ), .S(\SUMB[19][61] ) );
  FA1A S2_19_52 ( .A(\ab[19][52] ), .B(\CARRYB[18][52] ), .CI(\SUMB[18][53] ), 
        .CO(\CARRYB[19][52] ), .S(\SUMB[19][52] ) );
  FA1A S2_19_44 ( .A(\ab[19][44] ), .B(\CARRYB[18][44] ), .CI(\SUMB[18][45] ), 
        .CO(\CARRYB[19][44] ), .S(\SUMB[19][44] ) );
  FA1A S2_19_43 ( .A(\ab[19][43] ), .B(\CARRYB[18][43] ), .CI(\SUMB[18][44] ), 
        .CO(\CARRYB[19][43] ), .S(\SUMB[19][43] ) );
  FA1A S2_19_42 ( .A(\ab[19][42] ), .B(\CARRYB[18][42] ), .CI(\SUMB[18][43] ), 
        .CO(\CARRYB[19][42] ), .S(\SUMB[19][42] ) );
  FA1A S2_19_41 ( .A(\ab[19][41] ), .B(\CARRYB[18][41] ), .CI(\SUMB[18][42] ), 
        .CO(\CARRYB[19][41] ), .S(\SUMB[19][41] ) );
  FA1A S2_19_40 ( .A(\ab[19][40] ), .B(\CARRYB[18][40] ), .CI(\SUMB[18][41] ), 
        .CO(\CARRYB[19][40] ), .S(\SUMB[19][40] ) );
  FA1A S2_19_39 ( .A(\ab[19][39] ), .B(\CARRYB[18][39] ), .CI(\SUMB[18][40] ), 
        .CO(\CARRYB[19][39] ), .S(\SUMB[19][39] ) );
  FA1A S2_18_63 ( .A(\ab[18][63] ), .B(\CARRYB[17][63] ), .CI(\SUMB[17][64] ), 
        .CO(\CARRYB[18][63] ), .S(\SUMB[18][63] ) );
  FA1A S2_18_62 ( .A(\ab[18][62] ), .B(\CARRYB[17][62] ), .CI(\SUMB[17][63] ), 
        .CO(\CARRYB[18][62] ), .S(\SUMB[18][62] ) );
  FA1A S2_18_61 ( .A(\ab[18][61] ), .B(\CARRYB[17][61] ), .CI(\SUMB[17][62] ), 
        .CO(\CARRYB[18][61] ), .S(\SUMB[18][61] ) );
  FA1A S2_18_52 ( .A(\ab[18][52] ), .B(\CARRYB[17][52] ), .CI(\SUMB[17][53] ), 
        .CO(\CARRYB[18][52] ), .S(\SUMB[18][52] ) );
  FA1A S2_18_44 ( .A(\ab[18][44] ), .B(\CARRYB[17][44] ), .CI(\SUMB[17][45] ), 
        .CO(\CARRYB[18][44] ), .S(\SUMB[18][44] ) );
  FA1A S2_18_43 ( .A(\ab[18][43] ), .B(\CARRYB[17][43] ), .CI(\SUMB[17][44] ), 
        .CO(\CARRYB[18][43] ), .S(\SUMB[18][43] ) );
  FA1A S2_18_42 ( .A(\ab[18][42] ), .B(\CARRYB[17][42] ), .CI(\SUMB[17][43] ), 
        .CO(\CARRYB[18][42] ), .S(\SUMB[18][42] ) );
  FA1A S2_18_41 ( .A(\ab[18][41] ), .B(\CARRYB[17][41] ), .CI(\SUMB[17][42] ), 
        .CO(\CARRYB[18][41] ), .S(\SUMB[18][41] ) );
  FA1A S2_18_40 ( .A(\ab[18][40] ), .B(\CARRYB[17][40] ), .CI(\SUMB[17][41] ), 
        .CO(\CARRYB[18][40] ), .S(\SUMB[18][40] ) );
  FA1A S2_18_39 ( .A(\ab[18][39] ), .B(\CARRYB[17][39] ), .CI(\SUMB[17][40] ), 
        .CO(\CARRYB[18][39] ), .S(\SUMB[18][39] ) );
  FA1A S2_17_63 ( .A(\ab[17][63] ), .B(\CARRYB[16][63] ), .CI(\SUMB[16][64] ), 
        .CO(\CARRYB[17][63] ), .S(\SUMB[17][63] ) );
  FA1A S2_17_62 ( .A(\ab[17][62] ), .B(\CARRYB[16][62] ), .CI(\SUMB[16][63] ), 
        .CO(\CARRYB[17][62] ), .S(\SUMB[17][62] ) );
  FA1A S2_17_61 ( .A(\ab[17][61] ), .B(\CARRYB[16][61] ), .CI(\SUMB[16][62] ), 
        .CO(\CARRYB[17][61] ), .S(\SUMB[17][61] ) );
  FA1A S2_17_52 ( .A(\ab[17][52] ), .B(\CARRYB[16][52] ), .CI(\SUMB[16][53] ), 
        .CO(\CARRYB[17][52] ), .S(\SUMB[17][52] ) );
  FA1A S2_17_44 ( .A(\ab[17][44] ), .B(\CARRYB[16][44] ), .CI(\SUMB[16][45] ), 
        .CO(\CARRYB[17][44] ), .S(\SUMB[17][44] ) );
  FA1A S2_17_43 ( .A(\ab[17][43] ), .B(\CARRYB[16][43] ), .CI(\SUMB[16][44] ), 
        .CO(\CARRYB[17][43] ), .S(\SUMB[17][43] ) );
  FA1A S2_17_42 ( .A(\ab[17][42] ), .B(\CARRYB[16][42] ), .CI(\SUMB[16][43] ), 
        .CO(\CARRYB[17][42] ), .S(\SUMB[17][42] ) );
  FA1A S2_17_41 ( .A(\ab[17][41] ), .B(\CARRYB[16][41] ), .CI(\SUMB[16][42] ), 
        .CO(\CARRYB[17][41] ), .S(\SUMB[17][41] ) );
  FA1A S2_17_40 ( .A(\ab[17][40] ), .B(\CARRYB[16][40] ), .CI(\SUMB[16][41] ), 
        .CO(\CARRYB[17][40] ), .S(\SUMB[17][40] ) );
  FA1A S2_17_39 ( .A(\ab[17][39] ), .B(\CARRYB[16][39] ), .CI(\SUMB[16][40] ), 
        .CO(\CARRYB[17][39] ), .S(\SUMB[17][39] ) );
  FA1A S2_16_63 ( .A(\ab[16][63] ), .B(\CARRYB[15][63] ), .CI(\SUMB[15][64] ), 
        .CO(\CARRYB[16][63] ), .S(\SUMB[16][63] ) );
  FA1A S2_16_62 ( .A(\ab[16][62] ), .B(\CARRYB[15][62] ), .CI(\SUMB[15][63] ), 
        .CO(\CARRYB[16][62] ), .S(\SUMB[16][62] ) );
  FA1A S2_16_61 ( .A(\ab[16][61] ), .B(\CARRYB[15][61] ), .CI(\SUMB[15][62] ), 
        .CO(\CARRYB[16][61] ), .S(\SUMB[16][61] ) );
  FA1A S2_16_52 ( .A(\ab[16][52] ), .B(\CARRYB[15][52] ), .CI(\SUMB[15][53] ), 
        .CO(\CARRYB[16][52] ), .S(\SUMB[16][52] ) );
  FA1A S2_16_44 ( .A(\ab[16][44] ), .B(\CARRYB[15][44] ), .CI(\SUMB[15][45] ), 
        .CO(\CARRYB[16][44] ), .S(\SUMB[16][44] ) );
  FA1A S2_16_43 ( .A(\ab[16][43] ), .B(\CARRYB[15][43] ), .CI(\SUMB[15][44] ), 
        .CO(\CARRYB[16][43] ), .S(\SUMB[16][43] ) );
  FA1A S2_16_42 ( .A(\ab[16][42] ), .B(\CARRYB[15][42] ), .CI(\SUMB[15][43] ), 
        .CO(\CARRYB[16][42] ), .S(\SUMB[16][42] ) );
  FA1A S2_16_41 ( .A(\ab[16][41] ), .B(\CARRYB[15][41] ), .CI(\SUMB[15][42] ), 
        .CO(\CARRYB[16][41] ), .S(\SUMB[16][41] ) );
  FA1A S2_16_40 ( .A(\ab[16][40] ), .B(\CARRYB[15][40] ), .CI(\SUMB[15][41] ), 
        .CO(\CARRYB[16][40] ), .S(\SUMB[16][40] ) );
  FA1A S2_16_39 ( .A(\ab[16][39] ), .B(\CARRYB[15][39] ), .CI(\SUMB[15][40] ), 
        .CO(\CARRYB[16][39] ), .S(\SUMB[16][39] ) );
  FA1A S2_15_63 ( .A(\ab[15][63] ), .B(\CARRYB[14][63] ), .CI(\SUMB[14][64] ), 
        .CO(\CARRYB[15][63] ), .S(\SUMB[15][63] ) );
  FA1A S2_15_62 ( .A(\ab[15][62] ), .B(\CARRYB[14][62] ), .CI(\SUMB[14][63] ), 
        .CO(\CARRYB[15][62] ), .S(\SUMB[15][62] ) );
  FA1A S2_15_61 ( .A(\ab[15][61] ), .B(\CARRYB[14][61] ), .CI(\SUMB[14][62] ), 
        .CO(\CARRYB[15][61] ), .S(\SUMB[15][61] ) );
  FA1A S2_15_52 ( .A(\ab[15][52] ), .B(\CARRYB[14][52] ), .CI(\SUMB[14][53] ), 
        .CO(\CARRYB[15][52] ), .S(\SUMB[15][52] ) );
  FA1A S2_15_44 ( .A(\ab[15][44] ), .B(\CARRYB[14][44] ), .CI(\SUMB[14][45] ), 
        .CO(\CARRYB[15][44] ), .S(\SUMB[15][44] ) );
  FA1A S2_15_43 ( .A(\ab[15][43] ), .B(\CARRYB[14][43] ), .CI(\SUMB[14][44] ), 
        .CO(\CARRYB[15][43] ), .S(\SUMB[15][43] ) );
  FA1A S2_15_42 ( .A(\ab[15][42] ), .B(\CARRYB[14][42] ), .CI(\SUMB[14][43] ), 
        .CO(\CARRYB[15][42] ), .S(\SUMB[15][42] ) );
  FA1A S2_15_41 ( .A(\ab[15][41] ), .B(\CARRYB[14][41] ), .CI(\SUMB[14][42] ), 
        .CO(\CARRYB[15][41] ), .S(\SUMB[15][41] ) );
  FA1A S2_15_40 ( .A(\ab[15][40] ), .B(\CARRYB[14][40] ), .CI(\SUMB[14][41] ), 
        .CO(\CARRYB[15][40] ), .S(\SUMB[15][40] ) );
  FA1A S2_15_38 ( .A(\ab[15][38] ), .B(\CARRYB[14][38] ), .CI(\SUMB[14][39] ), 
        .CO(\CARRYB[15][38] ), .S(\SUMB[15][38] ) );
  FA1A S2_15_39 ( .A(\ab[15][39] ), .B(\CARRYB[14][39] ), .CI(\SUMB[14][40] ), 
        .CO(\CARRYB[15][39] ), .S(\SUMB[15][39] ) );
  FA1A S2_14_38 ( .A(\ab[14][38] ), .B(\CARRYB[13][38] ), .CI(\SUMB[13][39] ), 
        .CO(\CARRYB[14][38] ), .S(\SUMB[14][38] ) );
  FA1A S2_13_38 ( .A(\ab[13][38] ), .B(\CARRYB[12][38] ), .CI(\SUMB[12][39] ), 
        .CO(\CARRYB[13][38] ), .S(\SUMB[13][38] ) );
  FA1A S2_12_38 ( .A(\ab[12][38] ), .B(\CARRYB[11][38] ), .CI(\SUMB[11][39] ), 
        .CO(\CARRYB[12][38] ), .S(\SUMB[12][38] ) );
  FA1A S2_11_38 ( .A(\ab[11][38] ), .B(\CARRYB[10][38] ), .CI(\SUMB[10][39] ), 
        .CO(\CARRYB[11][38] ), .S(\SUMB[11][38] ) );
  FA1A S2_10_38 ( .A(\ab[10][38] ), .B(\CARRYB[9][38] ), .CI(\SUMB[9][39] ), 
        .CO(\CARRYB[10][38] ), .S(\SUMB[10][38] ) );
  FA1A S2_9_38 ( .A(\ab[9][38] ), .B(\CARRYB[8][38] ), .CI(\SUMB[8][39] ), 
        .CO(\CARRYB[9][38] ), .S(\SUMB[9][38] ) );
  FA1A S2_8_38 ( .A(\ab[8][38] ), .B(\CARRYB[7][38] ), .CI(\SUMB[7][39] ), 
        .CO(\CARRYB[8][38] ), .S(\SUMB[8][38] ) );
  FA1A S2_7_38 ( .A(\ab[7][38] ), .B(\CARRYB[6][38] ), .CI(\SUMB[6][39] ), 
        .CO(\CARRYB[7][38] ), .S(\SUMB[7][38] ) );
  FA1A S2_6_38 ( .A(\ab[6][38] ), .B(\CARRYB[5][38] ), .CI(\SUMB[5][39] ), 
        .CO(\CARRYB[6][38] ), .S(\SUMB[6][38] ) );
  FA1A S2_5_38 ( .A(\ab[5][38] ), .B(\CARRYB[4][38] ), .CI(\SUMB[4][39] ), 
        .CO(\CARRYB[5][38] ), .S(\SUMB[5][38] ) );
  FA1A S2_4_38 ( .A(\ab[4][38] ), .B(\CARRYB[3][38] ), .CI(\SUMB[3][39] ), 
        .CO(\CARRYB[4][38] ), .S(\SUMB[4][38] ) );
  FA1A S2_3_38 ( .A(\ab[3][38] ), .B(\CARRYB[2][38] ), .CI(\SUMB[2][39] ), 
        .CO(\CARRYB[3][38] ), .S(\SUMB[3][38] ) );
  FA1A S2_2_38 ( .A(\ab[2][38] ), .B(\CARRYB[1][38] ), .CI(\SUMB[1][39] ), 
        .CO(\CARRYB[2][38] ), .S(\SUMB[2][38] ) );
  FA1A S2_2_37 ( .A(\ab[2][37] ), .B(\CARRYB[1][37] ), .CI(\SUMB[1][38] ), 
        .CO(\CARRYB[2][37] ), .S(\SUMB[2][37] ) );
  FA1A S4_52 ( .A(\ab[29][52] ), .B(\CARRYB[28][52] ), .CI(\SUMB[28][53] ), 
        .CO(\CARRYB[29][52] ), .S(\SUMB[29][52] ) );
  FA1A S4_63 ( .A(\ab[29][63] ), .B(\CARRYB[28][63] ), .CI(\SUMB[28][64] ), 
        .CO(\CARRYB[29][63] ), .S(\SUMB[29][63] ) );
  FA1A S4_47 ( .A(\ab[29][47] ), .B(\CARRYB[28][47] ), .CI(\SUMB[28][48] ), 
        .CO(\CARRYB[29][47] ), .S(\SUMB[29][47] ) );
  FA1A S4_46 ( .A(\ab[29][46] ), .B(\CARRYB[28][46] ), .CI(\SUMB[28][47] ), 
        .CO(\CARRYB[29][46] ), .S(\SUMB[29][46] ) );
  FA1A S2_28_47 ( .A(\ab[28][47] ), .B(\CARRYB[27][47] ), .CI(\SUMB[27][48] ), 
        .CO(\CARRYB[28][47] ), .S(\SUMB[28][47] ) );
  FA1A S4_49 ( .A(\ab[29][49] ), .B(\CARRYB[28][49] ), .CI(\SUMB[28][50] ), 
        .CO(\CARRYB[29][49] ), .S(\SUMB[29][49] ) );
  FA1A S4_50 ( .A(\ab[29][50] ), .B(\CARRYB[28][50] ), .CI(\SUMB[28][51] ), 
        .CO(\CARRYB[29][50] ), .S(\SUMB[29][50] ) );
  FA1A S4_45 ( .A(\ab[29][45] ), .B(\CARRYB[28][45] ), .CI(\SUMB[28][46] ), 
        .CO(\CARRYB[29][45] ), .S(\SUMB[29][45] ) );
  FA1A S2_28_49 ( .A(\ab[28][49] ), .B(\CARRYB[27][49] ), .CI(\SUMB[27][50] ), 
        .CO(\CARRYB[28][49] ), .S(\SUMB[28][49] ) );
  FA1A S2_28_48 ( .A(\ab[28][48] ), .B(\CARRYB[27][48] ), .CI(\SUMB[27][49] ), 
        .CO(\CARRYB[28][48] ), .S(\SUMB[28][48] ) );
  FA1A S2_28_50 ( .A(\ab[28][50] ), .B(\CARRYB[27][50] ), .CI(\SUMB[27][51] ), 
        .CO(\CARRYB[28][50] ), .S(\SUMB[28][50] ) );
  FA1A S2_28_51 ( .A(\ab[28][51] ), .B(\CARRYB[27][51] ), .CI(\SUMB[27][52] ), 
        .CO(\CARRYB[28][51] ), .S(\SUMB[28][51] ) );
  FA1A S2_28_46 ( .A(\ab[28][46] ), .B(\CARRYB[27][46] ), .CI(\SUMB[27][47] ), 
        .CO(\CARRYB[28][46] ), .S(\SUMB[28][46] ) );
  FA1A S2_28_45 ( .A(\ab[28][45] ), .B(\CARRYB[27][45] ), .CI(\SUMB[27][46] ), 
        .CO(\CARRYB[28][45] ), .S(\SUMB[28][45] ) );
  FA1A S2_27_50 ( .A(\ab[27][50] ), .B(\CARRYB[26][50] ), .CI(\SUMB[26][51] ), 
        .CO(\CARRYB[27][50] ), .S(\SUMB[27][50] ) );
  FA1A S2_27_49 ( .A(\ab[27][49] ), .B(\CARRYB[26][49] ), .CI(\SUMB[26][50] ), 
        .CO(\CARRYB[27][49] ), .S(\SUMB[27][49] ) );
  FA1A S2_27_48 ( .A(\ab[27][48] ), .B(\CARRYB[26][48] ), .CI(\SUMB[26][49] ), 
        .CO(\CARRYB[27][48] ), .S(\SUMB[27][48] ) );
  FA1A S2_27_51 ( .A(\ab[27][51] ), .B(\CARRYB[26][51] ), .CI(\SUMB[26][52] ), 
        .CO(\CARRYB[27][51] ), .S(\SUMB[27][51] ) );
  FA1A S2_27_47 ( .A(\ab[27][47] ), .B(\CARRYB[26][47] ), .CI(\SUMB[26][48] ), 
        .CO(\CARRYB[27][47] ), .S(\SUMB[27][47] ) );
  FA1A S2_27_46 ( .A(\ab[27][46] ), .B(\CARRYB[26][46] ), .CI(\SUMB[26][47] ), 
        .CO(\CARRYB[27][46] ), .S(\SUMB[27][46] ) );
  FA1A S2_27_45 ( .A(\ab[27][45] ), .B(\CARRYB[26][45] ), .CI(\SUMB[26][46] ), 
        .CO(\CARRYB[27][45] ), .S(\SUMB[27][45] ) );
  FA1A S2_26_45 ( .A(\ab[26][45] ), .B(\CARRYB[25][45] ), .CI(\SUMB[25][46] ), 
        .CO(\CARRYB[26][45] ), .S(\SUMB[26][45] ) );
  FA1A S2_26_51 ( .A(\ab[26][51] ), .B(\CARRYB[25][51] ), .CI(\SUMB[25][52] ), 
        .CO(\CARRYB[26][51] ), .S(\SUMB[26][51] ) );
  FA1A S2_26_50 ( .A(\ab[26][50] ), .B(\CARRYB[25][50] ), .CI(\SUMB[25][51] ), 
        .CO(\CARRYB[26][50] ), .S(\SUMB[26][50] ) );
  FA1A S2_26_49 ( .A(\ab[26][49] ), .B(\CARRYB[25][49] ), .CI(\SUMB[25][50] ), 
        .CO(\CARRYB[26][49] ), .S(\SUMB[26][49] ) );
  FA1A S2_26_48 ( .A(\ab[26][48] ), .B(\CARRYB[25][48] ), .CI(\SUMB[25][49] ), 
        .CO(\CARRYB[26][48] ), .S(\SUMB[26][48] ) );
  FA1A S2_26_47 ( .A(\ab[26][47] ), .B(\CARRYB[25][47] ), .CI(\SUMB[25][48] ), 
        .CO(\CARRYB[26][47] ), .S(\SUMB[26][47] ) );
  FA1A S2_26_46 ( .A(\ab[26][46] ), .B(\CARRYB[25][46] ), .CI(\SUMB[25][47] ), 
        .CO(\CARRYB[26][46] ), .S(\SUMB[26][46] ) );
  FA1A S2_25_46 ( .A(\ab[25][46] ), .B(\CARRYB[24][46] ), .CI(\SUMB[24][47] ), 
        .CO(\CARRYB[25][46] ), .S(\SUMB[25][46] ) );
  FA1A S2_25_45 ( .A(\ab[25][45] ), .B(\CARRYB[24][45] ), .CI(\SUMB[24][46] ), 
        .CO(\CARRYB[25][45] ), .S(\SUMB[25][45] ) );
  FA1A S2_25_51 ( .A(\ab[25][51] ), .B(\CARRYB[24][51] ), .CI(\SUMB[24][52] ), 
        .CO(\CARRYB[25][51] ), .S(\SUMB[25][51] ) );
  FA1A S2_25_50 ( .A(\ab[25][50] ), .B(\CARRYB[24][50] ), .CI(\SUMB[24][51] ), 
        .CO(\CARRYB[25][50] ), .S(\SUMB[25][50] ) );
  FA1A S2_25_49 ( .A(\ab[25][49] ), .B(\CARRYB[24][49] ), .CI(\SUMB[24][50] ), 
        .CO(\CARRYB[25][49] ), .S(\SUMB[25][49] ) );
  FA1A S2_25_48 ( .A(\ab[25][48] ), .B(\CARRYB[24][48] ), .CI(\SUMB[24][49] ), 
        .CO(\CARRYB[25][48] ), .S(\SUMB[25][48] ) );
  FA1A S2_25_47 ( .A(\ab[25][47] ), .B(\CARRYB[24][47] ), .CI(\SUMB[24][48] ), 
        .CO(\CARRYB[25][47] ), .S(\SUMB[25][47] ) );
  FA1A S2_24_47 ( .A(\ab[24][47] ), .B(\CARRYB[23][47] ), .CI(\SUMB[23][48] ), 
        .CO(\CARRYB[24][47] ), .S(\SUMB[24][47] ) );
  FA1A S2_24_46 ( .A(\ab[24][46] ), .B(\CARRYB[23][46] ), .CI(\SUMB[23][47] ), 
        .CO(\CARRYB[24][46] ), .S(\SUMB[24][46] ) );
  FA1A S2_24_45 ( .A(\ab[24][45] ), .B(\CARRYB[23][45] ), .CI(\SUMB[23][46] ), 
        .CO(\CARRYB[24][45] ), .S(\SUMB[24][45] ) );
  FA1A S2_24_51 ( .A(\ab[24][51] ), .B(\CARRYB[23][51] ), .CI(\SUMB[23][52] ), 
        .CO(\CARRYB[24][51] ), .S(\SUMB[24][51] ) );
  FA1A S2_24_50 ( .A(\ab[24][50] ), .B(\CARRYB[23][50] ), .CI(\SUMB[23][51] ), 
        .CO(\CARRYB[24][50] ), .S(\SUMB[24][50] ) );
  FA1A S2_24_49 ( .A(\ab[24][49] ), .B(\CARRYB[23][49] ), .CI(\SUMB[23][50] ), 
        .CO(\CARRYB[24][49] ), .S(\SUMB[24][49] ) );
  FA1A S2_24_48 ( .A(\ab[24][48] ), .B(\CARRYB[23][48] ), .CI(\SUMB[23][49] ), 
        .CO(\CARRYB[24][48] ), .S(\SUMB[24][48] ) );
  FA1A S2_23_48 ( .A(\ab[23][48] ), .B(\CARRYB[22][48] ), .CI(\SUMB[22][49] ), 
        .CO(\CARRYB[23][48] ), .S(\SUMB[23][48] ) );
  FA1A S2_23_47 ( .A(\ab[23][47] ), .B(\CARRYB[22][47] ), .CI(\SUMB[22][48] ), 
        .CO(\CARRYB[23][47] ), .S(\SUMB[23][47] ) );
  FA1A S2_23_46 ( .A(\ab[23][46] ), .B(\CARRYB[22][46] ), .CI(\SUMB[22][47] ), 
        .CO(\CARRYB[23][46] ), .S(\SUMB[23][46] ) );
  FA1A S2_23_45 ( .A(\ab[23][45] ), .B(\CARRYB[22][45] ), .CI(\SUMB[22][46] ), 
        .CO(\CARRYB[23][45] ), .S(\SUMB[23][45] ) );
  FA1A S2_23_51 ( .A(\ab[23][51] ), .B(\CARRYB[22][51] ), .CI(\SUMB[22][52] ), 
        .CO(\CARRYB[23][51] ), .S(\SUMB[23][51] ) );
  FA1A S2_23_50 ( .A(\ab[23][50] ), .B(\CARRYB[22][50] ), .CI(\SUMB[22][51] ), 
        .CO(\CARRYB[23][50] ), .S(\SUMB[23][50] ) );
  FA1A S2_23_49 ( .A(\ab[23][49] ), .B(\CARRYB[22][49] ), .CI(\SUMB[22][50] ), 
        .CO(\CARRYB[23][49] ), .S(\SUMB[23][49] ) );
  FA1A S2_22_49 ( .A(\ab[22][49] ), .B(\CARRYB[21][49] ), .CI(\SUMB[21][50] ), 
        .CO(\CARRYB[22][49] ), .S(\SUMB[22][49] ) );
  FA1A S2_22_48 ( .A(\ab[22][48] ), .B(\CARRYB[21][48] ), .CI(\SUMB[21][49] ), 
        .CO(\CARRYB[22][48] ), .S(\SUMB[22][48] ) );
  FA1A S2_22_47 ( .A(\ab[22][47] ), .B(\CARRYB[21][47] ), .CI(\SUMB[21][48] ), 
        .CO(\CARRYB[22][47] ), .S(\SUMB[22][47] ) );
  FA1A S2_22_46 ( .A(\ab[22][46] ), .B(\CARRYB[21][46] ), .CI(\SUMB[21][47] ), 
        .CO(\CARRYB[22][46] ), .S(\SUMB[22][46] ) );
  FA1A S2_22_45 ( .A(\ab[22][45] ), .B(\CARRYB[21][45] ), .CI(\SUMB[21][46] ), 
        .CO(\CARRYB[22][45] ), .S(\SUMB[22][45] ) );
  FA1A S2_22_51 ( .A(\ab[22][51] ), .B(\CARRYB[21][51] ), .CI(\SUMB[21][52] ), 
        .CO(\CARRYB[22][51] ), .S(\SUMB[22][51] ) );
  FA1A S2_22_50 ( .A(\ab[22][50] ), .B(\CARRYB[21][50] ), .CI(\SUMB[21][51] ), 
        .CO(\CARRYB[22][50] ), .S(\SUMB[22][50] ) );
  FA1A S2_21_50 ( .A(\ab[21][50] ), .B(\CARRYB[20][50] ), .CI(\SUMB[20][51] ), 
        .CO(\CARRYB[21][50] ), .S(\SUMB[21][50] ) );
  FA1A S2_21_49 ( .A(\ab[21][49] ), .B(\CARRYB[20][49] ), .CI(\SUMB[20][50] ), 
        .CO(\CARRYB[21][49] ), .S(\SUMB[21][49] ) );
  FA1A S2_21_48 ( .A(\ab[21][48] ), .B(\CARRYB[20][48] ), .CI(\SUMB[20][49] ), 
        .CO(\CARRYB[21][48] ), .S(\SUMB[21][48] ) );
  FA1A S2_21_47 ( .A(\ab[21][47] ), .B(\CARRYB[20][47] ), .CI(\SUMB[20][48] ), 
        .CO(\CARRYB[21][47] ), .S(\SUMB[21][47] ) );
  FA1A S2_21_46 ( .A(\ab[21][46] ), .B(\CARRYB[20][46] ), .CI(\SUMB[20][47] ), 
        .CO(\CARRYB[21][46] ), .S(\SUMB[21][46] ) );
  FA1A S2_21_45 ( .A(\ab[21][45] ), .B(\CARRYB[20][45] ), .CI(\SUMB[20][46] ), 
        .CO(\CARRYB[21][45] ), .S(\SUMB[21][45] ) );
  FA1A S2_21_51 ( .A(\ab[21][51] ), .B(\CARRYB[20][51] ), .CI(\SUMB[20][52] ), 
        .CO(\CARRYB[21][51] ), .S(\SUMB[21][51] ) );
  FA1A S2_20_51 ( .A(\ab[20][51] ), .B(\CARRYB[19][51] ), .CI(\SUMB[19][52] ), 
        .CO(\CARRYB[20][51] ), .S(\SUMB[20][51] ) );
  FA1A S2_20_50 ( .A(\ab[20][50] ), .B(\CARRYB[19][50] ), .CI(\SUMB[19][51] ), 
        .CO(\CARRYB[20][50] ), .S(\SUMB[20][50] ) );
  FA1A S2_20_49 ( .A(\ab[20][49] ), .B(\CARRYB[19][49] ), .CI(\SUMB[19][50] ), 
        .CO(\CARRYB[20][49] ), .S(\SUMB[20][49] ) );
  FA1A S2_20_48 ( .A(\ab[20][48] ), .B(\CARRYB[19][48] ), .CI(\SUMB[19][49] ), 
        .CO(\CARRYB[20][48] ), .S(\SUMB[20][48] ) );
  FA1A S2_20_47 ( .A(\ab[20][47] ), .B(\CARRYB[19][47] ), .CI(\SUMB[19][48] ), 
        .CO(\CARRYB[20][47] ), .S(\SUMB[20][47] ) );
  FA1A S2_20_46 ( .A(\ab[20][46] ), .B(\CARRYB[19][46] ), .CI(\SUMB[19][47] ), 
        .CO(\CARRYB[20][46] ), .S(\SUMB[20][46] ) );
  FA1A S2_20_45 ( .A(\ab[20][45] ), .B(\CARRYB[19][45] ), .CI(\SUMB[19][46] ), 
        .CO(\CARRYB[20][45] ), .S(\SUMB[20][45] ) );
  FA1A S2_19_51 ( .A(\ab[19][51] ), .B(\CARRYB[18][51] ), .CI(\SUMB[18][52] ), 
        .CO(\CARRYB[19][51] ), .S(\SUMB[19][51] ) );
  FA1A S2_19_50 ( .A(\ab[19][50] ), .B(\CARRYB[18][50] ), .CI(\SUMB[18][51] ), 
        .CO(\CARRYB[19][50] ), .S(\SUMB[19][50] ) );
  FA1A S2_19_49 ( .A(\ab[19][49] ), .B(\CARRYB[18][49] ), .CI(\SUMB[18][50] ), 
        .CO(\CARRYB[19][49] ), .S(\SUMB[19][49] ) );
  FA1A S2_19_48 ( .A(\ab[19][48] ), .B(\CARRYB[18][48] ), .CI(\SUMB[18][49] ), 
        .CO(\CARRYB[19][48] ), .S(\SUMB[19][48] ) );
  FA1A S2_19_47 ( .A(\ab[19][47] ), .B(\CARRYB[18][47] ), .CI(\SUMB[18][48] ), 
        .CO(\CARRYB[19][47] ), .S(\SUMB[19][47] ) );
  FA1A S2_19_46 ( .A(\ab[19][46] ), .B(\CARRYB[18][46] ), .CI(\SUMB[18][47] ), 
        .CO(\CARRYB[19][46] ), .S(\SUMB[19][46] ) );
  FA1A S2_19_45 ( .A(\ab[19][45] ), .B(\CARRYB[18][45] ), .CI(\SUMB[18][46] ), 
        .CO(\CARRYB[19][45] ), .S(\SUMB[19][45] ) );
  FA1A S2_18_51 ( .A(\ab[18][51] ), .B(\CARRYB[17][51] ), .CI(\SUMB[17][52] ), 
        .CO(\CARRYB[18][51] ), .S(\SUMB[18][51] ) );
  FA1A S2_18_50 ( .A(\ab[18][50] ), .B(\CARRYB[17][50] ), .CI(\SUMB[17][51] ), 
        .CO(\CARRYB[18][50] ), .S(\SUMB[18][50] ) );
  FA1A S2_18_49 ( .A(\ab[18][49] ), .B(\CARRYB[17][49] ), .CI(\SUMB[17][50] ), 
        .CO(\CARRYB[18][49] ), .S(\SUMB[18][49] ) );
  FA1A S2_18_48 ( .A(\ab[18][48] ), .B(\CARRYB[17][48] ), .CI(\SUMB[17][49] ), 
        .CO(\CARRYB[18][48] ), .S(\SUMB[18][48] ) );
  FA1A S2_18_47 ( .A(\ab[18][47] ), .B(\CARRYB[17][47] ), .CI(\SUMB[17][48] ), 
        .CO(\CARRYB[18][47] ), .S(\SUMB[18][47] ) );
  FA1A S2_18_46 ( .A(\ab[18][46] ), .B(\CARRYB[17][46] ), .CI(\SUMB[17][47] ), 
        .CO(\CARRYB[18][46] ), .S(\SUMB[18][46] ) );
  FA1A S2_18_45 ( .A(\ab[18][45] ), .B(\CARRYB[17][45] ), .CI(\SUMB[17][46] ), 
        .CO(\CARRYB[18][45] ), .S(\SUMB[18][45] ) );
  FA1A S2_17_51 ( .A(\ab[17][51] ), .B(\CARRYB[16][51] ), .CI(\SUMB[16][52] ), 
        .CO(\CARRYB[17][51] ), .S(\SUMB[17][51] ) );
  FA1A S2_17_50 ( .A(\ab[17][50] ), .B(\CARRYB[16][50] ), .CI(\SUMB[16][51] ), 
        .CO(\CARRYB[17][50] ), .S(\SUMB[17][50] ) );
  FA1A S2_17_49 ( .A(\ab[17][49] ), .B(\CARRYB[16][49] ), .CI(\SUMB[16][50] ), 
        .CO(\CARRYB[17][49] ), .S(\SUMB[17][49] ) );
  FA1A S2_17_48 ( .A(\ab[17][48] ), .B(\CARRYB[16][48] ), .CI(\SUMB[16][49] ), 
        .CO(\CARRYB[17][48] ), .S(\SUMB[17][48] ) );
  FA1A S2_17_47 ( .A(\ab[17][47] ), .B(\CARRYB[16][47] ), .CI(\SUMB[16][48] ), 
        .CO(\CARRYB[17][47] ), .S(\SUMB[17][47] ) );
  FA1A S2_17_46 ( .A(\ab[17][46] ), .B(\CARRYB[16][46] ), .CI(\SUMB[16][47] ), 
        .CO(\CARRYB[17][46] ), .S(\SUMB[17][46] ) );
  FA1A S2_17_45 ( .A(\ab[17][45] ), .B(\CARRYB[16][45] ), .CI(\SUMB[16][46] ), 
        .CO(\CARRYB[17][45] ), .S(\SUMB[17][45] ) );
  FA1A S2_16_51 ( .A(\ab[16][51] ), .B(\CARRYB[15][51] ), .CI(\SUMB[15][52] ), 
        .CO(\CARRYB[16][51] ), .S(\SUMB[16][51] ) );
  FA1A S2_16_50 ( .A(\ab[16][50] ), .B(\CARRYB[15][50] ), .CI(\SUMB[15][51] ), 
        .CO(\CARRYB[16][50] ), .S(\SUMB[16][50] ) );
  FA1A S2_16_49 ( .A(\ab[16][49] ), .B(\CARRYB[15][49] ), .CI(\SUMB[15][50] ), 
        .CO(\CARRYB[16][49] ), .S(\SUMB[16][49] ) );
  FA1A S2_16_48 ( .A(\ab[16][48] ), .B(\CARRYB[15][48] ), .CI(\SUMB[15][49] ), 
        .CO(\CARRYB[16][48] ), .S(\SUMB[16][48] ) );
  FA1A S2_16_47 ( .A(\ab[16][47] ), .B(\CARRYB[15][47] ), .CI(\SUMB[15][48] ), 
        .CO(\CARRYB[16][47] ), .S(\SUMB[16][47] ) );
  FA1A S2_16_46 ( .A(\ab[16][46] ), .B(\CARRYB[15][46] ), .CI(\SUMB[15][47] ), 
        .CO(\CARRYB[16][46] ), .S(\SUMB[16][46] ) );
  FA1A S2_16_45 ( .A(\ab[16][45] ), .B(\CARRYB[15][45] ), .CI(\SUMB[15][46] ), 
        .CO(\CARRYB[16][45] ), .S(\SUMB[16][45] ) );
  FA1A S2_15_51 ( .A(\ab[15][51] ), .B(\CARRYB[14][51] ), .CI(\SUMB[14][52] ), 
        .CO(\CARRYB[15][51] ), .S(\SUMB[15][51] ) );
  FA1A S2_15_50 ( .A(\ab[15][50] ), .B(\CARRYB[14][50] ), .CI(\SUMB[14][51] ), 
        .CO(\CARRYB[15][50] ), .S(\SUMB[15][50] ) );
  FA1A S2_15_49 ( .A(\ab[15][49] ), .B(\CARRYB[14][49] ), .CI(\SUMB[14][50] ), 
        .CO(\CARRYB[15][49] ), .S(\SUMB[15][49] ) );
  FA1A S2_15_48 ( .A(\ab[15][48] ), .B(\CARRYB[14][48] ), .CI(\SUMB[14][49] ), 
        .CO(\CARRYB[15][48] ), .S(\SUMB[15][48] ) );
  FA1A S2_15_47 ( .A(\ab[15][47] ), .B(\CARRYB[14][47] ), .CI(\SUMB[14][48] ), 
        .CO(\CARRYB[15][47] ), .S(\SUMB[15][47] ) );
  FA1A S2_15_46 ( .A(\ab[15][46] ), .B(\CARRYB[14][46] ), .CI(\SUMB[14][47] ), 
        .CO(\CARRYB[15][46] ), .S(\SUMB[15][46] ) );
  FA1A S2_15_45 ( .A(\ab[15][45] ), .B(\CARRYB[14][45] ), .CI(\SUMB[14][46] ), 
        .CO(\CARRYB[15][45] ), .S(\SUMB[15][45] ) );
  FA1A S4_51 ( .A(\ab[29][51] ), .B(\CARRYB[28][51] ), .CI(\SUMB[28][52] ), 
        .CO(\CARRYB[29][51] ), .S(\SUMB[29][51] ) );
  FA1A S4_48 ( .A(\ab[29][48] ), .B(\CARRYB[28][48] ), .CI(\SUMB[28][49] ), 
        .CO(\CARRYB[29][48] ), .S(\SUMB[29][48] ) );
  FA1A S3_14_94 ( .A(\ab[14][94] ), .B(\CARRYB[13][94] ), .CI(\ab[13][95] ), 
        .CO(\CARRYB[14][94] ), .S(\SUMB[14][94] ) );
  FA1A S3_13_94 ( .A(\ab[13][94] ), .B(\CARRYB[12][94] ), .CI(\ab[12][95] ), 
        .CO(\CARRYB[13][94] ), .S(\SUMB[13][94] ) );
  FA1A S3_12_94 ( .A(\ab[12][94] ), .B(\CARRYB[11][94] ), .CI(\ab[11][95] ), 
        .CO(\CARRYB[12][94] ), .S(\SUMB[12][94] ) );
  FA1A S3_11_94 ( .A(\ab[11][94] ), .B(\CARRYB[10][94] ), .CI(\ab[10][95] ), 
        .CO(\CARRYB[11][94] ), .S(\SUMB[11][94] ) );
  FA1A S3_10_94 ( .A(\ab[10][94] ), .B(\CARRYB[9][94] ), .CI(\ab[9][95] ), 
        .CO(\CARRYB[10][94] ), .S(\SUMB[10][94] ) );
  FA1A S3_9_94 ( .A(\ab[9][94] ), .B(\CARRYB[8][94] ), .CI(\ab[8][95] ), .CO(
        \CARRYB[9][94] ), .S(\SUMB[9][94] ) );
  FA1A S3_8_94 ( .A(\ab[8][94] ), .B(\CARRYB[7][94] ), .CI(\ab[7][95] ), .CO(
        \CARRYB[8][94] ), .S(\SUMB[8][94] ) );
  FA1A S3_7_94 ( .A(\ab[7][94] ), .B(\CARRYB[6][94] ), .CI(\ab[6][95] ), .CO(
        \CARRYB[7][94] ), .S(\SUMB[7][94] ) );
  FA1A S3_6_94 ( .A(\ab[6][94] ), .B(\CARRYB[5][94] ), .CI(\ab[5][95] ), .CO(
        \CARRYB[6][94] ), .S(\SUMB[6][94] ) );
  FA1A S3_5_94 ( .A(\ab[5][94] ), .B(\CARRYB[4][94] ), .CI(\ab[4][95] ), .CO(
        \CARRYB[5][94] ), .S(\SUMB[5][94] ) );
  FA1A S3_4_94 ( .A(\ab[4][94] ), .B(\CARRYB[3][94] ), .CI(\ab[3][95] ), .CO(
        \CARRYB[4][94] ), .S(\SUMB[4][94] ) );
  FA1A S3_3_94 ( .A(\ab[3][94] ), .B(\CARRYB[2][94] ), .CI(\ab[2][95] ), .CO(
        \CARRYB[3][94] ), .S(\SUMB[3][94] ) );
  FA1A S3_2_94 ( .A(\ab[2][94] ), .B(\CARRYB[1][94] ), .CI(\ab[1][95] ), .CO(
        \CARRYB[2][94] ), .S(\SUMB[2][94] ) );
  FA1A S2_14_93 ( .A(\ab[14][93] ), .B(\CARRYB[13][93] ), .CI(\SUMB[13][94] ), 
        .CO(\CARRYB[14][93] ), .S(\SUMB[14][93] ) );
  FA1A S2_13_93 ( .A(\ab[13][93] ), .B(\CARRYB[12][93] ), .CI(\SUMB[12][94] ), 
        .CO(\CARRYB[13][93] ), .S(\SUMB[13][93] ) );
  FA1A S2_12_93 ( .A(\ab[12][93] ), .B(\CARRYB[11][93] ), .CI(\SUMB[11][94] ), 
        .CO(\CARRYB[12][93] ), .S(\SUMB[12][93] ) );
  FA1A S2_11_93 ( .A(\ab[11][93] ), .B(\CARRYB[10][93] ), .CI(\SUMB[10][94] ), 
        .CO(\CARRYB[11][93] ), .S(\SUMB[11][93] ) );
  FA1A S2_10_93 ( .A(\ab[10][93] ), .B(\CARRYB[9][93] ), .CI(\SUMB[9][94] ), 
        .CO(\CARRYB[10][93] ), .S(\SUMB[10][93] ) );
  FA1A S2_9_93 ( .A(\ab[9][93] ), .B(\CARRYB[8][93] ), .CI(\SUMB[8][94] ), 
        .CO(\CARRYB[9][93] ), .S(\SUMB[9][93] ) );
  FA1A S2_8_93 ( .A(\ab[8][93] ), .B(\CARRYB[7][93] ), .CI(\SUMB[7][94] ), 
        .CO(\CARRYB[8][93] ), .S(\SUMB[8][93] ) );
  FA1A S2_7_93 ( .A(\ab[7][93] ), .B(\CARRYB[6][93] ), .CI(\SUMB[6][94] ), 
        .CO(\CARRYB[7][93] ), .S(\SUMB[7][93] ) );
  FA1A S2_6_93 ( .A(\ab[6][93] ), .B(\CARRYB[5][93] ), .CI(\SUMB[5][94] ), 
        .CO(\CARRYB[6][93] ), .S(\SUMB[6][93] ) );
  FA1A S2_5_93 ( .A(\ab[5][93] ), .B(\CARRYB[4][93] ), .CI(\SUMB[4][94] ), 
        .CO(\CARRYB[5][93] ), .S(\SUMB[5][93] ) );
  FA1A S2_4_93 ( .A(\ab[4][93] ), .B(\CARRYB[3][93] ), .CI(\SUMB[3][94] ), 
        .CO(\CARRYB[4][93] ), .S(\SUMB[4][93] ) );
  FA1A S2_3_93 ( .A(\ab[3][93] ), .B(\CARRYB[2][93] ), .CI(\SUMB[2][94] ), 
        .CO(\CARRYB[3][93] ), .S(\SUMB[3][93] ) );
  FA1A S2_2_93 ( .A(\ab[2][93] ), .B(\CARRYB[1][93] ), .CI(\SUMB[1][94] ), 
        .CO(\CARRYB[2][93] ), .S(\SUMB[2][93] ) );
  FA1A S2_14_92 ( .A(\ab[14][92] ), .B(\CARRYB[13][92] ), .CI(\SUMB[13][93] ), 
        .CO(\CARRYB[14][92] ), .S(\SUMB[14][92] ) );
  FA1A S2_13_92 ( .A(\ab[13][92] ), .B(\CARRYB[12][92] ), .CI(\SUMB[12][93] ), 
        .CO(\CARRYB[13][92] ), .S(\SUMB[13][92] ) );
  FA1A S2_12_92 ( .A(\ab[12][92] ), .B(\CARRYB[11][92] ), .CI(\SUMB[11][93] ), 
        .CO(\CARRYB[12][92] ), .S(\SUMB[12][92] ) );
  FA1A S2_11_92 ( .A(\ab[11][92] ), .B(\CARRYB[10][92] ), .CI(\SUMB[10][93] ), 
        .CO(\CARRYB[11][92] ), .S(\SUMB[11][92] ) );
  FA1A S2_10_92 ( .A(\ab[10][92] ), .B(\CARRYB[9][92] ), .CI(\SUMB[9][93] ), 
        .CO(\CARRYB[10][92] ), .S(\SUMB[10][92] ) );
  FA1A S2_9_92 ( .A(\ab[9][92] ), .B(\CARRYB[8][92] ), .CI(\SUMB[8][93] ), 
        .CO(\CARRYB[9][92] ), .S(\SUMB[9][92] ) );
  FA1A S2_8_92 ( .A(\ab[8][92] ), .B(\CARRYB[7][92] ), .CI(\SUMB[7][93] ), 
        .CO(\CARRYB[8][92] ), .S(\SUMB[8][92] ) );
  FA1A S2_7_92 ( .A(\ab[7][92] ), .B(\CARRYB[6][92] ), .CI(\SUMB[6][93] ), 
        .CO(\CARRYB[7][92] ), .S(\SUMB[7][92] ) );
  FA1A S2_6_92 ( .A(\ab[6][92] ), .B(\CARRYB[5][92] ), .CI(\SUMB[5][93] ), 
        .CO(\CARRYB[6][92] ), .S(\SUMB[6][92] ) );
  FA1A S2_5_92 ( .A(\ab[5][92] ), .B(\CARRYB[4][92] ), .CI(\SUMB[4][93] ), 
        .CO(\CARRYB[5][92] ), .S(\SUMB[5][92] ) );
  FA1A S2_4_92 ( .A(\ab[4][92] ), .B(\CARRYB[3][92] ), .CI(\SUMB[3][93] ), 
        .CO(\CARRYB[4][92] ), .S(\SUMB[4][92] ) );
  FA1A S2_3_92 ( .A(\ab[3][92] ), .B(\CARRYB[2][92] ), .CI(\SUMB[2][93] ), 
        .CO(\CARRYB[3][92] ), .S(\SUMB[3][92] ) );
  FA1A S2_2_92 ( .A(\ab[2][92] ), .B(\CARRYB[1][92] ), .CI(\SUMB[1][93] ), 
        .CO(\CARRYB[2][92] ), .S(\SUMB[2][92] ) );
  FA1A S2_14_91 ( .A(\ab[14][91] ), .B(\CARRYB[13][91] ), .CI(\SUMB[13][92] ), 
        .CO(\CARRYB[14][91] ), .S(\SUMB[14][91] ) );
  FA1A S2_13_91 ( .A(\ab[13][91] ), .B(\CARRYB[12][91] ), .CI(\SUMB[12][92] ), 
        .CO(\CARRYB[13][91] ), .S(\SUMB[13][91] ) );
  FA1A S2_12_91 ( .A(\ab[12][91] ), .B(\CARRYB[11][91] ), .CI(\SUMB[11][92] ), 
        .CO(\CARRYB[12][91] ), .S(\SUMB[12][91] ) );
  FA1A S2_11_91 ( .A(\ab[11][91] ), .B(\CARRYB[10][91] ), .CI(\SUMB[10][92] ), 
        .CO(\CARRYB[11][91] ), .S(\SUMB[11][91] ) );
  FA1A S2_10_91 ( .A(\ab[10][91] ), .B(\CARRYB[9][91] ), .CI(\SUMB[9][92] ), 
        .CO(\CARRYB[10][91] ), .S(\SUMB[10][91] ) );
  FA1A S2_9_91 ( .A(\ab[9][91] ), .B(\CARRYB[8][91] ), .CI(\SUMB[8][92] ), 
        .CO(\CARRYB[9][91] ), .S(\SUMB[9][91] ) );
  FA1A S2_8_91 ( .A(\ab[8][91] ), .B(\CARRYB[7][91] ), .CI(\SUMB[7][92] ), 
        .CO(\CARRYB[8][91] ), .S(\SUMB[8][91] ) );
  FA1A S2_7_91 ( .A(\ab[7][91] ), .B(\CARRYB[6][91] ), .CI(\SUMB[6][92] ), 
        .CO(\CARRYB[7][91] ), .S(\SUMB[7][91] ) );
  FA1A S2_6_91 ( .A(\ab[6][91] ), .B(\CARRYB[5][91] ), .CI(\SUMB[5][92] ), 
        .CO(\CARRYB[6][91] ), .S(\SUMB[6][91] ) );
  FA1A S2_5_91 ( .A(\ab[5][91] ), .B(\CARRYB[4][91] ), .CI(\SUMB[4][92] ), 
        .CO(\CARRYB[5][91] ), .S(\SUMB[5][91] ) );
  FA1A S2_4_91 ( .A(\ab[4][91] ), .B(\CARRYB[3][91] ), .CI(\SUMB[3][92] ), 
        .CO(\CARRYB[4][91] ), .S(\SUMB[4][91] ) );
  FA1A S2_3_91 ( .A(\ab[3][91] ), .B(\CARRYB[2][91] ), .CI(\SUMB[2][92] ), 
        .CO(\CARRYB[3][91] ), .S(\SUMB[3][91] ) );
  FA1A S2_2_91 ( .A(\ab[2][91] ), .B(\CARRYB[1][91] ), .CI(\SUMB[1][92] ), 
        .CO(\CARRYB[2][91] ), .S(\SUMB[2][91] ) );
  FA1A S2_14_90 ( .A(\ab[14][90] ), .B(\CARRYB[13][90] ), .CI(\SUMB[13][91] ), 
        .CO(\CARRYB[14][90] ), .S(\SUMB[14][90] ) );
  FA1A S2_13_90 ( .A(\ab[13][90] ), .B(\CARRYB[12][90] ), .CI(\SUMB[12][91] ), 
        .CO(\CARRYB[13][90] ), .S(\SUMB[13][90] ) );
  FA1A S2_12_90 ( .A(\ab[12][90] ), .B(\CARRYB[11][90] ), .CI(\SUMB[11][91] ), 
        .CO(\CARRYB[12][90] ), .S(\SUMB[12][90] ) );
  FA1A S2_11_90 ( .A(\ab[11][90] ), .B(\CARRYB[10][90] ), .CI(\SUMB[10][91] ), 
        .CO(\CARRYB[11][90] ), .S(\SUMB[11][90] ) );
  FA1A S2_10_90 ( .A(\ab[10][90] ), .B(\CARRYB[9][90] ), .CI(\SUMB[9][91] ), 
        .CO(\CARRYB[10][90] ), .S(\SUMB[10][90] ) );
  FA1A S2_9_90 ( .A(\ab[9][90] ), .B(\CARRYB[8][90] ), .CI(\SUMB[8][91] ), 
        .CO(\CARRYB[9][90] ), .S(\SUMB[9][90] ) );
  FA1A S2_8_90 ( .A(\ab[8][90] ), .B(\CARRYB[7][90] ), .CI(\SUMB[7][91] ), 
        .CO(\CARRYB[8][90] ), .S(\SUMB[8][90] ) );
  FA1A S2_7_90 ( .A(\ab[7][90] ), .B(\CARRYB[6][90] ), .CI(\SUMB[6][91] ), 
        .CO(\CARRYB[7][90] ), .S(\SUMB[7][90] ) );
  FA1A S2_6_90 ( .A(\ab[6][90] ), .B(\CARRYB[5][90] ), .CI(\SUMB[5][91] ), 
        .CO(\CARRYB[6][90] ), .S(\SUMB[6][90] ) );
  FA1A S2_5_90 ( .A(\ab[5][90] ), .B(\CARRYB[4][90] ), .CI(\SUMB[4][91] ), 
        .CO(\CARRYB[5][90] ), .S(\SUMB[5][90] ) );
  FA1A S2_4_90 ( .A(\ab[4][90] ), .B(\CARRYB[3][90] ), .CI(\SUMB[3][91] ), 
        .CO(\CARRYB[4][90] ), .S(\SUMB[4][90] ) );
  FA1A S2_3_90 ( .A(\ab[3][90] ), .B(\CARRYB[2][90] ), .CI(\SUMB[2][91] ), 
        .CO(\CARRYB[3][90] ), .S(\SUMB[3][90] ) );
  FA1A S2_2_90 ( .A(\ab[2][90] ), .B(\CARRYB[1][90] ), .CI(\SUMB[1][91] ), 
        .CO(\CARRYB[2][90] ), .S(\SUMB[2][90] ) );
  FA1A S2_14_89 ( .A(\ab[14][89] ), .B(\CARRYB[13][89] ), .CI(\SUMB[13][90] ), 
        .CO(\CARRYB[14][89] ), .S(\SUMB[14][89] ) );
  FA1A S2_13_89 ( .A(\ab[13][89] ), .B(\CARRYB[12][89] ), .CI(\SUMB[12][90] ), 
        .CO(\CARRYB[13][89] ), .S(\SUMB[13][89] ) );
  FA1A S2_12_89 ( .A(\ab[12][89] ), .B(\CARRYB[11][89] ), .CI(\SUMB[11][90] ), 
        .CO(\CARRYB[12][89] ), .S(\SUMB[12][89] ) );
  FA1A S2_11_89 ( .A(\ab[11][89] ), .B(\CARRYB[10][89] ), .CI(\SUMB[10][90] ), 
        .CO(\CARRYB[11][89] ), .S(\SUMB[11][89] ) );
  FA1A S2_10_89 ( .A(\ab[10][89] ), .B(\CARRYB[9][89] ), .CI(\SUMB[9][90] ), 
        .CO(\CARRYB[10][89] ), .S(\SUMB[10][89] ) );
  FA1A S2_9_89 ( .A(\ab[9][89] ), .B(\CARRYB[8][89] ), .CI(\SUMB[8][90] ), 
        .CO(\CARRYB[9][89] ), .S(\SUMB[9][89] ) );
  FA1A S2_8_89 ( .A(\ab[8][89] ), .B(\CARRYB[7][89] ), .CI(\SUMB[7][90] ), 
        .CO(\CARRYB[8][89] ), .S(\SUMB[8][89] ) );
  FA1A S2_7_89 ( .A(\ab[7][89] ), .B(\CARRYB[6][89] ), .CI(\SUMB[6][90] ), 
        .CO(\CARRYB[7][89] ), .S(\SUMB[7][89] ) );
  FA1A S2_6_89 ( .A(\ab[6][89] ), .B(\CARRYB[5][89] ), .CI(\SUMB[5][90] ), 
        .CO(\CARRYB[6][89] ), .S(\SUMB[6][89] ) );
  FA1A S2_5_89 ( .A(\ab[5][89] ), .B(\CARRYB[4][89] ), .CI(\SUMB[4][90] ), 
        .CO(\CARRYB[5][89] ), .S(\SUMB[5][89] ) );
  FA1A S2_4_89 ( .A(\ab[4][89] ), .B(\CARRYB[3][89] ), .CI(\SUMB[3][90] ), 
        .CO(\CARRYB[4][89] ), .S(\SUMB[4][89] ) );
  FA1A S2_3_89 ( .A(\ab[3][89] ), .B(\CARRYB[2][89] ), .CI(\SUMB[2][90] ), 
        .CO(\CARRYB[3][89] ), .S(\SUMB[3][89] ) );
  FA1A S2_2_89 ( .A(\ab[2][89] ), .B(\CARRYB[1][89] ), .CI(\SUMB[1][90] ), 
        .CO(\CARRYB[2][89] ), .S(\SUMB[2][89] ) );
  FA1A S2_14_88 ( .A(\ab[14][88] ), .B(\CARRYB[13][88] ), .CI(\SUMB[13][89] ), 
        .CO(\CARRYB[14][88] ), .S(\SUMB[14][88] ) );
  FA1A S2_13_88 ( .A(\ab[13][88] ), .B(\CARRYB[12][88] ), .CI(\SUMB[12][89] ), 
        .CO(\CARRYB[13][88] ), .S(\SUMB[13][88] ) );
  FA1A S2_12_88 ( .A(\ab[12][88] ), .B(\CARRYB[11][88] ), .CI(\SUMB[11][89] ), 
        .CO(\CARRYB[12][88] ), .S(\SUMB[12][88] ) );
  FA1A S2_11_88 ( .A(\ab[11][88] ), .B(\CARRYB[10][88] ), .CI(\SUMB[10][89] ), 
        .CO(\CARRYB[11][88] ), .S(\SUMB[11][88] ) );
  FA1A S2_10_88 ( .A(\ab[10][88] ), .B(\CARRYB[9][88] ), .CI(\SUMB[9][89] ), 
        .CO(\CARRYB[10][88] ), .S(\SUMB[10][88] ) );
  FA1A S2_9_88 ( .A(\ab[9][88] ), .B(\CARRYB[8][88] ), .CI(\SUMB[8][89] ), 
        .CO(\CARRYB[9][88] ), .S(\SUMB[9][88] ) );
  FA1A S2_8_88 ( .A(\ab[8][88] ), .B(\CARRYB[7][88] ), .CI(\SUMB[7][89] ), 
        .CO(\CARRYB[8][88] ), .S(\SUMB[8][88] ) );
  FA1A S2_7_88 ( .A(\ab[7][88] ), .B(\CARRYB[6][88] ), .CI(\SUMB[6][89] ), 
        .CO(\CARRYB[7][88] ), .S(\SUMB[7][88] ) );
  FA1A S2_6_88 ( .A(\ab[6][88] ), .B(\CARRYB[5][88] ), .CI(\SUMB[5][89] ), 
        .CO(\CARRYB[6][88] ), .S(\SUMB[6][88] ) );
  FA1A S2_5_88 ( .A(\ab[5][88] ), .B(\CARRYB[4][88] ), .CI(\SUMB[4][89] ), 
        .CO(\CARRYB[5][88] ), .S(\SUMB[5][88] ) );
  FA1A S2_4_88 ( .A(\ab[4][88] ), .B(\CARRYB[3][88] ), .CI(\SUMB[3][89] ), 
        .CO(\CARRYB[4][88] ), .S(\SUMB[4][88] ) );
  FA1A S2_3_88 ( .A(\ab[3][88] ), .B(\CARRYB[2][88] ), .CI(\SUMB[2][89] ), 
        .CO(\CARRYB[3][88] ), .S(\SUMB[3][88] ) );
  FA1A S2_2_88 ( .A(\ab[2][88] ), .B(\CARRYB[1][88] ), .CI(\SUMB[1][89] ), 
        .CO(\CARRYB[2][88] ), .S(\SUMB[2][88] ) );
  FA1A S2_14_87 ( .A(\ab[14][87] ), .B(\CARRYB[13][87] ), .CI(\SUMB[13][88] ), 
        .CO(\CARRYB[14][87] ), .S(\SUMB[14][87] ) );
  FA1A S2_13_87 ( .A(\ab[13][87] ), .B(\CARRYB[12][87] ), .CI(\SUMB[12][88] ), 
        .CO(\CARRYB[13][87] ), .S(\SUMB[13][87] ) );
  FA1A S2_12_87 ( .A(\ab[12][87] ), .B(\CARRYB[11][87] ), .CI(\SUMB[11][88] ), 
        .CO(\CARRYB[12][87] ), .S(\SUMB[12][87] ) );
  FA1A S2_11_87 ( .A(\ab[11][87] ), .B(\CARRYB[10][87] ), .CI(\SUMB[10][88] ), 
        .CO(\CARRYB[11][87] ), .S(\SUMB[11][87] ) );
  FA1A S2_10_87 ( .A(\ab[10][87] ), .B(\CARRYB[9][87] ), .CI(\SUMB[9][88] ), 
        .CO(\CARRYB[10][87] ), .S(\SUMB[10][87] ) );
  FA1A S2_9_87 ( .A(\ab[9][87] ), .B(\CARRYB[8][87] ), .CI(\SUMB[8][88] ), 
        .CO(\CARRYB[9][87] ), .S(\SUMB[9][87] ) );
  FA1A S2_8_87 ( .A(\ab[8][87] ), .B(\CARRYB[7][87] ), .CI(\SUMB[7][88] ), 
        .CO(\CARRYB[8][87] ), .S(\SUMB[8][87] ) );
  FA1A S2_7_87 ( .A(\ab[7][87] ), .B(\CARRYB[6][87] ), .CI(\SUMB[6][88] ), 
        .CO(\CARRYB[7][87] ), .S(\SUMB[7][87] ) );
  FA1A S2_6_87 ( .A(\ab[6][87] ), .B(\CARRYB[5][87] ), .CI(\SUMB[5][88] ), 
        .CO(\CARRYB[6][87] ), .S(\SUMB[6][87] ) );
  FA1A S2_5_87 ( .A(\ab[5][87] ), .B(\CARRYB[4][87] ), .CI(\SUMB[4][88] ), 
        .CO(\CARRYB[5][87] ), .S(\SUMB[5][87] ) );
  FA1A S2_4_87 ( .A(\ab[4][87] ), .B(\CARRYB[3][87] ), .CI(\SUMB[3][88] ), 
        .CO(\CARRYB[4][87] ), .S(\SUMB[4][87] ) );
  FA1A S2_3_87 ( .A(\ab[3][87] ), .B(\CARRYB[2][87] ), .CI(\SUMB[2][88] ), 
        .CO(\CARRYB[3][87] ), .S(\SUMB[3][87] ) );
  FA1A S2_2_87 ( .A(\ab[2][87] ), .B(\CARRYB[1][87] ), .CI(\SUMB[1][88] ), 
        .CO(\CARRYB[2][87] ), .S(\SUMB[2][87] ) );
  FA1A S2_14_86 ( .A(\ab[14][86] ), .B(\CARRYB[13][86] ), .CI(\SUMB[13][87] ), 
        .CO(\CARRYB[14][86] ), .S(\SUMB[14][86] ) );
  FA1A S2_13_86 ( .A(\ab[13][86] ), .B(\CARRYB[12][86] ), .CI(\SUMB[12][87] ), 
        .CO(\CARRYB[13][86] ), .S(\SUMB[13][86] ) );
  FA1A S2_12_86 ( .A(\ab[12][86] ), .B(\CARRYB[11][86] ), .CI(\SUMB[11][87] ), 
        .CO(\CARRYB[12][86] ), .S(\SUMB[12][86] ) );
  FA1A S2_11_86 ( .A(\ab[11][86] ), .B(\CARRYB[10][86] ), .CI(\SUMB[10][87] ), 
        .CO(\CARRYB[11][86] ), .S(\SUMB[11][86] ) );
  FA1A S2_10_86 ( .A(\ab[10][86] ), .B(\CARRYB[9][86] ), .CI(\SUMB[9][87] ), 
        .CO(\CARRYB[10][86] ), .S(\SUMB[10][86] ) );
  FA1A S2_9_86 ( .A(\ab[9][86] ), .B(\CARRYB[8][86] ), .CI(\SUMB[8][87] ), 
        .CO(\CARRYB[9][86] ), .S(\SUMB[9][86] ) );
  FA1A S2_8_86 ( .A(\ab[8][86] ), .B(\CARRYB[7][86] ), .CI(\SUMB[7][87] ), 
        .CO(\CARRYB[8][86] ), .S(\SUMB[8][86] ) );
  FA1A S2_7_86 ( .A(\ab[7][86] ), .B(\CARRYB[6][86] ), .CI(\SUMB[6][87] ), 
        .CO(\CARRYB[7][86] ), .S(\SUMB[7][86] ) );
  FA1A S2_6_86 ( .A(\ab[6][86] ), .B(\CARRYB[5][86] ), .CI(\SUMB[5][87] ), 
        .CO(\CARRYB[6][86] ), .S(\SUMB[6][86] ) );
  FA1A S2_5_86 ( .A(\ab[5][86] ), .B(\CARRYB[4][86] ), .CI(\SUMB[4][87] ), 
        .CO(\CARRYB[5][86] ), .S(\SUMB[5][86] ) );
  FA1A S2_4_86 ( .A(\ab[4][86] ), .B(\CARRYB[3][86] ), .CI(\SUMB[3][87] ), 
        .CO(\CARRYB[4][86] ), .S(\SUMB[4][86] ) );
  FA1A S2_3_86 ( .A(\ab[3][86] ), .B(\CARRYB[2][86] ), .CI(\SUMB[2][87] ), 
        .CO(\CARRYB[3][86] ), .S(\SUMB[3][86] ) );
  FA1A S2_2_86 ( .A(\ab[2][86] ), .B(\CARRYB[1][86] ), .CI(\SUMB[1][87] ), 
        .CO(\CARRYB[2][86] ), .S(\SUMB[2][86] ) );
  FA1A S2_14_85 ( .A(\ab[14][85] ), .B(\CARRYB[13][85] ), .CI(\SUMB[13][86] ), 
        .CO(\CARRYB[14][85] ), .S(\SUMB[14][85] ) );
  FA1A S2_13_85 ( .A(\ab[13][85] ), .B(\CARRYB[12][85] ), .CI(\SUMB[12][86] ), 
        .CO(\CARRYB[13][85] ), .S(\SUMB[13][85] ) );
  FA1A S2_12_85 ( .A(\ab[12][85] ), .B(\CARRYB[11][85] ), .CI(\SUMB[11][86] ), 
        .CO(\CARRYB[12][85] ), .S(\SUMB[12][85] ) );
  FA1A S2_11_85 ( .A(\ab[11][85] ), .B(\CARRYB[10][85] ), .CI(\SUMB[10][86] ), 
        .CO(\CARRYB[11][85] ), .S(\SUMB[11][85] ) );
  FA1A S2_10_85 ( .A(\ab[10][85] ), .B(\CARRYB[9][85] ), .CI(\SUMB[9][86] ), 
        .CO(\CARRYB[10][85] ), .S(\SUMB[10][85] ) );
  FA1A S2_9_85 ( .A(\ab[9][85] ), .B(\CARRYB[8][85] ), .CI(\SUMB[8][86] ), 
        .CO(\CARRYB[9][85] ), .S(\SUMB[9][85] ) );
  FA1A S2_8_85 ( .A(\ab[8][85] ), .B(\CARRYB[7][85] ), .CI(\SUMB[7][86] ), 
        .CO(\CARRYB[8][85] ), .S(\SUMB[8][85] ) );
  FA1A S2_7_85 ( .A(\ab[7][85] ), .B(\CARRYB[6][85] ), .CI(\SUMB[6][86] ), 
        .CO(\CARRYB[7][85] ), .S(\SUMB[7][85] ) );
  FA1A S2_6_85 ( .A(\ab[6][85] ), .B(\CARRYB[5][85] ), .CI(\SUMB[5][86] ), 
        .CO(\CARRYB[6][85] ), .S(\SUMB[6][85] ) );
  FA1A S2_5_85 ( .A(\ab[5][85] ), .B(\CARRYB[4][85] ), .CI(\SUMB[4][86] ), 
        .CO(\CARRYB[5][85] ), .S(\SUMB[5][85] ) );
  FA1A S2_4_85 ( .A(\ab[4][85] ), .B(\CARRYB[3][85] ), .CI(\SUMB[3][86] ), 
        .CO(\CARRYB[4][85] ), .S(\SUMB[4][85] ) );
  FA1A S2_3_85 ( .A(\ab[3][85] ), .B(\CARRYB[2][85] ), .CI(\SUMB[2][86] ), 
        .CO(\CARRYB[3][85] ), .S(\SUMB[3][85] ) );
  FA1A S2_2_85 ( .A(\ab[2][85] ), .B(\CARRYB[1][85] ), .CI(\SUMB[1][86] ), 
        .CO(\CARRYB[2][85] ), .S(\SUMB[2][85] ) );
  FA1A S2_14_81 ( .A(\ab[14][81] ), .B(\CARRYB[13][81] ), .CI(\SUMB[13][82] ), 
        .CO(\CARRYB[14][81] ), .S(\SUMB[14][81] ) );
  FA1A S2_13_81 ( .A(\ab[13][81] ), .B(\CARRYB[12][81] ), .CI(\SUMB[12][82] ), 
        .CO(\CARRYB[13][81] ), .S(\SUMB[13][81] ) );
  FA1A S2_12_81 ( .A(\ab[12][81] ), .B(\CARRYB[11][81] ), .CI(\SUMB[11][82] ), 
        .CO(\CARRYB[12][81] ), .S(\SUMB[12][81] ) );
  FA1A S2_11_81 ( .A(\ab[11][81] ), .B(\CARRYB[10][81] ), .CI(\SUMB[10][82] ), 
        .CO(\CARRYB[11][81] ), .S(\SUMB[11][81] ) );
  FA1A S2_10_81 ( .A(\ab[10][81] ), .B(\CARRYB[9][81] ), .CI(\SUMB[9][82] ), 
        .CO(\CARRYB[10][81] ), .S(\SUMB[10][81] ) );
  FA1A S2_9_81 ( .A(\ab[9][81] ), .B(\CARRYB[8][81] ), .CI(\SUMB[8][82] ), 
        .CO(\CARRYB[9][81] ), .S(\SUMB[9][81] ) );
  FA1A S2_8_81 ( .A(\ab[8][81] ), .B(\CARRYB[7][81] ), .CI(\SUMB[7][82] ), 
        .CO(\CARRYB[8][81] ), .S(\SUMB[8][81] ) );
  FA1A S2_7_81 ( .A(\ab[7][81] ), .B(\CARRYB[6][81] ), .CI(\SUMB[6][82] ), 
        .CO(\CARRYB[7][81] ), .S(\SUMB[7][81] ) );
  FA1A S2_6_81 ( .A(\ab[6][81] ), .B(\CARRYB[5][81] ), .CI(\SUMB[5][82] ), 
        .CO(\CARRYB[6][81] ), .S(\SUMB[6][81] ) );
  FA1A S2_5_81 ( .A(\ab[5][81] ), .B(\CARRYB[4][81] ), .CI(\SUMB[4][82] ), 
        .CO(\CARRYB[5][81] ), .S(\SUMB[5][81] ) );
  FA1A S2_4_81 ( .A(\ab[4][81] ), .B(\CARRYB[3][81] ), .CI(\SUMB[3][82] ), 
        .CO(\CARRYB[4][81] ), .S(\SUMB[4][81] ) );
  FA1A S2_3_81 ( .A(\ab[3][81] ), .B(\CARRYB[2][81] ), .CI(\SUMB[2][82] ), 
        .CO(\CARRYB[3][81] ), .S(\SUMB[3][81] ) );
  FA1A S2_2_81 ( .A(\ab[2][81] ), .B(\CARRYB[1][81] ), .CI(\SUMB[1][82] ), 
        .CO(\CARRYB[2][81] ), .S(\SUMB[2][81] ) );
  FA1A S2_14_84 ( .A(\ab[14][84] ), .B(\CARRYB[13][84] ), .CI(\SUMB[13][85] ), 
        .CO(\CARRYB[14][84] ), .S(\SUMB[14][84] ) );
  FA1A S2_14_83 ( .A(\ab[14][83] ), .B(\CARRYB[13][83] ), .CI(\SUMB[13][84] ), 
        .CO(\CARRYB[14][83] ), .S(\SUMB[14][83] ) );
  FA1A S2_13_84 ( .A(\ab[13][84] ), .B(\CARRYB[12][84] ), .CI(\SUMB[12][85] ), 
        .CO(\CARRYB[13][84] ), .S(\SUMB[13][84] ) );
  FA1A S2_14_80 ( .A(\ab[14][80] ), .B(\CARRYB[13][80] ), .CI(\SUMB[13][81] ), 
        .CO(\CARRYB[14][80] ), .S(\SUMB[14][80] ) );
  FA1A S2_14_82 ( .A(\ab[14][82] ), .B(\CARRYB[13][82] ), .CI(\SUMB[13][83] ), 
        .CO(\CARRYB[14][82] ), .S(\SUMB[14][82] ) );
  FA1A S2_13_80 ( .A(\ab[13][80] ), .B(\CARRYB[12][80] ), .CI(\SUMB[12][81] ), 
        .CO(\CARRYB[13][80] ), .S(\SUMB[13][80] ) );
  FA1A S2_13_82 ( .A(\ab[13][82] ), .B(\CARRYB[12][82] ), .CI(\SUMB[12][83] ), 
        .CO(\CARRYB[13][82] ), .S(\SUMB[13][82] ) );
  FA1A S2_13_83 ( .A(\ab[13][83] ), .B(\CARRYB[12][83] ), .CI(\SUMB[12][84] ), 
        .CO(\CARRYB[13][83] ), .S(\SUMB[13][83] ) );
  FA1A S2_12_80 ( .A(\ab[12][80] ), .B(\CARRYB[11][80] ), .CI(\SUMB[11][81] ), 
        .CO(\CARRYB[12][80] ), .S(\SUMB[12][80] ) );
  FA1A S2_12_82 ( .A(\ab[12][82] ), .B(\CARRYB[11][82] ), .CI(\SUMB[11][83] ), 
        .CO(\CARRYB[12][82] ), .S(\SUMB[12][82] ) );
  FA1A S2_12_83 ( .A(\ab[12][83] ), .B(\CARRYB[11][83] ), .CI(\SUMB[11][84] ), 
        .CO(\CARRYB[12][83] ), .S(\SUMB[12][83] ) );
  FA1A S2_12_84 ( .A(\ab[12][84] ), .B(\CARRYB[11][84] ), .CI(\SUMB[11][85] ), 
        .CO(\CARRYB[12][84] ), .S(\SUMB[12][84] ) );
  FA1A S2_11_82 ( .A(\ab[11][82] ), .B(\CARRYB[10][82] ), .CI(\SUMB[10][83] ), 
        .CO(\CARRYB[11][82] ), .S(\SUMB[11][82] ) );
  FA1A S2_11_83 ( .A(\ab[11][83] ), .B(\CARRYB[10][83] ), .CI(\SUMB[10][84] ), 
        .CO(\CARRYB[11][83] ), .S(\SUMB[11][83] ) );
  FA1A S2_11_84 ( .A(\ab[11][84] ), .B(\CARRYB[10][84] ), .CI(\SUMB[10][85] ), 
        .CO(\CARRYB[11][84] ), .S(\SUMB[11][84] ) );
  FA1A S2_10_82 ( .A(\ab[10][82] ), .B(\CARRYB[9][82] ), .CI(\SUMB[9][83] ), 
        .CO(\CARRYB[10][82] ), .S(\SUMB[10][82] ) );
  FA1A S2_10_83 ( .A(\ab[10][83] ), .B(\CARRYB[9][83] ), .CI(\SUMB[9][84] ), 
        .CO(\CARRYB[10][83] ), .S(\SUMB[10][83] ) );
  FA1A S2_10_84 ( .A(\ab[10][84] ), .B(\CARRYB[9][84] ), .CI(\SUMB[9][85] ), 
        .CO(\CARRYB[10][84] ), .S(\SUMB[10][84] ) );
  FA1A S2_9_83 ( .A(\ab[9][83] ), .B(\CARRYB[8][83] ), .CI(\SUMB[8][84] ), 
        .CO(\CARRYB[9][83] ), .S(\SUMB[9][83] ) );
  FA1A S2_9_84 ( .A(\ab[9][84] ), .B(\CARRYB[8][84] ), .CI(\SUMB[8][85] ), 
        .CO(\CARRYB[9][84] ), .S(\SUMB[9][84] ) );
  FA1A S2_11_80 ( .A(\ab[11][80] ), .B(\CARRYB[10][80] ), .CI(\SUMB[10][81] ), 
        .CO(\CARRYB[11][80] ), .S(\SUMB[11][80] ) );
  FA1A S2_8_84 ( .A(\ab[8][84] ), .B(\CARRYB[7][84] ), .CI(\SUMB[7][85] ), 
        .CO(\CARRYB[8][84] ), .S(\SUMB[8][84] ) );
  FA1A S2_10_80 ( .A(\ab[10][80] ), .B(\CARRYB[9][80] ), .CI(\SUMB[9][81] ), 
        .CO(\CARRYB[10][80] ), .S(\SUMB[10][80] ) );
  FA1A S2_9_80 ( .A(\ab[9][80] ), .B(\CARRYB[8][80] ), .CI(\SUMB[8][81] ), 
        .CO(\CARRYB[9][80] ), .S(\SUMB[9][80] ) );
  FA1A S2_9_82 ( .A(\ab[9][82] ), .B(\CARRYB[8][82] ), .CI(\SUMB[8][83] ), 
        .CO(\CARRYB[9][82] ), .S(\SUMB[9][82] ) );
  FA1A S2_8_80 ( .A(\ab[8][80] ), .B(\CARRYB[7][80] ), .CI(\SUMB[7][81] ), 
        .CO(\CARRYB[8][80] ), .S(\SUMB[8][80] ) );
  FA1A S2_8_82 ( .A(\ab[8][82] ), .B(\CARRYB[7][82] ), .CI(\SUMB[7][83] ), 
        .CO(\CARRYB[8][82] ), .S(\SUMB[8][82] ) );
  FA1A S2_8_83 ( .A(\ab[8][83] ), .B(\CARRYB[7][83] ), .CI(\SUMB[7][84] ), 
        .CO(\CARRYB[8][83] ), .S(\SUMB[8][83] ) );
  FA1A S2_7_82 ( .A(\ab[7][82] ), .B(\CARRYB[6][82] ), .CI(\SUMB[6][83] ), 
        .CO(\CARRYB[7][82] ), .S(\SUMB[7][82] ) );
  FA1A S2_7_80 ( .A(\ab[7][80] ), .B(\CARRYB[6][80] ), .CI(\SUMB[6][81] ), 
        .CO(\CARRYB[7][80] ), .S(\SUMB[7][80] ) );
  FA1A S2_7_83 ( .A(\ab[7][83] ), .B(\CARRYB[6][83] ), .CI(\SUMB[6][84] ), 
        .CO(\CARRYB[7][83] ), .S(\SUMB[7][83] ) );
  FA1A S2_7_84 ( .A(\ab[7][84] ), .B(\CARRYB[6][84] ), .CI(\SUMB[6][85] ), 
        .CO(\CARRYB[7][84] ), .S(\SUMB[7][84] ) );
  FA1A S2_6_83 ( .A(\ab[6][83] ), .B(\CARRYB[5][83] ), .CI(\SUMB[5][84] ), 
        .CO(\CARRYB[6][83] ), .S(\SUMB[6][83] ) );
  FA1A S2_6_82 ( .A(\ab[6][82] ), .B(\CARRYB[5][82] ), .CI(\SUMB[5][83] ), 
        .CO(\CARRYB[6][82] ), .S(\SUMB[6][82] ) );
  FA1A S2_6_80 ( .A(\ab[6][80] ), .B(\CARRYB[5][80] ), .CI(\SUMB[5][81] ), 
        .CO(\CARRYB[6][80] ), .S(\SUMB[6][80] ) );
  FA1A S2_6_84 ( .A(\ab[6][84] ), .B(\CARRYB[5][84] ), .CI(\SUMB[5][85] ), 
        .CO(\CARRYB[6][84] ), .S(\SUMB[6][84] ) );
  FA1A S2_5_84 ( .A(\ab[5][84] ), .B(\CARRYB[4][84] ), .CI(\SUMB[4][85] ), 
        .CO(\CARRYB[5][84] ), .S(\SUMB[5][84] ) );
  FA1A S2_5_83 ( .A(\ab[5][83] ), .B(\CARRYB[4][83] ), .CI(\SUMB[4][84] ), 
        .CO(\CARRYB[5][83] ), .S(\SUMB[5][83] ) );
  FA1A S2_5_82 ( .A(\ab[5][82] ), .B(\CARRYB[4][82] ), .CI(\SUMB[4][83] ), 
        .CO(\CARRYB[5][82] ), .S(\SUMB[5][82] ) );
  FA1A S2_5_80 ( .A(\ab[5][80] ), .B(\CARRYB[4][80] ), .CI(\SUMB[4][81] ), 
        .CO(\CARRYB[5][80] ), .S(\SUMB[5][80] ) );
  FA1A S2_4_84 ( .A(\ab[4][84] ), .B(\CARRYB[3][84] ), .CI(\SUMB[3][85] ), 
        .CO(\CARRYB[4][84] ), .S(\SUMB[4][84] ) );
  FA1A S2_4_83 ( .A(\ab[4][83] ), .B(\CARRYB[3][83] ), .CI(\SUMB[3][84] ), 
        .CO(\CARRYB[4][83] ), .S(\SUMB[4][83] ) );
  FA1A S2_4_82 ( .A(\ab[4][82] ), .B(\CARRYB[3][82] ), .CI(\SUMB[3][83] ), 
        .CO(\CARRYB[4][82] ), .S(\SUMB[4][82] ) );
  FA1A S2_4_80 ( .A(\ab[4][80] ), .B(\CARRYB[3][80] ), .CI(\SUMB[3][81] ), 
        .CO(\CARRYB[4][80] ), .S(\SUMB[4][80] ) );
  FA1A S2_3_84 ( .A(\ab[3][84] ), .B(\CARRYB[2][84] ), .CI(\SUMB[2][85] ), 
        .CO(\CARRYB[3][84] ), .S(\SUMB[3][84] ) );
  FA1A S2_3_83 ( .A(\ab[3][83] ), .B(\CARRYB[2][83] ), .CI(\SUMB[2][84] ), 
        .CO(\CARRYB[3][83] ), .S(\SUMB[3][83] ) );
  FA1A S2_3_82 ( .A(\ab[3][82] ), .B(\CARRYB[2][82] ), .CI(\SUMB[2][83] ), 
        .CO(\CARRYB[3][82] ), .S(\SUMB[3][82] ) );
  FA1A S2_3_80 ( .A(\ab[3][80] ), .B(\CARRYB[2][80] ), .CI(\SUMB[2][81] ), 
        .CO(\CARRYB[3][80] ), .S(\SUMB[3][80] ) );
  FA1A S2_2_84 ( .A(\ab[2][84] ), .B(\CARRYB[1][84] ), .CI(\SUMB[1][85] ), 
        .CO(\CARRYB[2][84] ), .S(\SUMB[2][84] ) );
  FA1A S2_2_83 ( .A(\ab[2][83] ), .B(\CARRYB[1][83] ), .CI(\SUMB[1][84] ), 
        .CO(\CARRYB[2][83] ), .S(\SUMB[2][83] ) );
  FA1A S2_2_82 ( .A(\ab[2][82] ), .B(\CARRYB[1][82] ), .CI(\SUMB[1][83] ), 
        .CO(\CARRYB[2][82] ), .S(\SUMB[2][82] ) );
  FA1A S2_2_80 ( .A(\ab[2][80] ), .B(\CARRYB[1][80] ), .CI(\SUMB[1][81] ), 
        .CO(\CARRYB[2][80] ), .S(\SUMB[2][80] ) );
  FA1A S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FA1A S4_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), .CO(
        \CARRYB[29][0] ), .S(\SUMB[29][0] ) );
  FA1A S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FA1A S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FA1A S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(\A1[22] ) );
  FA1A S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FA1A S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA1A S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\A1[21] ) );
  FA1A S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA1A S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FA1A S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA1A S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA1A S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA1A S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_14_78 ( .A(\ab[14][78] ), .B(\CARRYB[13][78] ), .CI(\SUMB[13][79] ), 
        .CO(\CARRYB[14][78] ), .S(\SUMB[14][78] ) );
  FA1A S2_14_79 ( .A(\ab[14][79] ), .B(\CARRYB[13][79] ), .CI(\SUMB[13][80] ), 
        .CO(\CARRYB[14][79] ), .S(\SUMB[14][79] ) );
  FA1A S2_13_79 ( .A(\ab[13][79] ), .B(\CARRYB[12][79] ), .CI(\SUMB[12][80] ), 
        .CO(\CARRYB[13][79] ), .S(\SUMB[13][79] ) );
  FA1A S2_14_75 ( .A(\ab[14][75] ), .B(\CARRYB[13][75] ), .CI(\SUMB[13][76] ), 
        .CO(\CARRYB[14][75] ), .S(\SUMB[14][75] ) );
  FA1A S2_14_74 ( .A(\ab[14][74] ), .B(\CARRYB[13][74] ), .CI(\SUMB[13][75] ), 
        .CO(\CARRYB[14][74] ), .S(\SUMB[14][74] ) );
  FA1A S2_14_73 ( .A(\ab[14][73] ), .B(\CARRYB[13][73] ), .CI(\SUMB[13][74] ), 
        .CO(\CARRYB[14][73] ), .S(\SUMB[14][73] ) );
  FA1A S2_14_72 ( .A(\ab[14][72] ), .B(\CARRYB[13][72] ), .CI(\SUMB[13][73] ), 
        .CO(\CARRYB[14][72] ), .S(\SUMB[14][72] ) );
  FA1A S2_14_71 ( .A(\ab[14][71] ), .B(\CARRYB[13][71] ), .CI(\SUMB[13][72] ), 
        .CO(\CARRYB[14][71] ), .S(\SUMB[14][71] ) );
  FA1A S2_14_70 ( .A(\ab[14][70] ), .B(\CARRYB[13][70] ), .CI(\SUMB[13][71] ), 
        .CO(\CARRYB[14][70] ), .S(\SUMB[14][70] ) );
  FA1A S2_14_69 ( .A(\ab[14][69] ), .B(\CARRYB[13][69] ), .CI(\SUMB[13][70] ), 
        .CO(\CARRYB[14][69] ), .S(\SUMB[14][69] ) );
  FA1A S2_14_76 ( .A(\ab[14][76] ), .B(\CARRYB[13][76] ), .CI(\SUMB[13][77] ), 
        .CO(\CARRYB[14][76] ), .S(\SUMB[14][76] ) );
  FA1A S2_14_77 ( .A(\ab[14][77] ), .B(\CARRYB[13][77] ), .CI(\SUMB[13][78] ), 
        .CO(\CARRYB[14][77] ), .S(\SUMB[14][77] ) );
  FA1A S2_13_76 ( .A(\ab[13][76] ), .B(\CARRYB[12][76] ), .CI(\SUMB[12][77] ), 
        .CO(\CARRYB[13][76] ), .S(\SUMB[13][76] ) );
  FA1A S2_13_75 ( .A(\ab[13][75] ), .B(\CARRYB[12][75] ), .CI(\SUMB[12][76] ), 
        .CO(\CARRYB[13][75] ), .S(\SUMB[13][75] ) );
  FA1A S2_13_74 ( .A(\ab[13][74] ), .B(\CARRYB[12][74] ), .CI(\SUMB[12][75] ), 
        .CO(\CARRYB[13][74] ), .S(\SUMB[13][74] ) );
  FA1A S2_13_73 ( .A(\ab[13][73] ), .B(\CARRYB[12][73] ), .CI(\SUMB[12][74] ), 
        .CO(\CARRYB[13][73] ), .S(\SUMB[13][73] ) );
  FA1A S2_13_72 ( .A(\ab[13][72] ), .B(\CARRYB[12][72] ), .CI(\SUMB[12][73] ), 
        .CO(\CARRYB[13][72] ), .S(\SUMB[13][72] ) );
  FA1A S2_13_71 ( .A(\ab[13][71] ), .B(\CARRYB[12][71] ), .CI(\SUMB[12][72] ), 
        .CO(\CARRYB[13][71] ), .S(\SUMB[13][71] ) );
  FA1A S2_13_70 ( .A(\ab[13][70] ), .B(\CARRYB[12][70] ), .CI(\SUMB[12][71] ), 
        .CO(\CARRYB[13][70] ), .S(\SUMB[13][70] ) );
  FA1A S2_13_69 ( .A(\ab[13][69] ), .B(\CARRYB[12][69] ), .CI(\SUMB[12][70] ), 
        .CO(\CARRYB[13][69] ), .S(\SUMB[13][69] ) );
  FA1A S2_13_77 ( .A(\ab[13][77] ), .B(\CARRYB[12][77] ), .CI(\SUMB[12][78] ), 
        .CO(\CARRYB[13][77] ), .S(\SUMB[13][77] ) );
  FA1A S2_13_78 ( .A(\ab[13][78] ), .B(\CARRYB[12][78] ), .CI(\SUMB[12][79] ), 
        .CO(\CARRYB[13][78] ), .S(\SUMB[13][78] ) );
  FA1A S2_12_77 ( .A(\ab[12][77] ), .B(\CARRYB[11][77] ), .CI(\SUMB[11][78] ), 
        .CO(\CARRYB[12][77] ), .S(\SUMB[12][77] ) );
  FA1A S2_12_76 ( .A(\ab[12][76] ), .B(\CARRYB[11][76] ), .CI(\SUMB[11][77] ), 
        .CO(\CARRYB[12][76] ), .S(\SUMB[12][76] ) );
  FA1A S2_12_75 ( .A(\ab[12][75] ), .B(\CARRYB[11][75] ), .CI(\SUMB[11][76] ), 
        .CO(\CARRYB[12][75] ), .S(\SUMB[12][75] ) );
  FA1A S2_12_74 ( .A(\ab[12][74] ), .B(\CARRYB[11][74] ), .CI(\SUMB[11][75] ), 
        .CO(\CARRYB[12][74] ), .S(\SUMB[12][74] ) );
  FA1A S2_12_73 ( .A(\ab[12][73] ), .B(\CARRYB[11][73] ), .CI(\SUMB[11][74] ), 
        .CO(\CARRYB[12][73] ), .S(\SUMB[12][73] ) );
  FA1A S2_12_72 ( .A(\ab[12][72] ), .B(\CARRYB[11][72] ), .CI(\SUMB[11][73] ), 
        .CO(\CARRYB[12][72] ), .S(\SUMB[12][72] ) );
  FA1A S2_12_71 ( .A(\ab[12][71] ), .B(\CARRYB[11][71] ), .CI(\SUMB[11][72] ), 
        .CO(\CARRYB[12][71] ), .S(\SUMB[12][71] ) );
  FA1A S2_12_70 ( .A(\ab[12][70] ), .B(\CARRYB[11][70] ), .CI(\SUMB[11][71] ), 
        .CO(\CARRYB[12][70] ), .S(\SUMB[12][70] ) );
  FA1A S2_12_69 ( .A(\ab[12][69] ), .B(\CARRYB[11][69] ), .CI(\SUMB[11][70] ), 
        .CO(\CARRYB[12][69] ), .S(\SUMB[12][69] ) );
  FA1A S2_12_78 ( .A(\ab[12][78] ), .B(\CARRYB[11][78] ), .CI(\SUMB[11][79] ), 
        .CO(\CARRYB[12][78] ), .S(\SUMB[12][78] ) );
  FA1A S2_12_79 ( .A(\ab[12][79] ), .B(\CARRYB[11][79] ), .CI(\SUMB[11][80] ), 
        .CO(\CARRYB[12][79] ), .S(\SUMB[12][79] ) );
  FA1A S2_11_78 ( .A(\ab[11][78] ), .B(\CARRYB[10][78] ), .CI(\SUMB[10][79] ), 
        .CO(\CARRYB[11][78] ), .S(\SUMB[11][78] ) );
  FA1A S2_11_77 ( .A(\ab[11][77] ), .B(\CARRYB[10][77] ), .CI(\SUMB[10][78] ), 
        .CO(\CARRYB[11][77] ), .S(\SUMB[11][77] ) );
  FA1A S2_11_76 ( .A(\ab[11][76] ), .B(\CARRYB[10][76] ), .CI(\SUMB[10][77] ), 
        .CO(\CARRYB[11][76] ), .S(\SUMB[11][76] ) );
  FA1A S2_11_75 ( .A(\ab[11][75] ), .B(\CARRYB[10][75] ), .CI(\SUMB[10][76] ), 
        .CO(\CARRYB[11][75] ), .S(\SUMB[11][75] ) );
  FA1A S2_11_74 ( .A(\ab[11][74] ), .B(\CARRYB[10][74] ), .CI(\SUMB[10][75] ), 
        .CO(\CARRYB[11][74] ), .S(\SUMB[11][74] ) );
  FA1A S2_11_73 ( .A(\ab[11][73] ), .B(\CARRYB[10][73] ), .CI(\SUMB[10][74] ), 
        .CO(\CARRYB[11][73] ), .S(\SUMB[11][73] ) );
  FA1A S2_11_72 ( .A(\ab[11][72] ), .B(\CARRYB[10][72] ), .CI(\SUMB[10][73] ), 
        .CO(\CARRYB[11][72] ), .S(\SUMB[11][72] ) );
  FA1A S2_11_71 ( .A(\ab[11][71] ), .B(\CARRYB[10][71] ), .CI(\SUMB[10][72] ), 
        .CO(\CARRYB[11][71] ), .S(\SUMB[11][71] ) );
  FA1A S2_11_70 ( .A(\ab[11][70] ), .B(\CARRYB[10][70] ), .CI(\SUMB[10][71] ), 
        .CO(\CARRYB[11][70] ), .S(\SUMB[11][70] ) );
  FA1A S2_11_69 ( .A(\ab[11][69] ), .B(\CARRYB[10][69] ), .CI(\SUMB[10][70] ), 
        .CO(\CARRYB[11][69] ), .S(\SUMB[11][69] ) );
  FA1A S2_11_79 ( .A(\ab[11][79] ), .B(\CARRYB[10][79] ), .CI(\SUMB[10][80] ), 
        .CO(\CARRYB[11][79] ), .S(\SUMB[11][79] ) );
  FA1A S2_10_79 ( .A(\ab[10][79] ), .B(\CARRYB[9][79] ), .CI(\SUMB[9][80] ), 
        .CO(\CARRYB[10][79] ), .S(\SUMB[10][79] ) );
  FA1A S2_10_78 ( .A(\ab[10][78] ), .B(\CARRYB[9][78] ), .CI(\SUMB[9][79] ), 
        .CO(\CARRYB[10][78] ), .S(\SUMB[10][78] ) );
  FA1A S2_10_77 ( .A(\ab[10][77] ), .B(\CARRYB[9][77] ), .CI(\SUMB[9][78] ), 
        .CO(\CARRYB[10][77] ), .S(\SUMB[10][77] ) );
  FA1A S2_10_76 ( .A(\ab[10][76] ), .B(\CARRYB[9][76] ), .CI(\SUMB[9][77] ), 
        .CO(\CARRYB[10][76] ), .S(\SUMB[10][76] ) );
  FA1A S2_10_75 ( .A(\ab[10][75] ), .B(\CARRYB[9][75] ), .CI(\SUMB[9][76] ), 
        .CO(\CARRYB[10][75] ), .S(\SUMB[10][75] ) );
  FA1A S2_10_74 ( .A(\ab[10][74] ), .B(\CARRYB[9][74] ), .CI(\SUMB[9][75] ), 
        .CO(\CARRYB[10][74] ), .S(\SUMB[10][74] ) );
  FA1A S2_10_73 ( .A(\ab[10][73] ), .B(\CARRYB[9][73] ), .CI(\SUMB[9][74] ), 
        .CO(\CARRYB[10][73] ), .S(\SUMB[10][73] ) );
  FA1A S2_10_72 ( .A(\ab[10][72] ), .B(\CARRYB[9][72] ), .CI(\SUMB[9][73] ), 
        .CO(\CARRYB[10][72] ), .S(\SUMB[10][72] ) );
  FA1A S2_10_71 ( .A(\ab[10][71] ), .B(\CARRYB[9][71] ), .CI(\SUMB[9][72] ), 
        .CO(\CARRYB[10][71] ), .S(\SUMB[10][71] ) );
  FA1A S2_10_70 ( .A(\ab[10][70] ), .B(\CARRYB[9][70] ), .CI(\SUMB[9][71] ), 
        .CO(\CARRYB[10][70] ), .S(\SUMB[10][70] ) );
  FA1A S2_10_69 ( .A(\ab[10][69] ), .B(\CARRYB[9][69] ), .CI(\SUMB[9][70] ), 
        .CO(\CARRYB[10][69] ), .S(\SUMB[10][69] ) );
  FA1A S2_9_79 ( .A(\ab[9][79] ), .B(\CARRYB[8][79] ), .CI(\SUMB[8][80] ), 
        .CO(\CARRYB[9][79] ), .S(\SUMB[9][79] ) );
  FA1A S2_9_78 ( .A(\ab[9][78] ), .B(\CARRYB[8][78] ), .CI(\SUMB[8][79] ), 
        .CO(\CARRYB[9][78] ), .S(\SUMB[9][78] ) );
  FA1A S2_9_77 ( .A(\ab[9][77] ), .B(\CARRYB[8][77] ), .CI(\SUMB[8][78] ), 
        .CO(\CARRYB[9][77] ), .S(\SUMB[9][77] ) );
  FA1A S2_9_76 ( .A(\ab[9][76] ), .B(\CARRYB[8][76] ), .CI(\SUMB[8][77] ), 
        .CO(\CARRYB[9][76] ), .S(\SUMB[9][76] ) );
  FA1A S2_9_75 ( .A(\ab[9][75] ), .B(\CARRYB[8][75] ), .CI(\SUMB[8][76] ), 
        .CO(\CARRYB[9][75] ), .S(\SUMB[9][75] ) );
  FA1A S2_9_74 ( .A(\ab[9][74] ), .B(\CARRYB[8][74] ), .CI(\SUMB[8][75] ), 
        .CO(\CARRYB[9][74] ), .S(\SUMB[9][74] ) );
  FA1A S2_9_73 ( .A(\ab[9][73] ), .B(\CARRYB[8][73] ), .CI(\SUMB[8][74] ), 
        .CO(\CARRYB[9][73] ), .S(\SUMB[9][73] ) );
  FA1A S2_9_72 ( .A(\ab[9][72] ), .B(\CARRYB[8][72] ), .CI(\SUMB[8][73] ), 
        .CO(\CARRYB[9][72] ), .S(\SUMB[9][72] ) );
  FA1A S2_9_71 ( .A(\ab[9][71] ), .B(\CARRYB[8][71] ), .CI(\SUMB[8][72] ), 
        .CO(\CARRYB[9][71] ), .S(\SUMB[9][71] ) );
  FA1A S2_9_70 ( .A(\ab[9][70] ), .B(\CARRYB[8][70] ), .CI(\SUMB[8][71] ), 
        .CO(\CARRYB[9][70] ), .S(\SUMB[9][70] ) );
  FA1A S2_9_69 ( .A(\ab[9][69] ), .B(\CARRYB[8][69] ), .CI(\SUMB[8][70] ), 
        .CO(\CARRYB[9][69] ), .S(\SUMB[9][69] ) );
  FA1A S2_8_79 ( .A(\ab[8][79] ), .B(\CARRYB[7][79] ), .CI(\SUMB[7][80] ), 
        .CO(\CARRYB[8][79] ), .S(\SUMB[8][79] ) );
  FA1A S2_8_78 ( .A(\ab[8][78] ), .B(\CARRYB[7][78] ), .CI(\SUMB[7][79] ), 
        .CO(\CARRYB[8][78] ), .S(\SUMB[8][78] ) );
  FA1A S2_8_77 ( .A(\ab[8][77] ), .B(\CARRYB[7][77] ), .CI(\SUMB[7][78] ), 
        .CO(\CARRYB[8][77] ), .S(\SUMB[8][77] ) );
  FA1A S2_8_76 ( .A(\ab[8][76] ), .B(\CARRYB[7][76] ), .CI(\SUMB[7][77] ), 
        .CO(\CARRYB[8][76] ), .S(\SUMB[8][76] ) );
  FA1A S2_8_75 ( .A(\ab[8][75] ), .B(\CARRYB[7][75] ), .CI(\SUMB[7][76] ), 
        .CO(\CARRYB[8][75] ), .S(\SUMB[8][75] ) );
  FA1A S2_8_74 ( .A(\ab[8][74] ), .B(\CARRYB[7][74] ), .CI(\SUMB[7][75] ), 
        .CO(\CARRYB[8][74] ), .S(\SUMB[8][74] ) );
  FA1A S2_8_73 ( .A(\ab[8][73] ), .B(\CARRYB[7][73] ), .CI(\SUMB[7][74] ), 
        .CO(\CARRYB[8][73] ), .S(\SUMB[8][73] ) );
  FA1A S2_8_72 ( .A(\ab[8][72] ), .B(\CARRYB[7][72] ), .CI(\SUMB[7][73] ), 
        .CO(\CARRYB[8][72] ), .S(\SUMB[8][72] ) );
  FA1A S2_8_71 ( .A(\ab[8][71] ), .B(\CARRYB[7][71] ), .CI(\SUMB[7][72] ), 
        .CO(\CARRYB[8][71] ), .S(\SUMB[8][71] ) );
  FA1A S2_8_70 ( .A(\ab[8][70] ), .B(\CARRYB[7][70] ), .CI(\SUMB[7][71] ), 
        .CO(\CARRYB[8][70] ), .S(\SUMB[8][70] ) );
  FA1A S2_8_69 ( .A(\ab[8][69] ), .B(\CARRYB[7][69] ), .CI(\SUMB[7][70] ), 
        .CO(\CARRYB[8][69] ), .S(\SUMB[8][69] ) );
  FA1A S2_7_79 ( .A(\ab[7][79] ), .B(\CARRYB[6][79] ), .CI(\SUMB[6][80] ), 
        .CO(\CARRYB[7][79] ), .S(\SUMB[7][79] ) );
  FA1A S2_7_78 ( .A(\ab[7][78] ), .B(\CARRYB[6][78] ), .CI(\SUMB[6][79] ), 
        .CO(\CARRYB[7][78] ), .S(\SUMB[7][78] ) );
  FA1A S2_7_77 ( .A(\ab[7][77] ), .B(\CARRYB[6][77] ), .CI(\SUMB[6][78] ), 
        .CO(\CARRYB[7][77] ), .S(\SUMB[7][77] ) );
  FA1A S2_7_76 ( .A(\ab[7][76] ), .B(\CARRYB[6][76] ), .CI(\SUMB[6][77] ), 
        .CO(\CARRYB[7][76] ), .S(\SUMB[7][76] ) );
  FA1A S2_7_75 ( .A(\ab[7][75] ), .B(\CARRYB[6][75] ), .CI(\SUMB[6][76] ), 
        .CO(\CARRYB[7][75] ), .S(\SUMB[7][75] ) );
  FA1A S2_7_74 ( .A(\ab[7][74] ), .B(\CARRYB[6][74] ), .CI(\SUMB[6][75] ), 
        .CO(\CARRYB[7][74] ), .S(\SUMB[7][74] ) );
  FA1A S2_7_73 ( .A(\ab[7][73] ), .B(\CARRYB[6][73] ), .CI(\SUMB[6][74] ), 
        .CO(\CARRYB[7][73] ), .S(\SUMB[7][73] ) );
  FA1A S2_7_72 ( .A(\ab[7][72] ), .B(\CARRYB[6][72] ), .CI(\SUMB[6][73] ), 
        .CO(\CARRYB[7][72] ), .S(\SUMB[7][72] ) );
  FA1A S2_7_71 ( .A(\ab[7][71] ), .B(\CARRYB[6][71] ), .CI(\SUMB[6][72] ), 
        .CO(\CARRYB[7][71] ), .S(\SUMB[7][71] ) );
  FA1A S2_7_70 ( .A(\ab[7][70] ), .B(\CARRYB[6][70] ), .CI(\SUMB[6][71] ), 
        .CO(\CARRYB[7][70] ), .S(\SUMB[7][70] ) );
  FA1A S2_7_69 ( .A(\ab[7][69] ), .B(\CARRYB[6][69] ), .CI(\SUMB[6][70] ), 
        .CO(\CARRYB[7][69] ), .S(\SUMB[7][69] ) );
  FA1A S2_6_79 ( .A(\ab[6][79] ), .B(\CARRYB[5][79] ), .CI(\SUMB[5][80] ), 
        .CO(\CARRYB[6][79] ), .S(\SUMB[6][79] ) );
  FA1A S2_6_78 ( .A(\ab[6][78] ), .B(\CARRYB[5][78] ), .CI(\SUMB[5][79] ), 
        .CO(\CARRYB[6][78] ), .S(\SUMB[6][78] ) );
  FA1A S2_6_77 ( .A(\ab[6][77] ), .B(\CARRYB[5][77] ), .CI(\SUMB[5][78] ), 
        .CO(\CARRYB[6][77] ), .S(\SUMB[6][77] ) );
  FA1A S2_6_76 ( .A(\ab[6][76] ), .B(\CARRYB[5][76] ), .CI(\SUMB[5][77] ), 
        .CO(\CARRYB[6][76] ), .S(\SUMB[6][76] ) );
  FA1A S2_6_75 ( .A(\ab[6][75] ), .B(\CARRYB[5][75] ), .CI(\SUMB[5][76] ), 
        .CO(\CARRYB[6][75] ), .S(\SUMB[6][75] ) );
  FA1A S2_6_74 ( .A(\ab[6][74] ), .B(\CARRYB[5][74] ), .CI(\SUMB[5][75] ), 
        .CO(\CARRYB[6][74] ), .S(\SUMB[6][74] ) );
  FA1A S2_6_73 ( .A(\ab[6][73] ), .B(\CARRYB[5][73] ), .CI(\SUMB[5][74] ), 
        .CO(\CARRYB[6][73] ), .S(\SUMB[6][73] ) );
  FA1A S2_6_72 ( .A(\ab[6][72] ), .B(\CARRYB[5][72] ), .CI(\SUMB[5][73] ), 
        .CO(\CARRYB[6][72] ), .S(\SUMB[6][72] ) );
  FA1A S2_6_71 ( .A(\ab[6][71] ), .B(\CARRYB[5][71] ), .CI(\SUMB[5][72] ), 
        .CO(\CARRYB[6][71] ), .S(\SUMB[6][71] ) );
  FA1A S2_6_70 ( .A(\ab[6][70] ), .B(\CARRYB[5][70] ), .CI(\SUMB[5][71] ), 
        .CO(\CARRYB[6][70] ), .S(\SUMB[6][70] ) );
  FA1A S2_6_69 ( .A(\ab[6][69] ), .B(\CARRYB[5][69] ), .CI(\SUMB[5][70] ), 
        .CO(\CARRYB[6][69] ), .S(\SUMB[6][69] ) );
  FA1A S2_5_79 ( .A(\ab[5][79] ), .B(\CARRYB[4][79] ), .CI(\SUMB[4][80] ), 
        .CO(\CARRYB[5][79] ), .S(\SUMB[5][79] ) );
  FA1A S2_5_78 ( .A(\ab[5][78] ), .B(\CARRYB[4][78] ), .CI(\SUMB[4][79] ), 
        .CO(\CARRYB[5][78] ), .S(\SUMB[5][78] ) );
  FA1A S2_5_77 ( .A(\ab[5][77] ), .B(\CARRYB[4][77] ), .CI(\SUMB[4][78] ), 
        .CO(\CARRYB[5][77] ), .S(\SUMB[5][77] ) );
  FA1A S2_5_76 ( .A(\ab[5][76] ), .B(\CARRYB[4][76] ), .CI(\SUMB[4][77] ), 
        .CO(\CARRYB[5][76] ), .S(\SUMB[5][76] ) );
  FA1A S2_5_75 ( .A(\ab[5][75] ), .B(\CARRYB[4][75] ), .CI(\SUMB[4][76] ), 
        .CO(\CARRYB[5][75] ), .S(\SUMB[5][75] ) );
  FA1A S2_5_74 ( .A(\ab[5][74] ), .B(\CARRYB[4][74] ), .CI(\SUMB[4][75] ), 
        .CO(\CARRYB[5][74] ), .S(\SUMB[5][74] ) );
  FA1A S2_5_73 ( .A(\ab[5][73] ), .B(\CARRYB[4][73] ), .CI(\SUMB[4][74] ), 
        .CO(\CARRYB[5][73] ), .S(\SUMB[5][73] ) );
  FA1A S2_5_72 ( .A(\ab[5][72] ), .B(\CARRYB[4][72] ), .CI(\SUMB[4][73] ), 
        .CO(\CARRYB[5][72] ), .S(\SUMB[5][72] ) );
  FA1A S2_5_71 ( .A(\ab[5][71] ), .B(\CARRYB[4][71] ), .CI(\SUMB[4][72] ), 
        .CO(\CARRYB[5][71] ), .S(\SUMB[5][71] ) );
  FA1A S2_5_70 ( .A(\ab[5][70] ), .B(\CARRYB[4][70] ), .CI(\SUMB[4][71] ), 
        .CO(\CARRYB[5][70] ), .S(\SUMB[5][70] ) );
  FA1A S2_5_69 ( .A(\ab[5][69] ), .B(\CARRYB[4][69] ), .CI(\SUMB[4][70] ), 
        .CO(\CARRYB[5][69] ), .S(\SUMB[5][69] ) );
  FA1A S2_4_79 ( .A(\ab[4][79] ), .B(\CARRYB[3][79] ), .CI(\SUMB[3][80] ), 
        .CO(\CARRYB[4][79] ), .S(\SUMB[4][79] ) );
  FA1A S2_4_78 ( .A(\ab[4][78] ), .B(\CARRYB[3][78] ), .CI(\SUMB[3][79] ), 
        .CO(\CARRYB[4][78] ), .S(\SUMB[4][78] ) );
  FA1A S2_4_77 ( .A(\ab[4][77] ), .B(\CARRYB[3][77] ), .CI(\SUMB[3][78] ), 
        .CO(\CARRYB[4][77] ), .S(\SUMB[4][77] ) );
  FA1A S2_4_76 ( .A(\ab[4][76] ), .B(\CARRYB[3][76] ), .CI(\SUMB[3][77] ), 
        .CO(\CARRYB[4][76] ), .S(\SUMB[4][76] ) );
  FA1A S2_4_75 ( .A(\ab[4][75] ), .B(\CARRYB[3][75] ), .CI(\SUMB[3][76] ), 
        .CO(\CARRYB[4][75] ), .S(\SUMB[4][75] ) );
  FA1A S2_4_74 ( .A(\ab[4][74] ), .B(\CARRYB[3][74] ), .CI(\SUMB[3][75] ), 
        .CO(\CARRYB[4][74] ), .S(\SUMB[4][74] ) );
  FA1A S2_4_73 ( .A(\ab[4][73] ), .B(\CARRYB[3][73] ), .CI(\SUMB[3][74] ), 
        .CO(\CARRYB[4][73] ), .S(\SUMB[4][73] ) );
  FA1A S2_4_72 ( .A(\ab[4][72] ), .B(\CARRYB[3][72] ), .CI(\SUMB[3][73] ), 
        .CO(\CARRYB[4][72] ), .S(\SUMB[4][72] ) );
  FA1A S2_4_71 ( .A(\ab[4][71] ), .B(\CARRYB[3][71] ), .CI(\SUMB[3][72] ), 
        .CO(\CARRYB[4][71] ), .S(\SUMB[4][71] ) );
  FA1A S2_4_70 ( .A(\ab[4][70] ), .B(\CARRYB[3][70] ), .CI(\SUMB[3][71] ), 
        .CO(\CARRYB[4][70] ), .S(\SUMB[4][70] ) );
  FA1A S2_4_69 ( .A(\ab[4][69] ), .B(\CARRYB[3][69] ), .CI(\SUMB[3][70] ), 
        .CO(\CARRYB[4][69] ), .S(\SUMB[4][69] ) );
  FA1A S2_3_79 ( .A(\ab[3][79] ), .B(\CARRYB[2][79] ), .CI(\SUMB[2][80] ), 
        .CO(\CARRYB[3][79] ), .S(\SUMB[3][79] ) );
  FA1A S2_3_78 ( .A(\ab[3][78] ), .B(\CARRYB[2][78] ), .CI(\SUMB[2][79] ), 
        .CO(\CARRYB[3][78] ), .S(\SUMB[3][78] ) );
  FA1A S2_3_77 ( .A(\ab[3][77] ), .B(\CARRYB[2][77] ), .CI(\SUMB[2][78] ), 
        .CO(\CARRYB[3][77] ), .S(\SUMB[3][77] ) );
  FA1A S2_3_76 ( .A(\ab[3][76] ), .B(\CARRYB[2][76] ), .CI(\SUMB[2][77] ), 
        .CO(\CARRYB[3][76] ), .S(\SUMB[3][76] ) );
  FA1A S2_3_75 ( .A(\ab[3][75] ), .B(\CARRYB[2][75] ), .CI(\SUMB[2][76] ), 
        .CO(\CARRYB[3][75] ), .S(\SUMB[3][75] ) );
  FA1A S2_3_74 ( .A(\ab[3][74] ), .B(\CARRYB[2][74] ), .CI(\SUMB[2][75] ), 
        .CO(\CARRYB[3][74] ), .S(\SUMB[3][74] ) );
  FA1A S2_3_73 ( .A(\ab[3][73] ), .B(\CARRYB[2][73] ), .CI(\SUMB[2][74] ), 
        .CO(\CARRYB[3][73] ), .S(\SUMB[3][73] ) );
  FA1A S2_3_72 ( .A(\ab[3][72] ), .B(\CARRYB[2][72] ), .CI(\SUMB[2][73] ), 
        .CO(\CARRYB[3][72] ), .S(\SUMB[3][72] ) );
  FA1A S2_3_71 ( .A(\ab[3][71] ), .B(\CARRYB[2][71] ), .CI(\SUMB[2][72] ), 
        .CO(\CARRYB[3][71] ), .S(\SUMB[3][71] ) );
  FA1A S2_3_70 ( .A(\ab[3][70] ), .B(\CARRYB[2][70] ), .CI(\SUMB[2][71] ), 
        .CO(\CARRYB[3][70] ), .S(\SUMB[3][70] ) );
  FA1A S2_3_69 ( .A(\ab[3][69] ), .B(\CARRYB[2][69] ), .CI(\SUMB[2][70] ), 
        .CO(\CARRYB[3][69] ), .S(\SUMB[3][69] ) );
  FA1A S2_2_79 ( .A(\ab[2][79] ), .B(\CARRYB[1][79] ), .CI(\SUMB[1][80] ), 
        .CO(\CARRYB[2][79] ), .S(\SUMB[2][79] ) );
  FA1A S2_2_78 ( .A(\ab[2][78] ), .B(\CARRYB[1][78] ), .CI(\SUMB[1][79] ), 
        .CO(\CARRYB[2][78] ), .S(\SUMB[2][78] ) );
  FA1A S2_2_77 ( .A(\ab[2][77] ), .B(\CARRYB[1][77] ), .CI(\SUMB[1][78] ), 
        .CO(\CARRYB[2][77] ), .S(\SUMB[2][77] ) );
  FA1A S2_2_76 ( .A(\ab[2][76] ), .B(\CARRYB[1][76] ), .CI(\SUMB[1][77] ), 
        .CO(\CARRYB[2][76] ), .S(\SUMB[2][76] ) );
  FA1A S2_2_75 ( .A(\ab[2][75] ), .B(\CARRYB[1][75] ), .CI(\SUMB[1][76] ), 
        .CO(\CARRYB[2][75] ), .S(\SUMB[2][75] ) );
  FA1A S2_2_74 ( .A(\ab[2][74] ), .B(\CARRYB[1][74] ), .CI(\SUMB[1][75] ), 
        .CO(\CARRYB[2][74] ), .S(\SUMB[2][74] ) );
  FA1A S2_2_73 ( .A(\ab[2][73] ), .B(\CARRYB[1][73] ), .CI(\SUMB[1][74] ), 
        .CO(\CARRYB[2][73] ), .S(\SUMB[2][73] ) );
  FA1A S2_2_72 ( .A(\ab[2][72] ), .B(\CARRYB[1][72] ), .CI(\SUMB[1][73] ), 
        .CO(\CARRYB[2][72] ), .S(\SUMB[2][72] ) );
  FA1A S2_2_71 ( .A(\ab[2][71] ), .B(\CARRYB[1][71] ), .CI(\SUMB[1][72] ), 
        .CO(\CARRYB[2][71] ), .S(\SUMB[2][71] ) );
  FA1A S2_2_70 ( .A(\ab[2][70] ), .B(\CARRYB[1][70] ), .CI(\SUMB[1][71] ), 
        .CO(\CARRYB[2][70] ), .S(\SUMB[2][70] ) );
  FA1A S2_2_69 ( .A(\ab[2][69] ), .B(\CARRYB[1][69] ), .CI(\SUMB[1][70] ), 
        .CO(\CARRYB[2][69] ), .S(\SUMB[2][69] ) );
  FA1A S4_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), .CO(
        \CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA1A S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA1A S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA1A S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA1A S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA1A S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA1A S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA1A S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA1A S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1A S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1A S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA1A S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1A S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1A S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1A S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S4_30 ( .A(\ab[29][30] ), .B(\CARRYB[28][30] ), .CI(\SUMB[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FA1A S4_29 ( .A(\ab[29][29] ), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), 
        .CO(\CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_28_30 ( .A(\ab[28][30] ), .B(\CARRYB[27][30] ), .CI(\SUMB[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA1A S2_28_29 ( .A(\ab[28][29] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_27_30 ( .A(\ab[27][30] ), .B(\CARRYB[26][30] ), .CI(\SUMB[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_27_29 ( .A(\ab[27][29] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_26_29 ( .A(\ab[26][29] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA1A S2_26_30 ( .A(\ab[26][30] ), .B(\CARRYB[25][30] ), .CI(\SUMB[25][31] ), 
        .CO(\CARRYB[26][30] ), .S(\SUMB[26][30] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_25_30 ( .A(\ab[25][30] ), .B(\CARRYB[24][30] ), .CI(\SUMB[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_25_29 ( .A(\ab[25][29] ), .B(\CARRYB[24][29] ), .CI(\SUMB[24][30] ), 
        .CO(\CARRYB[25][29] ), .S(\SUMB[25][29] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_24_29 ( .A(\ab[24][29] ), .B(\CARRYB[23][29] ), .CI(\SUMB[23][30] ), 
        .CO(\CARRYB[24][29] ), .S(\SUMB[24][29] ) );
  FA1A S2_24_30 ( .A(\ab[24][30] ), .B(\CARRYB[23][30] ), .CI(\SUMB[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_23_30 ( .A(\ab[23][30] ), .B(\CARRYB[22][30] ), .CI(\SUMB[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_23_29 ( .A(\ab[23][29] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA1A S2_22_30 ( .A(\ab[22][30] ), .B(\CARRYB[21][30] ), .CI(\SUMB[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA1A S2_22_29 ( .A(\ab[22][29] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA1A S2_21_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\SUMB[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA1A S2_21_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA1A S2_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\SUMB[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA1A S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA1A S2_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\SUMB[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA1A S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA1A S2_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\SUMB[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA1A S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA1A S2_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\SUMB[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA1A S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA1A S2_14_68 ( .A(\ab[14][68] ), .B(\CARRYB[13][68] ), .CI(\SUMB[13][69] ), 
        .CO(\CARRYB[14][68] ), .S(\SUMB[14][68] ) );
  FA1A S2_14_67 ( .A(\ab[14][67] ), .B(\CARRYB[13][67] ), .CI(\SUMB[13][68] ), 
        .CO(\CARRYB[14][67] ), .S(\SUMB[14][67] ) );
  FA1A S2_14_66 ( .A(\ab[14][66] ), .B(\CARRYB[13][66] ), .CI(\SUMB[13][67] ), 
        .CO(\CARRYB[14][66] ), .S(\SUMB[14][66] ) );
  FA1A S2_14_65 ( .A(\ab[14][65] ), .B(\CARRYB[13][65] ), .CI(\SUMB[13][66] ), 
        .CO(\CARRYB[14][65] ), .S(\SUMB[14][65] ) );
  FA1A S2_14_64 ( .A(\ab[14][64] ), .B(\CARRYB[13][64] ), .CI(\SUMB[13][65] ), 
        .CO(\CARRYB[14][64] ), .S(\SUMB[14][64] ) );
  FA1A S2_14_60 ( .A(\ab[14][60] ), .B(\CARRYB[13][60] ), .CI(\SUMB[13][61] ), 
        .CO(\CARRYB[14][60] ), .S(\SUMB[14][60] ) );
  FA1A S2_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\SUMB[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA1A S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA1A S2_13_68 ( .A(\ab[13][68] ), .B(\CARRYB[12][68] ), .CI(\SUMB[12][69] ), 
        .CO(\CARRYB[13][68] ), .S(\SUMB[13][68] ) );
  FA1A S2_13_67 ( .A(\ab[13][67] ), .B(\CARRYB[12][67] ), .CI(\SUMB[12][68] ), 
        .CO(\CARRYB[13][67] ), .S(\SUMB[13][67] ) );
  FA1A S2_13_66 ( .A(\ab[13][66] ), .B(\CARRYB[12][66] ), .CI(\SUMB[12][67] ), 
        .CO(\CARRYB[13][66] ), .S(\SUMB[13][66] ) );
  FA1A S2_13_65 ( .A(\ab[13][65] ), .B(\CARRYB[12][65] ), .CI(\SUMB[12][66] ), 
        .CO(\CARRYB[13][65] ), .S(\SUMB[13][65] ) );
  FA1A S2_13_64 ( .A(\ab[13][64] ), .B(\CARRYB[12][64] ), .CI(\SUMB[12][65] ), 
        .CO(\CARRYB[13][64] ), .S(\SUMB[13][64] ) );
  FA1A S2_13_60 ( .A(\ab[13][60] ), .B(\CARRYB[12][60] ), .CI(\SUMB[12][61] ), 
        .CO(\CARRYB[13][60] ), .S(\SUMB[13][60] ) );
  FA1A S2_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\SUMB[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA1A S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA1A S2_12_68 ( .A(\ab[12][68] ), .B(\CARRYB[11][68] ), .CI(\SUMB[11][69] ), 
        .CO(\CARRYB[12][68] ), .S(\SUMB[12][68] ) );
  FA1A S2_12_67 ( .A(\ab[12][67] ), .B(\CARRYB[11][67] ), .CI(\SUMB[11][68] ), 
        .CO(\CARRYB[12][67] ), .S(\SUMB[12][67] ) );
  FA1A S2_12_66 ( .A(\ab[12][66] ), .B(\CARRYB[11][66] ), .CI(\SUMB[11][67] ), 
        .CO(\CARRYB[12][66] ), .S(\SUMB[12][66] ) );
  FA1A S2_12_65 ( .A(\ab[12][65] ), .B(\CARRYB[11][65] ), .CI(\SUMB[11][66] ), 
        .CO(\CARRYB[12][65] ), .S(\SUMB[12][65] ) );
  FA1A S2_12_64 ( .A(\ab[12][64] ), .B(\CARRYB[11][64] ), .CI(\SUMB[11][65] ), 
        .CO(\CARRYB[12][64] ), .S(\SUMB[12][64] ) );
  FA1A S2_12_60 ( .A(\ab[12][60] ), .B(\CARRYB[11][60] ), .CI(\SUMB[11][61] ), 
        .CO(\CARRYB[12][60] ), .S(\SUMB[12][60] ) );
  FA1A S2_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\SUMB[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA1A S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA1A S2_11_68 ( .A(\ab[11][68] ), .B(\CARRYB[10][68] ), .CI(\SUMB[10][69] ), 
        .CO(\CARRYB[11][68] ), .S(\SUMB[11][68] ) );
  FA1A S2_11_67 ( .A(\ab[11][67] ), .B(\CARRYB[10][67] ), .CI(\SUMB[10][68] ), 
        .CO(\CARRYB[11][67] ), .S(\SUMB[11][67] ) );
  FA1A S2_11_66 ( .A(\ab[11][66] ), .B(\CARRYB[10][66] ), .CI(\SUMB[10][67] ), 
        .CO(\CARRYB[11][66] ), .S(\SUMB[11][66] ) );
  FA1A S2_11_65 ( .A(\ab[11][65] ), .B(\CARRYB[10][65] ), .CI(\SUMB[10][66] ), 
        .CO(\CARRYB[11][65] ), .S(\SUMB[11][65] ) );
  FA1A S2_11_64 ( .A(\ab[11][64] ), .B(\CARRYB[10][64] ), .CI(\SUMB[10][65] ), 
        .CO(\CARRYB[11][64] ), .S(\SUMB[11][64] ) );
  FA1A S2_11_60 ( .A(\ab[11][60] ), .B(\CARRYB[10][60] ), .CI(\SUMB[10][61] ), 
        .CO(\CARRYB[11][60] ), .S(\SUMB[11][60] ) );
  FA1A S2_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\SUMB[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA1A S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA1A S2_10_68 ( .A(\ab[10][68] ), .B(\CARRYB[9][68] ), .CI(\SUMB[9][69] ), 
        .CO(\CARRYB[10][68] ), .S(\SUMB[10][68] ) );
  FA1A S2_10_67 ( .A(\ab[10][67] ), .B(\CARRYB[9][67] ), .CI(\SUMB[9][68] ), 
        .CO(\CARRYB[10][67] ), .S(\SUMB[10][67] ) );
  FA1A S2_10_66 ( .A(\ab[10][66] ), .B(\CARRYB[9][66] ), .CI(\SUMB[9][67] ), 
        .CO(\CARRYB[10][66] ), .S(\SUMB[10][66] ) );
  FA1A S2_10_65 ( .A(\ab[10][65] ), .B(\CARRYB[9][65] ), .CI(\SUMB[9][66] ), 
        .CO(\CARRYB[10][65] ), .S(\SUMB[10][65] ) );
  FA1A S2_10_64 ( .A(\ab[10][64] ), .B(\CARRYB[9][64] ), .CI(\SUMB[9][65] ), 
        .CO(\CARRYB[10][64] ), .S(\SUMB[10][64] ) );
  FA1A S2_10_60 ( .A(\ab[10][60] ), .B(\CARRYB[9][60] ), .CI(\SUMB[9][61] ), 
        .CO(\CARRYB[10][60] ), .S(\SUMB[10][60] ) );
  FA1A S2_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\SUMB[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA1A S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA1A S2_9_68 ( .A(\ab[9][68] ), .B(\CARRYB[8][68] ), .CI(\SUMB[8][69] ), 
        .CO(\CARRYB[9][68] ), .S(\SUMB[9][68] ) );
  FA1A S2_9_67 ( .A(\ab[9][67] ), .B(\CARRYB[8][67] ), .CI(\SUMB[8][68] ), 
        .CO(\CARRYB[9][67] ), .S(\SUMB[9][67] ) );
  FA1A S2_9_66 ( .A(\ab[9][66] ), .B(\CARRYB[8][66] ), .CI(\SUMB[8][67] ), 
        .CO(\CARRYB[9][66] ), .S(\SUMB[9][66] ) );
  FA1A S2_9_65 ( .A(\ab[9][65] ), .B(\CARRYB[8][65] ), .CI(\SUMB[8][66] ), 
        .CO(\CARRYB[9][65] ), .S(\SUMB[9][65] ) );
  FA1A S2_9_64 ( .A(\ab[9][64] ), .B(\CARRYB[8][64] ), .CI(\SUMB[8][65] ), 
        .CO(\CARRYB[9][64] ), .S(\SUMB[9][64] ) );
  FA1A S2_9_60 ( .A(\ab[9][60] ), .B(\CARRYB[8][60] ), .CI(\SUMB[8][61] ), 
        .CO(\CARRYB[9][60] ), .S(\SUMB[9][60] ) );
  FA1A S2_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\SUMB[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA1A S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1A S2_8_68 ( .A(\ab[8][68] ), .B(\CARRYB[7][68] ), .CI(\SUMB[7][69] ), 
        .CO(\CARRYB[8][68] ), .S(\SUMB[8][68] ) );
  FA1A S2_8_67 ( .A(\ab[8][67] ), .B(\CARRYB[7][67] ), .CI(\SUMB[7][68] ), 
        .CO(\CARRYB[8][67] ), .S(\SUMB[8][67] ) );
  FA1A S2_8_66 ( .A(\ab[8][66] ), .B(\CARRYB[7][66] ), .CI(\SUMB[7][67] ), 
        .CO(\CARRYB[8][66] ), .S(\SUMB[8][66] ) );
  FA1A S2_8_65 ( .A(\ab[8][65] ), .B(\CARRYB[7][65] ), .CI(\SUMB[7][66] ), 
        .CO(\CARRYB[8][65] ), .S(\SUMB[8][65] ) );
  FA1A S2_8_64 ( .A(\ab[8][64] ), .B(\CARRYB[7][64] ), .CI(\SUMB[7][65] ), 
        .CO(\CARRYB[8][64] ), .S(\SUMB[8][64] ) );
  FA1A S2_8_60 ( .A(\ab[8][60] ), .B(\CARRYB[7][60] ), .CI(\SUMB[7][61] ), 
        .CO(\CARRYB[8][60] ), .S(\SUMB[8][60] ) );
  FA1A S2_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\SUMB[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA1A S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1A S2_7_68 ( .A(\ab[7][68] ), .B(\CARRYB[6][68] ), .CI(\SUMB[6][69] ), 
        .CO(\CARRYB[7][68] ), .S(\SUMB[7][68] ) );
  FA1A S2_7_67 ( .A(\ab[7][67] ), .B(\CARRYB[6][67] ), .CI(\SUMB[6][68] ), 
        .CO(\CARRYB[7][67] ), .S(\SUMB[7][67] ) );
  FA1A S2_7_66 ( .A(\ab[7][66] ), .B(\CARRYB[6][66] ), .CI(\SUMB[6][67] ), 
        .CO(\CARRYB[7][66] ), .S(\SUMB[7][66] ) );
  FA1A S2_7_65 ( .A(\ab[7][65] ), .B(\CARRYB[6][65] ), .CI(\SUMB[6][66] ), 
        .CO(\CARRYB[7][65] ), .S(\SUMB[7][65] ) );
  FA1A S2_7_64 ( .A(\ab[7][64] ), .B(\CARRYB[6][64] ), .CI(\SUMB[6][65] ), 
        .CO(\CARRYB[7][64] ), .S(\SUMB[7][64] ) );
  FA1A S2_7_60 ( .A(\ab[7][60] ), .B(\CARRYB[6][60] ), .CI(\SUMB[6][61] ), 
        .CO(\CARRYB[7][60] ), .S(\SUMB[7][60] ) );
  FA1A S2_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\SUMB[8][31] ), 
        .CO(\CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA1A S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1A S2_6_68 ( .A(\ab[6][68] ), .B(\CARRYB[5][68] ), .CI(\SUMB[5][69] ), 
        .CO(\CARRYB[6][68] ), .S(\SUMB[6][68] ) );
  FA1A S2_6_67 ( .A(\ab[6][67] ), .B(\CARRYB[5][67] ), .CI(\SUMB[5][68] ), 
        .CO(\CARRYB[6][67] ), .S(\SUMB[6][67] ) );
  FA1A S2_6_66 ( .A(\ab[6][66] ), .B(\CARRYB[5][66] ), .CI(\SUMB[5][67] ), 
        .CO(\CARRYB[6][66] ), .S(\SUMB[6][66] ) );
  FA1A S2_6_65 ( .A(\ab[6][65] ), .B(\CARRYB[5][65] ), .CI(\SUMB[5][66] ), 
        .CO(\CARRYB[6][65] ), .S(\SUMB[6][65] ) );
  FA1A S2_6_64 ( .A(\ab[6][64] ), .B(\CARRYB[5][64] ), .CI(\SUMB[5][65] ), 
        .CO(\CARRYB[6][64] ), .S(\SUMB[6][64] ) );
  FA1A S2_6_60 ( .A(\ab[6][60] ), .B(\CARRYB[5][60] ), .CI(\SUMB[5][61] ), 
        .CO(\CARRYB[6][60] ), .S(\SUMB[6][60] ) );
  FA1A S2_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\SUMB[7][31] ), 
        .CO(\CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA1A S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1A S2_5_68 ( .A(\ab[5][68] ), .B(\CARRYB[4][68] ), .CI(\SUMB[4][69] ), 
        .CO(\CARRYB[5][68] ), .S(\SUMB[5][68] ) );
  FA1A S2_5_67 ( .A(\ab[5][67] ), .B(\CARRYB[4][67] ), .CI(\SUMB[4][68] ), 
        .CO(\CARRYB[5][67] ), .S(\SUMB[5][67] ) );
  FA1A S2_5_66 ( .A(\ab[5][66] ), .B(\CARRYB[4][66] ), .CI(\SUMB[4][67] ), 
        .CO(\CARRYB[5][66] ), .S(\SUMB[5][66] ) );
  FA1A S2_5_65 ( .A(\ab[5][65] ), .B(\CARRYB[4][65] ), .CI(\SUMB[4][66] ), 
        .CO(\CARRYB[5][65] ), .S(\SUMB[5][65] ) );
  FA1A S2_5_64 ( .A(\ab[5][64] ), .B(\CARRYB[4][64] ), .CI(\SUMB[4][65] ), 
        .CO(\CARRYB[5][64] ), .S(\SUMB[5][64] ) );
  FA1A S2_5_60 ( .A(\ab[5][60] ), .B(\CARRYB[4][60] ), .CI(\SUMB[4][61] ), 
        .CO(\CARRYB[5][60] ), .S(\SUMB[5][60] ) );
  FA1A S2_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\SUMB[6][31] ), 
        .CO(\CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA1A S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1A S2_4_68 ( .A(\ab[4][68] ), .B(\CARRYB[3][68] ), .CI(\SUMB[3][69] ), 
        .CO(\CARRYB[4][68] ), .S(\SUMB[4][68] ) );
  FA1A S2_4_67 ( .A(\ab[4][67] ), .B(\CARRYB[3][67] ), .CI(\SUMB[3][68] ), 
        .CO(\CARRYB[4][67] ), .S(\SUMB[4][67] ) );
  FA1A S2_4_66 ( .A(\ab[4][66] ), .B(\CARRYB[3][66] ), .CI(\SUMB[3][67] ), 
        .CO(\CARRYB[4][66] ), .S(\SUMB[4][66] ) );
  FA1A S2_4_65 ( .A(\ab[4][65] ), .B(\CARRYB[3][65] ), .CI(\SUMB[3][66] ), 
        .CO(\CARRYB[4][65] ), .S(\SUMB[4][65] ) );
  FA1A S2_4_64 ( .A(\ab[4][64] ), .B(\CARRYB[3][64] ), .CI(\SUMB[3][65] ), 
        .CO(\CARRYB[4][64] ), .S(\SUMB[4][64] ) );
  FA1A S2_4_60 ( .A(\ab[4][60] ), .B(\CARRYB[3][60] ), .CI(\SUMB[3][61] ), 
        .CO(\CARRYB[4][60] ), .S(\SUMB[4][60] ) );
  FA1A S2_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\SUMB[5][31] ), 
        .CO(\CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA1A S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA1A S2_3_68 ( .A(\ab[3][68] ), .B(\CARRYB[2][68] ), .CI(\SUMB[2][69] ), 
        .CO(\CARRYB[3][68] ), .S(\SUMB[3][68] ) );
  FA1A S2_3_67 ( .A(\ab[3][67] ), .B(\CARRYB[2][67] ), .CI(\SUMB[2][68] ), 
        .CO(\CARRYB[3][67] ), .S(\SUMB[3][67] ) );
  FA1A S2_3_66 ( .A(\ab[3][66] ), .B(\CARRYB[2][66] ), .CI(\SUMB[2][67] ), 
        .CO(\CARRYB[3][66] ), .S(\SUMB[3][66] ) );
  FA1A S2_3_65 ( .A(\ab[3][65] ), .B(\CARRYB[2][65] ), .CI(\SUMB[2][66] ), 
        .CO(\CARRYB[3][65] ), .S(\SUMB[3][65] ) );
  FA1A S2_3_64 ( .A(\ab[3][64] ), .B(\CARRYB[2][64] ), .CI(\SUMB[2][65] ), 
        .CO(\CARRYB[3][64] ), .S(\SUMB[3][64] ) );
  FA1A S2_3_60 ( .A(\ab[3][60] ), .B(\CARRYB[2][60] ), .CI(\SUMB[2][61] ), 
        .CO(\CARRYB[3][60] ), .S(\SUMB[3][60] ) );
  FA1A S2_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\SUMB[4][31] ), 
        .CO(\CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA1A S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA1A S2_2_68 ( .A(\ab[2][68] ), .B(\CARRYB[1][68] ), .CI(\SUMB[1][69] ), 
        .CO(\CARRYB[2][68] ), .S(\SUMB[2][68] ) );
  FA1A S2_2_67 ( .A(\ab[2][67] ), .B(\CARRYB[1][67] ), .CI(\SUMB[1][68] ), 
        .CO(\CARRYB[2][67] ), .S(\SUMB[2][67] ) );
  FA1A S2_2_66 ( .A(\ab[2][66] ), .B(\CARRYB[1][66] ), .CI(\SUMB[1][67] ), 
        .CO(\CARRYB[2][66] ), .S(\SUMB[2][66] ) );
  FA1A S2_2_65 ( .A(\ab[2][65] ), .B(\CARRYB[1][65] ), .CI(\SUMB[1][66] ), 
        .CO(\CARRYB[2][65] ), .S(\SUMB[2][65] ) );
  FA1A S2_2_64 ( .A(\ab[2][64] ), .B(\CARRYB[1][64] ), .CI(\SUMB[1][65] ), 
        .CO(\CARRYB[2][64] ), .S(\SUMB[2][64] ) );
  FA1A S2_2_60 ( .A(\ab[2][60] ), .B(\CARRYB[1][60] ), .CI(\SUMB[1][61] ), 
        .CO(\CARRYB[2][60] ), .S(\SUMB[2][60] ) );
  FA1A S2_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\SUMB[3][31] ), 
        .CO(\CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA1A S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\SUMB[3][30] ), 
        .CO(\CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1A S2_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .CI(\SUMB[2][31] ), 
        .CO(\CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA1A S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1A S2_2_30 ( .A(\ab[2][30] ), .B(\CARRYB[1][30] ), .CI(\SUMB[1][31] ), 
        .CO(\CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  FA1A S2_2_29 ( .A(\ab[2][29] ), .B(\CARRYB[1][29] ), .CI(\SUMB[1][30] ), 
        .CO(\CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1A S4_33 ( .A(\ab[29][33] ), .B(\CARRYB[28][33] ), .CI(\SUMB[28][34] ), 
        .CO(\CARRYB[29][33] ), .S(\SUMB[29][33] ) );
  FA1A S4_34 ( .A(\ab[29][34] ), .B(\CARRYB[28][34] ), .CI(\SUMB[28][35] ), 
        .CO(\CARRYB[29][34] ), .S(\SUMB[29][34] ) );
  FA1A S4_31 ( .A(\ab[29][31] ), .B(\CARRYB[28][31] ), .CI(\SUMB[28][32] ), 
        .CO(\CARRYB[29][31] ), .S(\SUMB[29][31] ) );
  FA1A S2_28_33 ( .A(\ab[28][33] ), .B(\CARRYB[27][33] ), .CI(\SUMB[27][34] ), 
        .CO(\CARRYB[28][33] ), .S(\SUMB[28][33] ) );
  FA1A S2_28_32 ( .A(\ab[28][32] ), .B(\CARRYB[27][32] ), .CI(\SUMB[27][33] ), 
        .CO(\CARRYB[28][32] ), .S(\SUMB[28][32] ) );
  FA1A S2_28_34 ( .A(\ab[28][34] ), .B(\CARRYB[27][34] ), .CI(\SUMB[27][35] ), 
        .CO(\CARRYB[28][34] ), .S(\SUMB[28][34] ) );
  FA1A S4_37 ( .A(\ab[29][37] ), .B(\CARRYB[28][37] ), .CI(\SUMB[28][38] ), 
        .CO(\CARRYB[29][37] ), .S(\SUMB[29][37] ) );
  FA1A S2_27_34 ( .A(\ab[27][34] ), .B(\CARRYB[26][34] ), .CI(\SUMB[26][35] ), 
        .CO(\CARRYB[27][34] ), .S(\SUMB[27][34] ) );
  FA1A S2_27_33 ( .A(\ab[27][33] ), .B(\CARRYB[26][33] ), .CI(\SUMB[26][34] ), 
        .CO(\CARRYB[27][33] ), .S(\SUMB[27][33] ) );
  FA1A S2_28_37 ( .A(\ab[28][37] ), .B(\CARRYB[27][37] ), .CI(\SUMB[27][38] ), 
        .CO(\CARRYB[28][37] ), .S(\SUMB[28][37] ) );
  FA1A S2_28_36 ( .A(\ab[28][36] ), .B(\CARRYB[27][36] ), .CI(\SUMB[27][37] ), 
        .CO(\CARRYB[28][36] ), .S(\SUMB[28][36] ) );
  FA1A S2_28_35 ( .A(\ab[28][35] ), .B(\CARRYB[27][35] ), .CI(\SUMB[27][36] ), 
        .CO(\CARRYB[28][35] ), .S(\SUMB[28][35] ) );
  FA1A S2_26_34 ( .A(\ab[26][34] ), .B(\CARRYB[25][34] ), .CI(\SUMB[25][35] ), 
        .CO(\CARRYB[26][34] ), .S(\SUMB[26][34] ) );
  FA1A S2_28_31 ( .A(\ab[28][31] ), .B(\CARRYB[27][31] ), .CI(\SUMB[27][32] ), 
        .CO(\CARRYB[28][31] ), .S(\SUMB[28][31] ) );
  FA1A S4_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), .CO(
        \CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA1A S2_27_37 ( .A(\ab[27][37] ), .B(\CARRYB[26][37] ), .CI(\SUMB[26][38] ), 
        .CO(\CARRYB[27][37] ), .S(\SUMB[27][37] ) );
  FA1A S2_27_36 ( .A(\ab[27][36] ), .B(\CARRYB[26][36] ), .CI(\SUMB[26][37] ), 
        .CO(\CARRYB[27][36] ), .S(\SUMB[27][36] ) );
  FA1A S2_27_35 ( .A(\ab[27][35] ), .B(\CARRYB[26][35] ), .CI(\SUMB[26][36] ), 
        .CO(\CARRYB[27][35] ), .S(\SUMB[27][35] ) );
  FA1A S2_27_32 ( .A(\ab[27][32] ), .B(\CARRYB[26][32] ), .CI(\SUMB[26][33] ), 
        .CO(\CARRYB[27][32] ), .S(\SUMB[27][32] ) );
  FA1A S2_27_31 ( .A(\ab[27][31] ), .B(\CARRYB[26][31] ), .CI(\SUMB[26][32] ), 
        .CO(\CARRYB[27][31] ), .S(\SUMB[27][31] ) );
  FA1A S4_27 ( .A(\ab[29][27] ), .B(\CARRYB[28][27] ), .CI(\SUMB[28][28] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA1A S4_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), .CO(
        \CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA1A S4_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), .CO(
        \CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA1A S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA1A S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA1A S2_26_37 ( .A(\ab[26][37] ), .B(\CARRYB[25][37] ), .CI(\SUMB[25][38] ), 
        .CO(\CARRYB[26][37] ), .S(\SUMB[26][37] ) );
  FA1A S2_26_36 ( .A(\ab[26][36] ), .B(\CARRYB[25][36] ), .CI(\SUMB[25][37] ), 
        .CO(\CARRYB[26][36] ), .S(\SUMB[26][36] ) );
  FA1A S2_28_38 ( .A(\ab[28][38] ), .B(\CARRYB[27][38] ), .CI(\SUMB[27][39] ), 
        .CO(\CARRYB[28][38] ), .S(\SUMB[28][38] ) );
  FA1A S2_26_35 ( .A(\ab[26][35] ), .B(\CARRYB[25][35] ), .CI(\SUMB[25][36] ), 
        .CO(\CARRYB[26][35] ), .S(\SUMB[26][35] ) );
  FA1A S2_26_33 ( .A(\ab[26][33] ), .B(\CARRYB[25][33] ), .CI(\SUMB[25][34] ), 
        .CO(\CARRYB[26][33] ), .S(\SUMB[26][33] ) );
  FA1A S2_26_32 ( .A(\ab[26][32] ), .B(\CARRYB[25][32] ), .CI(\SUMB[25][33] ), 
        .CO(\CARRYB[26][32] ), .S(\SUMB[26][32] ) );
  FA1A S2_26_31 ( .A(\ab[26][31] ), .B(\CARRYB[25][31] ), .CI(\SUMB[25][32] ), 
        .CO(\CARRYB[26][31] ), .S(\SUMB[26][31] ) );
  FA1A S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA1A S2_28_28 ( .A(\ab[28][28] ), .B(\CARRYB[27][28] ), .CI(\SUMB[27][29] ), 
        .CO(\CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA1A S4_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA1A S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA1A S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA1A S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA1A S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA1A S2_25_37 ( .A(\ab[25][37] ), .B(\CARRYB[24][37] ), .CI(\SUMB[24][38] ), 
        .CO(\CARRYB[25][37] ), .S(\SUMB[25][37] ) );
  FA1A S2_25_36 ( .A(\ab[25][36] ), .B(\CARRYB[24][36] ), .CI(\SUMB[24][37] ), 
        .CO(\CARRYB[25][36] ), .S(\SUMB[25][36] ) );
  FA1A S2_27_38 ( .A(\ab[27][38] ), .B(\CARRYB[26][38] ), .CI(\SUMB[26][39] ), 
        .CO(\CARRYB[27][38] ), .S(\SUMB[27][38] ) );
  FA1A S2_25_35 ( .A(\ab[25][35] ), .B(\CARRYB[24][35] ), .CI(\SUMB[24][36] ), 
        .CO(\CARRYB[25][35] ), .S(\SUMB[25][35] ) );
  FA1A S2_25_34 ( .A(\ab[25][34] ), .B(\CARRYB[24][34] ), .CI(\SUMB[24][35] ), 
        .CO(\CARRYB[25][34] ), .S(\SUMB[25][34] ) );
  FA1A S2_25_33 ( .A(\ab[25][33] ), .B(\CARRYB[24][33] ), .CI(\SUMB[24][34] ), 
        .CO(\CARRYB[25][33] ), .S(\SUMB[25][33] ) );
  FA1A S2_25_32 ( .A(\ab[25][32] ), .B(\CARRYB[24][32] ), .CI(\SUMB[24][33] ), 
        .CO(\CARRYB[25][32] ), .S(\SUMB[25][32] ) );
  FA1A S2_27_28 ( .A(\ab[27][28] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), 
        .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FA1A S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA1A S2_28_26 ( .A(\ab[28][26] ), .B(\CARRYB[27][26] ), .CI(\SUMB[27][27] ), 
        .CO(\CARRYB[28][26] ), .S(\SUMB[28][26] ) );
  FA1A S4_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA1A S4_22 ( .A(\ab[29][22] ), .B(\CARRYB[28][22] ), .CI(\SUMB[28][23] ), 
        .CO(\CARRYB[29][22] ), .S(\SUMB[29][22] ) );
  FA1A S4_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA1A S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA1A S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA1A S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA1A S2_28_7 ( .A(\ab[28][7] ), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA1A S2_28_6 ( .A(\ab[28][6] ), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA1A S2_24_37 ( .A(\ab[24][37] ), .B(\CARRYB[23][37] ), .CI(\SUMB[23][38] ), 
        .CO(\CARRYB[24][37] ), .S(\SUMB[24][37] ) );
  FA1A S2_24_36 ( .A(\ab[24][36] ), .B(\CARRYB[23][36] ), .CI(\SUMB[23][37] ), 
        .CO(\CARRYB[24][36] ), .S(\SUMB[24][36] ) );
  FA1A S2_26_38 ( .A(\ab[26][38] ), .B(\CARRYB[25][38] ), .CI(\SUMB[25][39] ), 
        .CO(\CARRYB[26][38] ), .S(\SUMB[26][38] ) );
  FA1A S2_24_35 ( .A(\ab[24][35] ), .B(\CARRYB[23][35] ), .CI(\SUMB[23][36] ), 
        .CO(\CARRYB[24][35] ), .S(\SUMB[24][35] ) );
  FA1A S2_24_34 ( .A(\ab[24][34] ), .B(\CARRYB[23][34] ), .CI(\SUMB[23][35] ), 
        .CO(\CARRYB[24][34] ), .S(\SUMB[24][34] ) );
  FA1A S2_24_33 ( .A(\ab[24][33] ), .B(\CARRYB[23][33] ), .CI(\SUMB[23][34] ), 
        .CO(\CARRYB[24][33] ), .S(\SUMB[24][33] ) );
  FA1A S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA1A S2_27_27 ( .A(\ab[27][27] ), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), 
        .CO(\CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA1A S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA1A S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA1A S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA1A S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA1A S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA1A S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA1A S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA1A S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA1A S2_27_7 ( .A(\ab[27][7] ), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA1A S2_27_6 ( .A(\ab[27][6] ), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA1A S2_23_37 ( .A(\ab[23][37] ), .B(\CARRYB[22][37] ), .CI(\SUMB[22][38] ), 
        .CO(\CARRYB[23][37] ), .S(\SUMB[23][37] ) );
  FA1A S2_23_36 ( .A(\ab[23][36] ), .B(\CARRYB[22][36] ), .CI(\SUMB[22][37] ), 
        .CO(\CARRYB[23][36] ), .S(\SUMB[23][36] ) );
  FA1A S2_25_38 ( .A(\ab[25][38] ), .B(\CARRYB[24][38] ), .CI(\SUMB[24][39] ), 
        .CO(\CARRYB[25][38] ), .S(\SUMB[25][38] ) );
  FA1A S2_23_35 ( .A(\ab[23][35] ), .B(\CARRYB[22][35] ), .CI(\SUMB[22][36] ), 
        .CO(\CARRYB[23][35] ), .S(\SUMB[23][35] ) );
  FA1A S2_23_34 ( .A(\ab[23][34] ), .B(\CARRYB[22][34] ), .CI(\SUMB[22][35] ), 
        .CO(\CARRYB[23][34] ), .S(\SUMB[23][34] ) );
  FA1A S2_25_31 ( .A(\ab[25][31] ), .B(\CARRYB[24][31] ), .CI(\SUMB[24][32] ), 
        .CO(\CARRYB[25][31] ), .S(\SUMB[25][31] ) );
  FA1A S2_26_27 ( .A(\ab[26][27] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), 
        .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FA1A S2_26_28 ( .A(\ab[26][28] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), 
        .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FA1A S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA1A S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA1A S2_27_23 ( .A(\ab[27][23] ), .B(\CARRYB[26][23] ), .CI(\SUMB[26][24] ), 
        .CO(\CARRYB[27][23] ), .S(\SUMB[27][23] ) );
  FA1A S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), 
        .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FA1A S2_27_21 ( .A(\ab[27][21] ), .B(\CARRYB[26][21] ), .CI(\SUMB[26][22] ), 
        .CO(\CARRYB[27][21] ), .S(\SUMB[27][21] ) );
  FA1A S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA1A S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA1A S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA1A S2_26_8 ( .A(\ab[26][8] ), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA1A S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA1A S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA1A S2_22_37 ( .A(\ab[22][37] ), .B(\CARRYB[21][37] ), .CI(\SUMB[21][38] ), 
        .CO(\CARRYB[22][37] ), .S(\SUMB[22][37] ) );
  FA1A S2_22_36 ( .A(\ab[22][36] ), .B(\CARRYB[21][36] ), .CI(\SUMB[21][37] ), 
        .CO(\CARRYB[22][36] ), .S(\SUMB[22][36] ) );
  FA1A S2_24_38 ( .A(\ab[24][38] ), .B(\CARRYB[23][38] ), .CI(\SUMB[23][39] ), 
        .CO(\CARRYB[24][38] ), .S(\SUMB[24][38] ) );
  FA1A S2_22_35 ( .A(\ab[22][35] ), .B(\CARRYB[21][35] ), .CI(\SUMB[21][36] ), 
        .CO(\CARRYB[22][35] ), .S(\SUMB[22][35] ) );
  FA1A S2_24_31 ( .A(\ab[24][31] ), .B(\CARRYB[23][31] ), .CI(\SUMB[23][32] ), 
        .CO(\CARRYB[24][31] ), .S(\SUMB[24][31] ) );
  FA1A S2_24_32 ( .A(\ab[24][32] ), .B(\CARRYB[23][32] ), .CI(\SUMB[23][33] ), 
        .CO(\CARRYB[24][32] ), .S(\SUMB[24][32] ) );
  FA1A S2_25_28 ( .A(\ab[25][28] ), .B(\CARRYB[24][28] ), .CI(\SUMB[24][29] ), 
        .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FA1A S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), 
        .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA1A S2_26_25 ( .A(\ab[26][25] ), .B(\CARRYB[25][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA1A S2_26_24 ( .A(\ab[26][24] ), .B(\CARRYB[25][24] ), .CI(\SUMB[25][25] ), 
        .CO(\CARRYB[26][24] ), .S(\SUMB[26][24] ) );
  FA1A S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA1A S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA1A S2_26_21 ( .A(\ab[26][21] ), .B(\CARRYB[25][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA1A S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA1A S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA1A S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA1A S2_25_8 ( .A(\ab[25][8] ), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA1A S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA1A S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA1A S2_21_37 ( .A(\ab[21][37] ), .B(\CARRYB[20][37] ), .CI(\SUMB[20][38] ), 
        .CO(\CARRYB[21][37] ), .S(\SUMB[21][37] ) );
  FA1A S2_21_36 ( .A(\ab[21][36] ), .B(\CARRYB[20][36] ), .CI(\SUMB[20][37] ), 
        .CO(\CARRYB[21][36] ), .S(\SUMB[21][36] ) );
  FA1A S2_23_38 ( .A(\ab[23][38] ), .B(\CARRYB[22][38] ), .CI(\SUMB[22][39] ), 
        .CO(\CARRYB[23][38] ), .S(\SUMB[23][38] ) );
  FA1A S2_23_32 ( .A(\ab[23][32] ), .B(\CARRYB[22][32] ), .CI(\SUMB[22][33] ), 
        .CO(\CARRYB[23][32] ), .S(\SUMB[23][32] ) );
  FA1A S2_23_33 ( .A(\ab[23][33] ), .B(\CARRYB[22][33] ), .CI(\SUMB[22][34] ), 
        .CO(\CARRYB[23][33] ), .S(\SUMB[23][33] ) );
  FA1A S2_25_27 ( .A(\ab[25][27] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA1A S2_25_26 ( .A(\ab[25][26] ), .B(\CARRYB[24][26] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA1A S2_25_25 ( .A(\ab[25][25] ), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), 
        .CO(\CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA1A S2_25_24 ( .A(\ab[25][24] ), .B(\CARRYB[24][24] ), .CI(\SUMB[24][25] ), 
        .CO(\CARRYB[25][24] ), .S(\SUMB[25][24] ) );
  FA1A S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA1A S2_25_22 ( .A(\ab[25][22] ), .B(\CARRYB[24][22] ), .CI(\SUMB[24][23] ), 
        .CO(\CARRYB[25][22] ), .S(\SUMB[25][22] ) );
  FA1A S2_25_21 ( .A(\ab[25][21] ), .B(\CARRYB[24][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA1A S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA1A S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA1A S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA1A S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA1A S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA1A S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA1A S2_20_37 ( .A(\ab[20][37] ), .B(\CARRYB[19][37] ), .CI(\SUMB[19][38] ), 
        .CO(\CARRYB[20][37] ), .S(\SUMB[20][37] ) );
  FA1A S2_22_38 ( .A(\ab[22][38] ), .B(\CARRYB[21][38] ), .CI(\SUMB[21][39] ), 
        .CO(\CARRYB[22][38] ), .S(\SUMB[22][38] ) );
  FA1A S2_22_33 ( .A(\ab[22][33] ), .B(\CARRYB[21][33] ), .CI(\SUMB[21][34] ), 
        .CO(\CARRYB[22][33] ), .S(\SUMB[22][33] ) );
  FA1A S2_22_34 ( .A(\ab[22][34] ), .B(\CARRYB[21][34] ), .CI(\SUMB[21][35] ), 
        .CO(\CARRYB[22][34] ), .S(\SUMB[22][34] ) );
  FA1A S2_23_31 ( .A(\ab[23][31] ), .B(\CARRYB[22][31] ), .CI(\SUMB[22][32] ), 
        .CO(\CARRYB[23][31] ), .S(\SUMB[23][31] ) );
  FA1A S2_24_28 ( .A(\ab[24][28] ), .B(\CARRYB[23][28] ), .CI(\SUMB[23][29] ), 
        .CO(\CARRYB[24][28] ), .S(\SUMB[24][28] ) );
  FA1A S2_24_27 ( .A(\ab[24][27] ), .B(\CARRYB[23][27] ), .CI(\SUMB[23][28] ), 
        .CO(\CARRYB[24][27] ), .S(\SUMB[24][27] ) );
  FA1A S2_24_26 ( .A(\ab[24][26] ), .B(\CARRYB[23][26] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA1A S2_24_25 ( .A(\ab[24][25] ), .B(\CARRYB[23][25] ), .CI(\SUMB[23][26] ), 
        .CO(\CARRYB[24][25] ), .S(\SUMB[24][25] ) );
  FA1A S2_24_24 ( .A(\ab[24][24] ), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), 
        .CO(\CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA1A S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA1A S2_24_22 ( .A(\ab[24][22] ), .B(\CARRYB[23][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA1A S2_24_21 ( .A(\ab[24][21] ), .B(\CARRYB[23][21] ), .CI(\SUMB[23][22] ), 
        .CO(\CARRYB[24][21] ), .S(\SUMB[24][21] ) );
  FA1A S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA1A S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1A S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1A S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA1A S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA1A S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA1A S2_21_38 ( .A(\ab[21][38] ), .B(\CARRYB[20][38] ), .CI(\SUMB[20][39] ), 
        .CO(\CARRYB[21][38] ), .S(\SUMB[21][38] ) );
  FA1A S2_21_34 ( .A(\ab[21][34] ), .B(\CARRYB[20][34] ), .CI(\SUMB[20][35] ), 
        .CO(\CARRYB[21][34] ), .S(\SUMB[21][34] ) );
  FA1A S2_21_35 ( .A(\ab[21][35] ), .B(\CARRYB[20][35] ), .CI(\SUMB[20][36] ), 
        .CO(\CARRYB[21][35] ), .S(\SUMB[21][35] ) );
  FA1A S2_22_31 ( .A(\ab[22][31] ), .B(\CARRYB[21][31] ), .CI(\SUMB[21][32] ), 
        .CO(\CARRYB[22][31] ), .S(\SUMB[22][31] ) );
  FA1A S2_22_32 ( .A(\ab[22][32] ), .B(\CARRYB[21][32] ), .CI(\SUMB[21][33] ), 
        .CO(\CARRYB[22][32] ), .S(\SUMB[22][32] ) );
  FA1A S2_23_28 ( .A(\ab[23][28] ), .B(\CARRYB[22][28] ), .CI(\SUMB[22][29] ), 
        .CO(\CARRYB[23][28] ), .S(\SUMB[23][28] ) );
  FA1A S2_23_27 ( .A(\ab[23][27] ), .B(\CARRYB[22][27] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA1A S2_23_26 ( .A(\ab[23][26] ), .B(\CARRYB[22][26] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA1A S2_23_25 ( .A(\ab[23][25] ), .B(\CARRYB[22][25] ), .CI(\SUMB[22][26] ), 
        .CO(\CARRYB[23][25] ), .S(\SUMB[23][25] ) );
  FA1A S2_23_24 ( .A(\ab[23][24] ), .B(\CARRYB[22][24] ), .CI(\SUMB[22][25] ), 
        .CO(\CARRYB[23][24] ), .S(\SUMB[23][24] ) );
  FA1A S2_23_23 ( .A(\ab[23][23] ), .B(\CARRYB[22][23] ), .CI(\SUMB[22][24] ), 
        .CO(\CARRYB[23][23] ), .S(\SUMB[23][23] ) );
  FA1A S2_23_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA1A S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA1A S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1A S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1A S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA1A S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA1A S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA1A S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA1A S2_20_38 ( .A(\ab[20][38] ), .B(\CARRYB[19][38] ), .CI(\SUMB[19][39] ), 
        .CO(\CARRYB[20][38] ), .S(\SUMB[20][38] ) );
  FA1A S2_20_35 ( .A(\ab[20][35] ), .B(\CARRYB[19][35] ), .CI(\SUMB[19][36] ), 
        .CO(\CARRYB[20][35] ), .S(\SUMB[20][35] ) );
  FA1A S2_20_36 ( .A(\ab[20][36] ), .B(\CARRYB[19][36] ), .CI(\SUMB[19][37] ), 
        .CO(\CARRYB[20][36] ), .S(\SUMB[20][36] ) );
  FA1A S2_21_32 ( .A(\ab[21][32] ), .B(\CARRYB[20][32] ), .CI(\SUMB[20][33] ), 
        .CO(\CARRYB[21][32] ), .S(\SUMB[21][32] ) );
  FA1A S2_21_33 ( .A(\ab[21][33] ), .B(\CARRYB[20][33] ), .CI(\SUMB[20][34] ), 
        .CO(\CARRYB[21][33] ), .S(\SUMB[21][33] ) );
  FA1A S2_22_28 ( .A(\ab[22][28] ), .B(\CARRYB[21][28] ), .CI(\SUMB[21][29] ), 
        .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FA1A S2_22_27 ( .A(\ab[22][27] ), .B(\CARRYB[21][27] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA1A S2_22_26 ( .A(\ab[22][26] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA1A S2_22_25 ( .A(\ab[22][25] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA1A S2_22_24 ( .A(\ab[22][24] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA1A S2_22_23 ( .A(\ab[22][23] ), .B(\CARRYB[21][23] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA1A S2_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA1A S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA1A S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA1A S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1A S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1A S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1A S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA1A S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA1A S2_19_38 ( .A(\ab[19][38] ), .B(\CARRYB[18][38] ), .CI(\SUMB[18][39] ), 
        .CO(\CARRYB[19][38] ), .S(\SUMB[19][38] ) );
  FA1A S2_19_36 ( .A(\ab[19][36] ), .B(\CARRYB[18][36] ), .CI(\SUMB[18][37] ), 
        .CO(\CARRYB[19][36] ), .S(\SUMB[19][36] ) );
  FA1A S2_19_37 ( .A(\ab[19][37] ), .B(\CARRYB[18][37] ), .CI(\SUMB[18][38] ), 
        .CO(\CARRYB[19][37] ), .S(\SUMB[19][37] ) );
  FA1A S2_20_33 ( .A(\ab[20][33] ), .B(\CARRYB[19][33] ), .CI(\SUMB[19][34] ), 
        .CO(\CARRYB[20][33] ), .S(\SUMB[20][33] ) );
  FA1A S2_20_34 ( .A(\ab[20][34] ), .B(\CARRYB[19][34] ), .CI(\SUMB[19][35] ), 
        .CO(\CARRYB[20][34] ), .S(\SUMB[20][34] ) );
  FA1A S2_21_31 ( .A(\ab[21][31] ), .B(\CARRYB[20][31] ), .CI(\SUMB[20][32] ), 
        .CO(\CARRYB[21][31] ), .S(\SUMB[21][31] ) );
  FA1A S2_21_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA1A S2_21_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA1A S2_21_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA1A S2_21_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA1A S2_21_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA1A S2_21_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA1A S2_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA1A S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA1A S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1A S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1A S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1A S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA1A S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1A S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1A S2_18_38 ( .A(\ab[18][38] ), .B(\CARRYB[17][38] ), .CI(\SUMB[17][39] ), 
        .CO(\CARRYB[18][38] ), .S(\SUMB[18][38] ) );
  FA1A S2_18_37 ( .A(\ab[18][37] ), .B(\CARRYB[17][37] ), .CI(\SUMB[17][38] ), 
        .CO(\CARRYB[18][37] ), .S(\SUMB[18][37] ) );
  FA1A S2_19_34 ( .A(\ab[19][34] ), .B(\CARRYB[18][34] ), .CI(\SUMB[18][35] ), 
        .CO(\CARRYB[19][34] ), .S(\SUMB[19][34] ) );
  FA1A S2_19_35 ( .A(\ab[19][35] ), .B(\CARRYB[18][35] ), .CI(\SUMB[18][36] ), 
        .CO(\CARRYB[19][35] ), .S(\SUMB[19][35] ) );
  FA1A S2_20_32 ( .A(\ab[20][32] ), .B(\CARRYB[19][32] ), .CI(\SUMB[19][33] ), 
        .CO(\CARRYB[20][32] ), .S(\SUMB[20][32] ) );
  FA1A S2_20_31 ( .A(\ab[20][31] ), .B(\CARRYB[19][31] ), .CI(\SUMB[19][32] ), 
        .CO(\CARRYB[20][31] ), .S(\SUMB[20][31] ) );
  FA1A S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA1A S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA1A S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA1A S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA1A S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA1A S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA1A S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA1A S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA1A S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA1A S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1A S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1A S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1A S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA1A S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1A S2_17_38 ( .A(\ab[17][38] ), .B(\CARRYB[16][38] ), .CI(\SUMB[16][39] ), 
        .CO(\CARRYB[17][38] ), .S(\SUMB[17][38] ) );
  FA1A S2_18_35 ( .A(\ab[18][35] ), .B(\CARRYB[17][35] ), .CI(\SUMB[17][36] ), 
        .CO(\CARRYB[18][35] ), .S(\SUMB[18][35] ) );
  FA1A S2_18_36 ( .A(\ab[18][36] ), .B(\CARRYB[17][36] ), .CI(\SUMB[17][37] ), 
        .CO(\CARRYB[18][36] ), .S(\SUMB[18][36] ) );
  FA1A S2_19_33 ( .A(\ab[19][33] ), .B(\CARRYB[18][33] ), .CI(\SUMB[18][34] ), 
        .CO(\CARRYB[19][33] ), .S(\SUMB[19][33] ) );
  FA1A S2_19_32 ( .A(\ab[19][32] ), .B(\CARRYB[18][32] ), .CI(\SUMB[18][33] ), 
        .CO(\CARRYB[19][32] ), .S(\SUMB[19][32] ) );
  FA1A S2_19_31 ( .A(\ab[19][31] ), .B(\CARRYB[18][31] ), .CI(\SUMB[18][32] ), 
        .CO(\CARRYB[19][31] ), .S(\SUMB[19][31] ) );
  FA1A S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA1A S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA1A S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA1A S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA1A S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA1A S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA1A S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA1A S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA1A S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1A S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1A S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1A S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA1A S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1A S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA1A S2_17_36 ( .A(\ab[17][36] ), .B(\CARRYB[16][36] ), .CI(\SUMB[16][37] ), 
        .CO(\CARRYB[17][36] ), .S(\SUMB[17][36] ) );
  FA1A S2_17_37 ( .A(\ab[17][37] ), .B(\CARRYB[16][37] ), .CI(\SUMB[16][38] ), 
        .CO(\CARRYB[17][37] ), .S(\SUMB[17][37] ) );
  FA1A S2_18_34 ( .A(\ab[18][34] ), .B(\CARRYB[17][34] ), .CI(\SUMB[17][35] ), 
        .CO(\CARRYB[18][34] ), .S(\SUMB[18][34] ) );
  FA1A S2_18_33 ( .A(\ab[18][33] ), .B(\CARRYB[17][33] ), .CI(\SUMB[17][34] ), 
        .CO(\CARRYB[18][33] ), .S(\SUMB[18][33] ) );
  FA1A S2_18_32 ( .A(\ab[18][32] ), .B(\CARRYB[17][32] ), .CI(\SUMB[17][33] ), 
        .CO(\CARRYB[18][32] ), .S(\SUMB[18][32] ) );
  FA1A S2_18_31 ( .A(\ab[18][31] ), .B(\CARRYB[17][31] ), .CI(\SUMB[17][32] ), 
        .CO(\CARRYB[18][31] ), .S(\SUMB[18][31] ) );
  FA1A S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA1A S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA1A S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA1A S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA1A S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA1A S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA1A S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA1A S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA1A S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1A S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1A S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1A S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1A S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1A S2_16_37 ( .A(\ab[16][37] ), .B(\CARRYB[15][37] ), .CI(\SUMB[15][38] ), 
        .CO(\CARRYB[16][37] ), .S(\SUMB[16][37] ) );
  FA1A S2_16_38 ( .A(\ab[16][38] ), .B(\CARRYB[15][38] ), .CI(\SUMB[15][39] ), 
        .CO(\CARRYB[16][38] ), .S(\SUMB[16][38] ) );
  FA1A S2_17_35 ( .A(\ab[17][35] ), .B(\CARRYB[16][35] ), .CI(\SUMB[16][36] ), 
        .CO(\CARRYB[17][35] ), .S(\SUMB[17][35] ) );
  FA1A S2_17_34 ( .A(\ab[17][34] ), .B(\CARRYB[16][34] ), .CI(\SUMB[16][35] ), 
        .CO(\CARRYB[17][34] ), .S(\SUMB[17][34] ) );
  FA1A S2_17_33 ( .A(\ab[17][33] ), .B(\CARRYB[16][33] ), .CI(\SUMB[16][34] ), 
        .CO(\CARRYB[17][33] ), .S(\SUMB[17][33] ) );
  FA1A S2_17_32 ( .A(\ab[17][32] ), .B(\CARRYB[16][32] ), .CI(\SUMB[16][33] ), 
        .CO(\CARRYB[17][32] ), .S(\SUMB[17][32] ) );
  FA1A S2_17_31 ( .A(\ab[17][31] ), .B(\CARRYB[16][31] ), .CI(\SUMB[16][32] ), 
        .CO(\CARRYB[17][31] ), .S(\SUMB[17][31] ) );
  FA1A S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA1A S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA1A S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA1A S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA1A S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA1A S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA1A S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA1A S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA1A S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1A S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1A S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1A S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1A S2_14_63 ( .A(\ab[14][63] ), .B(\CARRYB[13][63] ), .CI(\SUMB[13][64] ), 
        .CO(\CARRYB[14][63] ), .S(\SUMB[14][63] ) );
  FA1A S2_14_62 ( .A(\ab[14][62] ), .B(\CARRYB[13][62] ), .CI(\SUMB[13][63] ), 
        .CO(\CARRYB[14][62] ), .S(\SUMB[14][62] ) );
  FA1A S2_14_61 ( .A(\ab[14][61] ), .B(\CARRYB[13][61] ), .CI(\SUMB[13][62] ), 
        .CO(\CARRYB[14][61] ), .S(\SUMB[14][61] ) );
  FA1A S2_16_36 ( .A(\ab[16][36] ), .B(\CARRYB[15][36] ), .CI(\SUMB[15][37] ), 
        .CO(\CARRYB[16][36] ), .S(\SUMB[16][36] ) );
  FA1A S2_16_35 ( .A(\ab[16][35] ), .B(\CARRYB[15][35] ), .CI(\SUMB[15][36] ), 
        .CO(\CARRYB[16][35] ), .S(\SUMB[16][35] ) );
  FA1A S2_16_34 ( .A(\ab[16][34] ), .B(\CARRYB[15][34] ), .CI(\SUMB[15][35] ), 
        .CO(\CARRYB[16][34] ), .S(\SUMB[16][34] ) );
  FA1A S2_16_33 ( .A(\ab[16][33] ), .B(\CARRYB[15][33] ), .CI(\SUMB[15][34] ), 
        .CO(\CARRYB[16][33] ), .S(\SUMB[16][33] ) );
  FA1A S2_16_32 ( .A(\ab[16][32] ), .B(\CARRYB[15][32] ), .CI(\SUMB[15][33] ), 
        .CO(\CARRYB[16][32] ), .S(\SUMB[16][32] ) );
  FA1A S2_16_31 ( .A(\ab[16][31] ), .B(\CARRYB[15][31] ), .CI(\SUMB[15][32] ), 
        .CO(\CARRYB[16][31] ), .S(\SUMB[16][31] ) );
  FA1A S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA1A S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA1A S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA1A S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA1A S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA1A S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA1A S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA1A S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA1A S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1A S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1A S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA1A S2_13_63 ( .A(\ab[13][63] ), .B(\CARRYB[12][63] ), .CI(\SUMB[12][64] ), 
        .CO(\CARRYB[13][63] ), .S(\SUMB[13][63] ) );
  FA1A S2_13_62 ( .A(\ab[13][62] ), .B(\CARRYB[12][62] ), .CI(\SUMB[12][63] ), 
        .CO(\CARRYB[13][62] ), .S(\SUMB[13][62] ) );
  FA1A S2_13_61 ( .A(\ab[13][61] ), .B(\CARRYB[12][61] ), .CI(\SUMB[12][62] ), 
        .CO(\CARRYB[13][61] ), .S(\SUMB[13][61] ) );
  FA1A S2_15_37 ( .A(\ab[15][37] ), .B(\CARRYB[14][37] ), .CI(\SUMB[14][38] ), 
        .CO(\CARRYB[15][37] ), .S(\SUMB[15][37] ) );
  FA1A S2_15_36 ( .A(\ab[15][36] ), .B(\CARRYB[14][36] ), .CI(\SUMB[14][37] ), 
        .CO(\CARRYB[15][36] ), .S(\SUMB[15][36] ) );
  FA1A S2_15_35 ( .A(\ab[15][35] ), .B(\CARRYB[14][35] ), .CI(\SUMB[14][36] ), 
        .CO(\CARRYB[15][35] ), .S(\SUMB[15][35] ) );
  FA1A S2_15_34 ( .A(\ab[15][34] ), .B(\CARRYB[14][34] ), .CI(\SUMB[14][35] ), 
        .CO(\CARRYB[15][34] ), .S(\SUMB[15][34] ) );
  FA1A S2_15_33 ( .A(\ab[15][33] ), .B(\CARRYB[14][33] ), .CI(\SUMB[14][34] ), 
        .CO(\CARRYB[15][33] ), .S(\SUMB[15][33] ) );
  FA1A S2_15_32 ( .A(\ab[15][32] ), .B(\CARRYB[14][32] ), .CI(\SUMB[14][33] ), 
        .CO(\CARRYB[15][32] ), .S(\SUMB[15][32] ) );
  FA1A S2_15_31 ( .A(\ab[15][31] ), .B(\CARRYB[14][31] ), .CI(\SUMB[14][32] ), 
        .CO(\CARRYB[15][31] ), .S(\SUMB[15][31] ) );
  FA1A S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA1A S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA1A S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA1A S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA1A S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA1A S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA1A S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA1A S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S2_12_63 ( .A(\ab[12][63] ), .B(\CARRYB[11][63] ), .CI(\SUMB[11][64] ), 
        .CO(\CARRYB[12][63] ), .S(\SUMB[12][63] ) );
  FA1A S2_12_62 ( .A(\ab[12][62] ), .B(\CARRYB[11][62] ), .CI(\SUMB[11][63] ), 
        .CO(\CARRYB[12][62] ), .S(\SUMB[12][62] ) );
  FA1A S2_12_61 ( .A(\ab[12][61] ), .B(\CARRYB[11][61] ), .CI(\SUMB[11][62] ), 
        .CO(\CARRYB[12][61] ), .S(\SUMB[12][61] ) );
  FA1A S2_14_37 ( .A(\ab[14][37] ), .B(\CARRYB[13][37] ), .CI(\SUMB[13][38] ), 
        .CO(\CARRYB[14][37] ), .S(\SUMB[14][37] ) );
  FA1A S2_14_36 ( .A(\ab[14][36] ), .B(\CARRYB[13][36] ), .CI(\SUMB[13][37] ), 
        .CO(\CARRYB[14][36] ), .S(\SUMB[14][36] ) );
  FA1A S2_14_35 ( .A(\ab[14][35] ), .B(\CARRYB[13][35] ), .CI(\SUMB[13][36] ), 
        .CO(\CARRYB[14][35] ), .S(\SUMB[14][35] ) );
  FA1A S2_14_34 ( .A(\ab[14][34] ), .B(\CARRYB[13][34] ), .CI(\SUMB[13][35] ), 
        .CO(\CARRYB[14][34] ), .S(\SUMB[14][34] ) );
  FA1A S2_14_33 ( .A(\ab[14][33] ), .B(\CARRYB[13][33] ), .CI(\SUMB[13][34] ), 
        .CO(\CARRYB[14][33] ), .S(\SUMB[14][33] ) );
  FA1A S2_14_32 ( .A(\ab[14][32] ), .B(\CARRYB[13][32] ), .CI(\SUMB[13][33] ), 
        .CO(\CARRYB[14][32] ), .S(\SUMB[14][32] ) );
  FA1A S2_14_31 ( .A(\ab[14][31] ), .B(\CARRYB[13][31] ), .CI(\SUMB[13][32] ), 
        .CO(\CARRYB[14][31] ), .S(\SUMB[14][31] ) );
  FA1A S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA1A S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA1A S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA1A S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA1A S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA1A S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA1A S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA1A S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_11_63 ( .A(\ab[11][63] ), .B(\CARRYB[10][63] ), .CI(\SUMB[10][64] ), 
        .CO(\CARRYB[11][63] ), .S(\SUMB[11][63] ) );
  FA1A S2_11_62 ( .A(\ab[11][62] ), .B(\CARRYB[10][62] ), .CI(\SUMB[10][63] ), 
        .CO(\CARRYB[11][62] ), .S(\SUMB[11][62] ) );
  FA1A S2_11_61 ( .A(\ab[11][61] ), .B(\CARRYB[10][61] ), .CI(\SUMB[10][62] ), 
        .CO(\CARRYB[11][61] ), .S(\SUMB[11][61] ) );
  FA1A S2_13_37 ( .A(\ab[13][37] ), .B(\CARRYB[12][37] ), .CI(\SUMB[12][38] ), 
        .CO(\CARRYB[13][37] ), .S(\SUMB[13][37] ) );
  FA1A S2_13_36 ( .A(\ab[13][36] ), .B(\CARRYB[12][36] ), .CI(\SUMB[12][37] ), 
        .CO(\CARRYB[13][36] ), .S(\SUMB[13][36] ) );
  FA1A S2_13_35 ( .A(\ab[13][35] ), .B(\CARRYB[12][35] ), .CI(\SUMB[12][36] ), 
        .CO(\CARRYB[13][35] ), .S(\SUMB[13][35] ) );
  FA1A S2_13_34 ( .A(\ab[13][34] ), .B(\CARRYB[12][34] ), .CI(\SUMB[12][35] ), 
        .CO(\CARRYB[13][34] ), .S(\SUMB[13][34] ) );
  FA1A S2_13_33 ( .A(\ab[13][33] ), .B(\CARRYB[12][33] ), .CI(\SUMB[12][34] ), 
        .CO(\CARRYB[13][33] ), .S(\SUMB[13][33] ) );
  FA1A S2_13_32 ( .A(\ab[13][32] ), .B(\CARRYB[12][32] ), .CI(\SUMB[12][33] ), 
        .CO(\CARRYB[13][32] ), .S(\SUMB[13][32] ) );
  FA1A S2_13_31 ( .A(\ab[13][31] ), .B(\CARRYB[12][31] ), .CI(\SUMB[12][32] ), 
        .CO(\CARRYB[13][31] ), .S(\SUMB[13][31] ) );
  FA1A S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA1A S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA1A S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA1A S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA1A S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA1A S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA1A S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA1A S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_10_63 ( .A(\ab[10][63] ), .B(\CARRYB[9][63] ), .CI(\SUMB[9][64] ), 
        .CO(\CARRYB[10][63] ), .S(\SUMB[10][63] ) );
  FA1A S2_10_62 ( .A(\ab[10][62] ), .B(\CARRYB[9][62] ), .CI(\SUMB[9][63] ), 
        .CO(\CARRYB[10][62] ), .S(\SUMB[10][62] ) );
  FA1A S2_10_61 ( .A(\ab[10][61] ), .B(\CARRYB[9][61] ), .CI(\SUMB[9][62] ), 
        .CO(\CARRYB[10][61] ), .S(\SUMB[10][61] ) );
  FA1A S2_12_37 ( .A(\ab[12][37] ), .B(\CARRYB[11][37] ), .CI(\SUMB[11][38] ), 
        .CO(\CARRYB[12][37] ), .S(\SUMB[12][37] ) );
  FA1A S2_12_36 ( .A(\ab[12][36] ), .B(\CARRYB[11][36] ), .CI(\SUMB[11][37] ), 
        .CO(\CARRYB[12][36] ), .S(\SUMB[12][36] ) );
  FA1A S2_12_35 ( .A(\ab[12][35] ), .B(\CARRYB[11][35] ), .CI(\SUMB[11][36] ), 
        .CO(\CARRYB[12][35] ), .S(\SUMB[12][35] ) );
  FA1A S2_12_34 ( .A(\ab[12][34] ), .B(\CARRYB[11][34] ), .CI(\SUMB[11][35] ), 
        .CO(\CARRYB[12][34] ), .S(\SUMB[12][34] ) );
  FA1A S2_12_33 ( .A(\ab[12][33] ), .B(\CARRYB[11][33] ), .CI(\SUMB[11][34] ), 
        .CO(\CARRYB[12][33] ), .S(\SUMB[12][33] ) );
  FA1A S2_12_32 ( .A(\ab[12][32] ), .B(\CARRYB[11][32] ), .CI(\SUMB[11][33] ), 
        .CO(\CARRYB[12][32] ), .S(\SUMB[12][32] ) );
  FA1A S2_12_31 ( .A(\ab[12][31] ), .B(\CARRYB[11][31] ), .CI(\SUMB[11][32] ), 
        .CO(\CARRYB[12][31] ), .S(\SUMB[12][31] ) );
  FA1A S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA1A S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA1A S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA1A S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA1A S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA1A S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA1A S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA1A S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_9_63 ( .A(\ab[9][63] ), .B(\CARRYB[8][63] ), .CI(\SUMB[8][64] ), 
        .CO(\CARRYB[9][63] ), .S(\SUMB[9][63] ) );
  FA1A S2_9_62 ( .A(\ab[9][62] ), .B(\CARRYB[8][62] ), .CI(\SUMB[8][63] ), 
        .CO(\CARRYB[9][62] ), .S(\SUMB[9][62] ) );
  FA1A S2_9_61 ( .A(\ab[9][61] ), .B(\CARRYB[8][61] ), .CI(\SUMB[8][62] ), 
        .CO(\CARRYB[9][61] ), .S(\SUMB[9][61] ) );
  FA1A S2_11_37 ( .A(\ab[11][37] ), .B(\CARRYB[10][37] ), .CI(\SUMB[10][38] ), 
        .CO(\CARRYB[11][37] ), .S(\SUMB[11][37] ) );
  FA1A S2_11_36 ( .A(\ab[11][36] ), .B(\CARRYB[10][36] ), .CI(\SUMB[10][37] ), 
        .CO(\CARRYB[11][36] ), .S(\SUMB[11][36] ) );
  FA1A S2_11_35 ( .A(\ab[11][35] ), .B(\CARRYB[10][35] ), .CI(\SUMB[10][36] ), 
        .CO(\CARRYB[11][35] ), .S(\SUMB[11][35] ) );
  FA1A S2_11_34 ( .A(\ab[11][34] ), .B(\CARRYB[10][34] ), .CI(\SUMB[10][35] ), 
        .CO(\CARRYB[11][34] ), .S(\SUMB[11][34] ) );
  FA1A S2_11_33 ( .A(\ab[11][33] ), .B(\CARRYB[10][33] ), .CI(\SUMB[10][34] ), 
        .CO(\CARRYB[11][33] ), .S(\SUMB[11][33] ) );
  FA1A S2_11_32 ( .A(\ab[11][32] ), .B(\CARRYB[10][32] ), .CI(\SUMB[10][33] ), 
        .CO(\CARRYB[11][32] ), .S(\SUMB[11][32] ) );
  FA1A S2_11_31 ( .A(\ab[11][31] ), .B(\CARRYB[10][31] ), .CI(\SUMB[10][32] ), 
        .CO(\CARRYB[11][31] ), .S(\SUMB[11][31] ) );
  FA1A S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1A S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA1A S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1A S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1A S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1A S2_11_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1A S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1A S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_8_63 ( .A(\ab[8][63] ), .B(\CARRYB[7][63] ), .CI(\SUMB[7][64] ), 
        .CO(\CARRYB[8][63] ), .S(\SUMB[8][63] ) );
  FA1A S2_8_62 ( .A(\ab[8][62] ), .B(\CARRYB[7][62] ), .CI(\SUMB[7][63] ), 
        .CO(\CARRYB[8][62] ), .S(\SUMB[8][62] ) );
  FA1A S2_8_61 ( .A(\ab[8][61] ), .B(\CARRYB[7][61] ), .CI(\SUMB[7][62] ), 
        .CO(\CARRYB[8][61] ), .S(\SUMB[8][61] ) );
  FA1A S2_10_37 ( .A(\ab[10][37] ), .B(\CARRYB[9][37] ), .CI(\SUMB[9][38] ), 
        .CO(\CARRYB[10][37] ), .S(\SUMB[10][37] ) );
  FA1A S2_10_36 ( .A(\ab[10][36] ), .B(\CARRYB[9][36] ), .CI(\SUMB[9][37] ), 
        .CO(\CARRYB[10][36] ), .S(\SUMB[10][36] ) );
  FA1A S2_10_35 ( .A(\ab[10][35] ), .B(\CARRYB[9][35] ), .CI(\SUMB[9][36] ), 
        .CO(\CARRYB[10][35] ), .S(\SUMB[10][35] ) );
  FA1A S2_10_34 ( .A(\ab[10][34] ), .B(\CARRYB[9][34] ), .CI(\SUMB[9][35] ), 
        .CO(\CARRYB[10][34] ), .S(\SUMB[10][34] ) );
  FA1A S2_10_33 ( .A(\ab[10][33] ), .B(\CARRYB[9][33] ), .CI(\SUMB[9][34] ), 
        .CO(\CARRYB[10][33] ), .S(\SUMB[10][33] ) );
  FA1A S2_10_32 ( .A(\ab[10][32] ), .B(\CARRYB[9][32] ), .CI(\SUMB[9][33] ), 
        .CO(\CARRYB[10][32] ), .S(\SUMB[10][32] ) );
  FA1A S2_10_31 ( .A(\ab[10][31] ), .B(\CARRYB[9][31] ), .CI(\SUMB[9][32] ), 
        .CO(\CARRYB[10][31] ), .S(\SUMB[10][31] ) );
  FA1A S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1A S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA1A S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA1A S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1A S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1A S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA1A S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA1A S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_7_63 ( .A(\ab[7][63] ), .B(\CARRYB[6][63] ), .CI(\SUMB[6][64] ), 
        .CO(\CARRYB[7][63] ), .S(\SUMB[7][63] ) );
  FA1A S2_7_62 ( .A(\ab[7][62] ), .B(\CARRYB[6][62] ), .CI(\SUMB[6][63] ), 
        .CO(\CARRYB[7][62] ), .S(\SUMB[7][62] ) );
  FA1A S2_7_61 ( .A(\ab[7][61] ), .B(\CARRYB[6][61] ), .CI(\SUMB[6][62] ), 
        .CO(\CARRYB[7][61] ), .S(\SUMB[7][61] ) );
  FA1A S2_9_37 ( .A(\ab[9][37] ), .B(\CARRYB[8][37] ), .CI(\SUMB[8][38] ), 
        .CO(\CARRYB[9][37] ), .S(\SUMB[9][37] ) );
  FA1A S2_9_36 ( .A(\ab[9][36] ), .B(\CARRYB[8][36] ), .CI(\SUMB[8][37] ), 
        .CO(\CARRYB[9][36] ), .S(\SUMB[9][36] ) );
  FA1A S2_9_35 ( .A(\ab[9][35] ), .B(\CARRYB[8][35] ), .CI(\SUMB[8][36] ), 
        .CO(\CARRYB[9][35] ), .S(\SUMB[9][35] ) );
  FA1A S2_9_34 ( .A(\ab[9][34] ), .B(\CARRYB[8][34] ), .CI(\SUMB[8][35] ), 
        .CO(\CARRYB[9][34] ), .S(\SUMB[9][34] ) );
  FA1A S2_9_33 ( .A(\ab[9][33] ), .B(\CARRYB[8][33] ), .CI(\SUMB[8][34] ), 
        .CO(\CARRYB[9][33] ), .S(\SUMB[9][33] ) );
  FA1A S2_9_32 ( .A(\ab[9][32] ), .B(\CARRYB[8][32] ), .CI(\SUMB[8][33] ), 
        .CO(\CARRYB[9][32] ), .S(\SUMB[9][32] ) );
  FA1A S2_9_31 ( .A(\ab[9][31] ), .B(\CARRYB[8][31] ), .CI(\SUMB[8][32] ), 
        .CO(\CARRYB[9][31] ), .S(\SUMB[9][31] ) );
  FA1A S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1A S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1A S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1A S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1A S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1A S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA1A S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_6_63 ( .A(\ab[6][63] ), .B(\CARRYB[5][63] ), .CI(\SUMB[5][64] ), 
        .CO(\CARRYB[6][63] ), .S(\SUMB[6][63] ) );
  FA1A S2_6_62 ( .A(\ab[6][62] ), .B(\CARRYB[5][62] ), .CI(\SUMB[5][63] ), 
        .CO(\CARRYB[6][62] ), .S(\SUMB[6][62] ) );
  FA1A S2_6_61 ( .A(\ab[6][61] ), .B(\CARRYB[5][61] ), .CI(\SUMB[5][62] ), 
        .CO(\CARRYB[6][61] ), .S(\SUMB[6][61] ) );
  FA1A S2_8_37 ( .A(\ab[8][37] ), .B(\CARRYB[7][37] ), .CI(\SUMB[7][38] ), 
        .CO(\CARRYB[8][37] ), .S(\SUMB[8][37] ) );
  FA1A S2_8_36 ( .A(\ab[8][36] ), .B(\CARRYB[7][36] ), .CI(\SUMB[7][37] ), 
        .CO(\CARRYB[8][36] ), .S(\SUMB[8][36] ) );
  FA1A S2_8_35 ( .A(\ab[8][35] ), .B(\CARRYB[7][35] ), .CI(\SUMB[7][36] ), 
        .CO(\CARRYB[8][35] ), .S(\SUMB[8][35] ) );
  FA1A S2_8_34 ( .A(\ab[8][34] ), .B(\CARRYB[7][34] ), .CI(\SUMB[7][35] ), 
        .CO(\CARRYB[8][34] ), .S(\SUMB[8][34] ) );
  FA1A S2_8_33 ( .A(\ab[8][33] ), .B(\CARRYB[7][33] ), .CI(\SUMB[7][34] ), 
        .CO(\CARRYB[8][33] ), .S(\SUMB[8][33] ) );
  FA1A S2_8_32 ( .A(\ab[8][32] ), .B(\CARRYB[7][32] ), .CI(\SUMB[7][33] ), 
        .CO(\CARRYB[8][32] ), .S(\SUMB[8][32] ) );
  FA1A S2_8_31 ( .A(\ab[8][31] ), .B(\CARRYB[7][31] ), .CI(\SUMB[7][32] ), 
        .CO(\CARRYB[8][31] ), .S(\SUMB[8][31] ) );
  FA1A S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA1A S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1A S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1A S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1A S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1A S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1A S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1A S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_5_63 ( .A(\ab[5][63] ), .B(\CARRYB[4][63] ), .CI(\SUMB[4][64] ), 
        .CO(\CARRYB[5][63] ), .S(\SUMB[5][63] ) );
  FA1A S2_5_62 ( .A(\ab[5][62] ), .B(\CARRYB[4][62] ), .CI(\SUMB[4][63] ), 
        .CO(\CARRYB[5][62] ), .S(\SUMB[5][62] ) );
  FA1A S2_5_61 ( .A(\ab[5][61] ), .B(\CARRYB[4][61] ), .CI(\SUMB[4][62] ), 
        .CO(\CARRYB[5][61] ), .S(\SUMB[5][61] ) );
  FA1A S2_7_37 ( .A(\ab[7][37] ), .B(\CARRYB[6][37] ), .CI(\SUMB[6][38] ), 
        .CO(\CARRYB[7][37] ), .S(\SUMB[7][37] ) );
  FA1A S2_7_36 ( .A(\ab[7][36] ), .B(\CARRYB[6][36] ), .CI(\SUMB[6][37] ), 
        .CO(\CARRYB[7][36] ), .S(\SUMB[7][36] ) );
  FA1A S2_7_35 ( .A(\ab[7][35] ), .B(\CARRYB[6][35] ), .CI(\SUMB[6][36] ), 
        .CO(\CARRYB[7][35] ), .S(\SUMB[7][35] ) );
  FA1A S2_7_34 ( .A(\ab[7][34] ), .B(\CARRYB[6][34] ), .CI(\SUMB[6][35] ), 
        .CO(\CARRYB[7][34] ), .S(\SUMB[7][34] ) );
  FA1A S2_7_33 ( .A(\ab[7][33] ), .B(\CARRYB[6][33] ), .CI(\SUMB[6][34] ), 
        .CO(\CARRYB[7][33] ), .S(\SUMB[7][33] ) );
  FA1A S2_7_32 ( .A(\ab[7][32] ), .B(\CARRYB[6][32] ), .CI(\SUMB[6][33] ), 
        .CO(\CARRYB[7][32] ), .S(\SUMB[7][32] ) );
  FA1A S2_7_31 ( .A(\ab[7][31] ), .B(\CARRYB[6][31] ), .CI(\SUMB[6][32] ), 
        .CO(\CARRYB[7][31] ), .S(\SUMB[7][31] ) );
  FA1A S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA1A S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1A S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA1A S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA1A S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA1A S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA1A S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA1A S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_4_63 ( .A(\ab[4][63] ), .B(\CARRYB[3][63] ), .CI(\SUMB[3][64] ), 
        .CO(\CARRYB[4][63] ), .S(\SUMB[4][63] ) );
  FA1A S2_4_62 ( .A(\ab[4][62] ), .B(\CARRYB[3][62] ), .CI(\SUMB[3][63] ), 
        .CO(\CARRYB[4][62] ), .S(\SUMB[4][62] ) );
  FA1A S2_4_61 ( .A(\ab[4][61] ), .B(\CARRYB[3][61] ), .CI(\SUMB[3][62] ), 
        .CO(\CARRYB[4][61] ), .S(\SUMB[4][61] ) );
  FA1A S2_6_37 ( .A(\ab[6][37] ), .B(\CARRYB[5][37] ), .CI(\SUMB[5][38] ), 
        .CO(\CARRYB[6][37] ), .S(\SUMB[6][37] ) );
  FA1A S2_6_36 ( .A(\ab[6][36] ), .B(\CARRYB[5][36] ), .CI(\SUMB[5][37] ), 
        .CO(\CARRYB[6][36] ), .S(\SUMB[6][36] ) );
  FA1A S2_6_35 ( .A(\ab[6][35] ), .B(\CARRYB[5][35] ), .CI(\SUMB[5][36] ), 
        .CO(\CARRYB[6][35] ), .S(\SUMB[6][35] ) );
  FA1A S2_6_34 ( .A(\ab[6][34] ), .B(\CARRYB[5][34] ), .CI(\SUMB[5][35] ), 
        .CO(\CARRYB[6][34] ), .S(\SUMB[6][34] ) );
  FA1A S2_6_33 ( .A(\ab[6][33] ), .B(\CARRYB[5][33] ), .CI(\SUMB[5][34] ), 
        .CO(\CARRYB[6][33] ), .S(\SUMB[6][33] ) );
  FA1A S2_6_32 ( .A(\ab[6][32] ), .B(\CARRYB[5][32] ), .CI(\SUMB[5][33] ), 
        .CO(\CARRYB[6][32] ), .S(\SUMB[6][32] ) );
  FA1A S2_6_31 ( .A(\ab[6][31] ), .B(\CARRYB[5][31] ), .CI(\SUMB[5][32] ), 
        .CO(\CARRYB[6][31] ), .S(\SUMB[6][31] ) );
  FA1A S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1A S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA1A S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA1A S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA1A S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1A S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1A S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA1A S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_3_63 ( .A(\ab[3][63] ), .B(\CARRYB[2][63] ), .CI(\SUMB[2][64] ), 
        .CO(\CARRYB[3][63] ), .S(\SUMB[3][63] ) );
  FA1A S2_3_62 ( .A(\ab[3][62] ), .B(\CARRYB[2][62] ), .CI(\SUMB[2][63] ), 
        .CO(\CARRYB[3][62] ), .S(\SUMB[3][62] ) );
  FA1A S2_3_61 ( .A(\ab[3][61] ), .B(\CARRYB[2][61] ), .CI(\SUMB[2][62] ), 
        .CO(\CARRYB[3][61] ), .S(\SUMB[3][61] ) );
  FA1A S2_5_37 ( .A(\ab[5][37] ), .B(\CARRYB[4][37] ), .CI(\SUMB[4][38] ), 
        .CO(\CARRYB[5][37] ), .S(\SUMB[5][37] ) );
  FA1A S2_5_36 ( .A(\ab[5][36] ), .B(\CARRYB[4][36] ), .CI(\SUMB[4][37] ), 
        .CO(\CARRYB[5][36] ), .S(\SUMB[5][36] ) );
  FA1A S2_5_35 ( .A(\ab[5][35] ), .B(\CARRYB[4][35] ), .CI(\SUMB[4][36] ), 
        .CO(\CARRYB[5][35] ), .S(\SUMB[5][35] ) );
  FA1A S2_5_34 ( .A(\ab[5][34] ), .B(\CARRYB[4][34] ), .CI(\SUMB[4][35] ), 
        .CO(\CARRYB[5][34] ), .S(\SUMB[5][34] ) );
  FA1A S2_5_33 ( .A(\ab[5][33] ), .B(\CARRYB[4][33] ), .CI(\SUMB[4][34] ), 
        .CO(\CARRYB[5][33] ), .S(\SUMB[5][33] ) );
  FA1A S2_5_32 ( .A(\ab[5][32] ), .B(\CARRYB[4][32] ), .CI(\SUMB[4][33] ), 
        .CO(\CARRYB[5][32] ), .S(\SUMB[5][32] ) );
  FA1A S2_5_31 ( .A(\ab[5][31] ), .B(\CARRYB[4][31] ), .CI(\SUMB[4][32] ), 
        .CO(\CARRYB[5][31] ), .S(\SUMB[5][31] ) );
  FA1A S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA1A S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA1A S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1A S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1A S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1A S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1A S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_2_63 ( .A(\ab[2][63] ), .B(\CARRYB[1][63] ), .CI(\SUMB[1][64] ), 
        .CO(\CARRYB[2][63] ), .S(\SUMB[2][63] ) );
  FA1A S2_2_62 ( .A(\ab[2][62] ), .B(\CARRYB[1][62] ), .CI(\SUMB[1][63] ), 
        .CO(\CARRYB[2][62] ), .S(\SUMB[2][62] ) );
  FA1A S2_2_61 ( .A(\ab[2][61] ), .B(\CARRYB[1][61] ), .CI(\SUMB[1][62] ), 
        .CO(\CARRYB[2][61] ), .S(\SUMB[2][61] ) );
  FA1A S2_4_37 ( .A(\ab[4][37] ), .B(\CARRYB[3][37] ), .CI(\SUMB[3][38] ), 
        .CO(\CARRYB[4][37] ), .S(\SUMB[4][37] ) );
  FA1A S2_4_36 ( .A(\ab[4][36] ), .B(\CARRYB[3][36] ), .CI(\SUMB[3][37] ), 
        .CO(\CARRYB[4][36] ), .S(\SUMB[4][36] ) );
  FA1A S2_4_35 ( .A(\ab[4][35] ), .B(\CARRYB[3][35] ), .CI(\SUMB[3][36] ), 
        .CO(\CARRYB[4][35] ), .S(\SUMB[4][35] ) );
  FA1A S2_4_34 ( .A(\ab[4][34] ), .B(\CARRYB[3][34] ), .CI(\SUMB[3][35] ), 
        .CO(\CARRYB[4][34] ), .S(\SUMB[4][34] ) );
  FA1A S2_4_33 ( .A(\ab[4][33] ), .B(\CARRYB[3][33] ), .CI(\SUMB[3][34] ), 
        .CO(\CARRYB[4][33] ), .S(\SUMB[4][33] ) );
  FA1A S2_4_32 ( .A(\ab[4][32] ), .B(\CARRYB[3][32] ), .CI(\SUMB[3][33] ), 
        .CO(\CARRYB[4][32] ), .S(\SUMB[4][32] ) );
  FA1A S2_4_31 ( .A(\ab[4][31] ), .B(\CARRYB[3][31] ), .CI(\SUMB[3][32] ), 
        .CO(\CARRYB[4][31] ), .S(\SUMB[4][31] ) );
  FA1A S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1A S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1A S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1A S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1A S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1A S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA1A S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA1A S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_3_37 ( .A(\ab[3][37] ), .B(\CARRYB[2][37] ), .CI(\SUMB[2][38] ), 
        .CO(\CARRYB[3][37] ), .S(\SUMB[3][37] ) );
  FA1A S2_3_36 ( .A(\ab[3][36] ), .B(\CARRYB[2][36] ), .CI(\SUMB[2][37] ), 
        .CO(\CARRYB[3][36] ), .S(\SUMB[3][36] ) );
  FA1A S2_3_35 ( .A(\ab[3][35] ), .B(\CARRYB[2][35] ), .CI(\SUMB[2][36] ), 
        .CO(\CARRYB[3][35] ), .S(\SUMB[3][35] ) );
  FA1A S2_3_34 ( .A(\ab[3][34] ), .B(\CARRYB[2][34] ), .CI(\SUMB[2][35] ), 
        .CO(\CARRYB[3][34] ), .S(\SUMB[3][34] ) );
  FA1A S2_3_33 ( .A(\ab[3][33] ), .B(\CARRYB[2][33] ), .CI(\SUMB[2][34] ), 
        .CO(\CARRYB[3][33] ), .S(\SUMB[3][33] ) );
  FA1A S2_3_32 ( .A(\ab[3][32] ), .B(\CARRYB[2][32] ), .CI(\SUMB[2][33] ), 
        .CO(\CARRYB[3][32] ), .S(\SUMB[3][32] ) );
  FA1A S2_3_31 ( .A(\ab[3][31] ), .B(\CARRYB[2][31] ), .CI(\SUMB[2][32] ), 
        .CO(\CARRYB[3][31] ), .S(\SUMB[3][31] ) );
  FA1A S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA1A S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1A S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1A S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA1A S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA1A S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA1A S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA1A S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_2_36 ( .A(\ab[2][36] ), .B(\CARRYB[1][36] ), .CI(\SUMB[1][37] ), 
        .CO(\CARRYB[2][36] ), .S(\SUMB[2][36] ) );
  FA1A S2_2_35 ( .A(\ab[2][35] ), .B(\CARRYB[1][35] ), .CI(\SUMB[1][36] ), 
        .CO(\CARRYB[2][35] ), .S(\SUMB[2][35] ) );
  FA1A S2_2_34 ( .A(\ab[2][34] ), .B(\CARRYB[1][34] ), .CI(\SUMB[1][35] ), 
        .CO(\CARRYB[2][34] ), .S(\SUMB[2][34] ) );
  FA1A S2_2_33 ( .A(\ab[2][33] ), .B(\CARRYB[1][33] ), .CI(\SUMB[1][34] ), 
        .CO(\CARRYB[2][33] ), .S(\SUMB[2][33] ) );
  FA1A S2_2_32 ( .A(\ab[2][32] ), .B(\CARRYB[1][32] ), .CI(\SUMB[1][33] ), 
        .CO(\CARRYB[2][32] ), .S(\SUMB[2][32] ) );
  FA1A S2_2_31 ( .A(\ab[2][31] ), .B(\CARRYB[1][31] ), .CI(\SUMB[1][32] ), 
        .CO(\CARRYB[2][31] ), .S(\SUMB[2][31] ) );
  FA1A S2_2_28 ( .A(\ab[2][28] ), .B(\CARRYB[1][28] ), .CI(\SUMB[1][29] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FA1A S2_2_27 ( .A(\ab[2][27] ), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1A S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1A S2_2_25 ( .A(\ab[2][25] ), .B(\CARRYB[1][25] ), .CI(\SUMB[1][26] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1A S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), 
        .CO(\CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA1A S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1A S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA1A S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), 
        .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA1A S4_32 ( .A(\ab[29][32] ), .B(\CARRYB[28][32] ), .CI(\SUMB[28][33] ), 
        .CO(\CARRYB[29][32] ), .S(\SUMB[29][32] ) );
  FA1A S4_36 ( .A(\ab[29][36] ), .B(\CARRYB[28][36] ), .CI(\SUMB[28][37] ), 
        .CO(\CARRYB[29][36] ), .S(\SUMB[29][36] ) );
  FA1A S4_35 ( .A(\ab[29][35] ), .B(\CARRYB[28][35] ), .CI(\SUMB[28][36] ), 
        .CO(\CARRYB[29][35] ), .S(\SUMB[29][35] ) );
  FA1A S4_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA1A S4_3 ( .A(\ab[29][3] ), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), .CO(
        \CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA1A S4_38 ( .A(\ab[29][38] ), .B(\CARRYB[28][38] ), .CI(\SUMB[28][39] ), 
        .CO(\CARRYB[29][38] ), .S(\SUMB[29][38] ) );
  FA1A S4_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA1A S4_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), .CO(
        \CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA1A S4_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), 
        .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FA1A S4_6 ( .A(\ab[29][6] ), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), .CO(
        \CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA1A S4_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), 
        .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA1A S4_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA1A S4_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA1A S4_5 ( .A(\ab[29][5] ), .B(\CARRYB[28][5] ), .CI(\SUMB[28][6] ), .CO(
        \CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA1A S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA1A S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), 
        .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA1A S2_28_12 ( .A(\ab[28][12] ), .B(\CARRYB[27][12] ), .CI(\SUMB[27][13] ), 
        .CO(\CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA1A S2_28_5 ( .A(\ab[28][5] ), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA1A S4_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA1A S4_14 ( .A(\ab[29][14] ), .B(\CARRYB[28][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA1A S4_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), 
        .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA1A S4_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA1A S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), 
        .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA1A S2_27_5 ( .A(\ab[27][5] ), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA1A S4_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), .CO(
        \CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA1A S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA1A S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA1A S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA1A S2_28_14 ( .A(\ab[28][14] ), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA1A S2_28_13 ( .A(\ab[28][13] ), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), 
        .CO(\CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA1A S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA1A S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA1A S2_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA1A S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA1A S2_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\SUMB[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA1A S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA1A S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA1A S2_27_15 ( .A(\ab[27][15] ), .B(\CARRYB[26][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA1A S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA1A S2_27_13 ( .A(\ab[27][13] ), .B(\CARRYB[26][13] ), .CI(\SUMB[26][14] ), 
        .CO(\CARRYB[27][13] ), .S(\SUMB[27][13] ) );
  FA1A S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA1A S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA1A S2_27_11 ( .A(\ab[27][11] ), .B(\CARRYB[26][11] ), .CI(\SUMB[26][12] ), 
        .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FA1A S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA1A S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA1A S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA1A S2_26_18 ( .A(\ab[26][18] ), .B(\CARRYB[25][18] ), .CI(\SUMB[25][19] ), 
        .CO(\CARRYB[26][18] ), .S(\SUMB[26][18] ) );
  FA1A S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA1A S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA1A S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA1A S2_26_14 ( .A(\ab[26][14] ), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), 
        .CO(\CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA1A S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), 
        .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA1A S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA1A S2_26_12 ( .A(\ab[26][12] ), .B(\CARRYB[25][12] ), .CI(\SUMB[25][13] ), 
        .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FA1A S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), 
        .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA1A S2_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA1A S2_26_9 ( .A(\ab[26][9] ), .B(\CARRYB[25][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA1A S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA1A S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA1A S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA1A S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA1A S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA1A S2_25_14 ( .A(\ab[25][14] ), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), 
        .CO(\CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA1A S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA1A S2_25_13 ( .A(\ab[25][13] ), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), 
        .CO(\CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA1A S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), 
        .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA1A S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), 
        .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA1A S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA1A S2_25_9 ( .A(\ab[25][9] ), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA1A S2_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\SUMB[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA1A S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA1A S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA1A S2_24_16 ( .A(\ab[24][16] ), .B(\CARRYB[23][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA1A S2_24_15 ( .A(\ab[24][15] ), .B(\CARRYB[23][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA1A S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA1A S2_24_14 ( .A(\ab[24][14] ), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), 
        .CO(\CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA1A S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), 
        .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA1A S2_24_12 ( .A(\ab[24][12] ), .B(\CARRYB[23][12] ), .CI(\SUMB[23][13] ), 
        .CO(\CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA1A S2_24_11 ( .A(\ab[24][11] ), .B(\CARRYB[23][11] ), .CI(\SUMB[23][12] ), 
        .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA1A S2_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA1A S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA1A S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA1A S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA1A S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA1A S2_23_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA1A S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1A S2_23_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA1A S2_23_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA1A S2_23_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA1A S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA1A S2_23_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA1A S2_23_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA1A S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA1A S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA1A S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA1A S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA1A S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA1A S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA1A S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA1A S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA1A S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA1A S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA1A S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA1A S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA1A S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA1A S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA1A S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA1A S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1A S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA1A S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA1A S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA1A S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA1A S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA1A S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA1A S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA1A S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1A S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1A S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA1A S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1A S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA1A S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA1A S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA1A S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA1A S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA1A S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA1A S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA1A S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA1A S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA1A S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1A S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA1A S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1A S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA1A S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA1A S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA1A S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA1A S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA1A S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA1A S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA1A S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA1A S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA1A S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA1A S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1A S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA1A S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA1A S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA1A S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA1A S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA1A S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA1A S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA1A S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA1A S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA1A S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA1A S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA1A S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1A S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA1A S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA1A S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA1A S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA1A S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA1A S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA1A S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA1A S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA1A S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA1A S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA1A S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1A S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA1A S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA1A S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA1A S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA1A S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA1A S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA1A S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA1A S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA1A S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA1A S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1A S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA1A S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA1A S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA1A S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA1A S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA1A S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA1A S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA1A S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA1A S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA1A S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1A S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA1A S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA1A S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA1A S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA1A S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA1A S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA1A S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA1A S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA1A S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA1A S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA1A S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA1A S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA1A S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1A S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1A S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1A S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1A S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1A S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1A S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1A S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1A S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1A S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1A S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1A S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1A S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA1A S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1A S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1A S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1A S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA1A S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1A S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1A S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1A S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1A S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1A S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1A S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1A S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1A S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1A S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1A S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA1A S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1A S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1A S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1A S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1A S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1A S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1A S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1A S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1A S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1A S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1A S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S4_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA1A S4_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA1A S4_12 ( .A(\ab[29][12] ), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), 
        .CO(\CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA1A S4_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA1A S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA1A S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA1A S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA1A S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA1A S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA1A S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA1A S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA1A S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA1A S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA1A S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA1A S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA1A S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA1A S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA1A S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA1A S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA1A S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA1A S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA1A S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1A S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1A S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1A S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA1A S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1A S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1A S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA1A S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1A S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  AN2P U2 ( .A(n173), .B(n305), .Z(n3) );
  IVDA U3 ( .A(n557), .Z(n4) );
  IVP U4 ( .A(A[22]), .Z(n557) );
  IVP U5 ( .A(n10), .Z(n8) );
  IVP U6 ( .A(n10), .Z(n9) );
  IVP U7 ( .A(n10), .Z(n7) );
  IVP U8 ( .A(n10), .Z(n6) );
  IVP U9 ( .A(n10), .Z(n5) );
  IVP U10 ( .A(n181), .Z(n174) );
  IVP U11 ( .A(n172), .Z(n165) );
  IVP U12 ( .A(n181), .Z(n176) );
  IVP U13 ( .A(n181), .Z(n177) );
  IVP U14 ( .A(n181), .Z(n173) );
  IVP U15 ( .A(n172), .Z(n164) );
  IVP U16 ( .A(n181), .Z(n175) );
  IVP U17 ( .A(n172), .Z(n167) );
  IVP U18 ( .A(n190), .Z(n183) );
  IVP U19 ( .A(n190), .Z(n185) );
  IVP U20 ( .A(n172), .Z(n168) );
  IVP U21 ( .A(n181), .Z(n178) );
  IVP U22 ( .A(n190), .Z(n186) );
  IVP U23 ( .A(n190), .Z(n182) );
  IVP U24 ( .A(n172), .Z(n166) );
  IVP U25 ( .A(n190), .Z(n184) );
  IVP U26 ( .A(n172), .Z(n169) );
  IVP U27 ( .A(n199), .Z(n192) );
  IVP U28 ( .A(n181), .Z(n179) );
  IVP U29 ( .A(n190), .Z(n187) );
  IVP U30 ( .A(n199), .Z(n193) );
  IVP U31 ( .A(n199), .Z(n194) );
  IVP U32 ( .A(n172), .Z(n170) );
  IVP U33 ( .A(n199), .Z(n191) );
  IVP U34 ( .A(n190), .Z(n188) );
  IVP U35 ( .A(n199), .Z(n195) );
  IVP U36 ( .A(n181), .Z(n180) );
  IVP U37 ( .A(n208), .Z(n201) );
  IVP U38 ( .A(n199), .Z(n196) );
  IVP U39 ( .A(n172), .Z(n171) );
  IVP U40 ( .A(n208), .Z(n203) );
  IVP U41 ( .A(n208), .Z(n204) );
  IVP U42 ( .A(n190), .Z(n189) );
  IVP U43 ( .A(n208), .Z(n200) );
  IVP U44 ( .A(n208), .Z(n202) );
  IVP U45 ( .A(n199), .Z(n197) );
  IVP U46 ( .A(n208), .Z(n205) );
  IVP U47 ( .A(n217), .Z(n210) );
  IVP U48 ( .A(n199), .Z(n198) );
  IVP U49 ( .A(n217), .Z(n211) );
  IVP U50 ( .A(n217), .Z(n212) );
  IVP U51 ( .A(n217), .Z(n209) );
  IVP U52 ( .A(n208), .Z(n206) );
  IVP U53 ( .A(n217), .Z(n213) );
  IVP U54 ( .A(n226), .Z(n219) );
  IVP U55 ( .A(n217), .Z(n214) );
  IVP U56 ( .A(n208), .Z(n207) );
  IVP U57 ( .A(n226), .Z(n221) );
  IVP U58 ( .A(n226), .Z(n222) );
  IVP U59 ( .A(n226), .Z(n218) );
  IVP U60 ( .A(n226), .Z(n220) );
  IVP U61 ( .A(n235), .Z(n228) );
  IVP U62 ( .A(n235), .Z(n230) );
  IVP U63 ( .A(n217), .Z(n215) );
  IVP U64 ( .A(n235), .Z(n227) );
  IVP U65 ( .A(n226), .Z(n223) );
  IVP U66 ( .A(n235), .Z(n231) );
  IVP U67 ( .A(n235), .Z(n229) );
  IVP U68 ( .A(n217), .Z(n216) );
  IVP U69 ( .A(n244), .Z(n237) );
  IVP U70 ( .A(n226), .Z(n224) );
  IVP U71 ( .A(n235), .Z(n232) );
  IVP U72 ( .A(n244), .Z(n239) );
  IVP U73 ( .A(n235), .Z(n233) );
  IVP U74 ( .A(n244), .Z(n240) );
  IVP U75 ( .A(n226), .Z(n225) );
  IVP U76 ( .A(n244), .Z(n236) );
  IVP U77 ( .A(n244), .Z(n238) );
  IVP U78 ( .A(n244), .Z(n241) );
  IVP U79 ( .A(n253), .Z(n246) );
  IVP U80 ( .A(n235), .Z(n234) );
  IVP U81 ( .A(n253), .Z(n245) );
  IVP U82 ( .A(n253), .Z(n248) );
  IVP U83 ( .A(n244), .Z(n242) );
  IVP U84 ( .A(n253), .Z(n249) );
  IVP U85 ( .A(n253), .Z(n247) );
  IVP U86 ( .A(n262), .Z(n255) );
  IVP U87 ( .A(n253), .Z(n250) );
  IVP U88 ( .A(n244), .Z(n243) );
  IVP U89 ( .A(n262), .Z(n254) );
  IVP U90 ( .A(n262), .Z(n256) );
  IVP U91 ( .A(n262), .Z(n257) );
  IVP U92 ( .A(n262), .Z(n258) );
  IVP U93 ( .A(n271), .Z(n264) );
  IVP U94 ( .A(n253), .Z(n251) );
  IVP U95 ( .A(n262), .Z(n259) );
  IVP U96 ( .A(n271), .Z(n263) );
  IVP U97 ( .A(n262), .Z(n260) );
  IVP U98 ( .A(n271), .Z(n266) );
  IVP U99 ( .A(n271), .Z(n267) );
  IVP U100 ( .A(n253), .Z(n252) );
  IVP U101 ( .A(n271), .Z(n265) );
  IVP U102 ( .A(n271), .Z(n268) );
  IVP U103 ( .A(n280), .Z(n273) );
  IVP U104 ( .A(n262), .Z(n261) );
  IVP U105 ( .A(n280), .Z(n274) );
  IVP U106 ( .A(n280), .Z(n275) );
  IVP U107 ( .A(n280), .Z(n276) );
  IVP U108 ( .A(n271), .Z(n269) );
  IVP U109 ( .A(n280), .Z(n272) );
  IVP U110 ( .A(n289), .Z(n282) );
  IVP U111 ( .A(n289), .Z(n281) );
  IVP U112 ( .A(n280), .Z(n277) );
  IVP U113 ( .A(n289), .Z(n285) );
  IVP U114 ( .A(n271), .Z(n270) );
  IVP U115 ( .A(n289), .Z(n283) );
  IVP U116 ( .A(n289), .Z(n284) );
  IVP U117 ( .A(n289), .Z(n286) );
  IVP U118 ( .A(n280), .Z(n278) );
  IVP U119 ( .A(n298), .Z(n291) );
  IVP U120 ( .A(n298), .Z(n293) );
  IVP U121 ( .A(n298), .Z(n294) );
  IVP U122 ( .A(n289), .Z(n287) );
  IVP U123 ( .A(n280), .Z(n279) );
  IVP U124 ( .A(n298), .Z(n290) );
  IVP U125 ( .A(n298), .Z(n292) );
  IVP U126 ( .A(n549), .Z(n10) );
  IVP U127 ( .A(n298), .Z(n295) );
  IVP U128 ( .A(n289), .Z(n288) );
  IVP U129 ( .A(n549), .Z(n13) );
  IVP U130 ( .A(n298), .Z(n296) );
  IVP U131 ( .A(n549), .Z(n12) );
  IVP U132 ( .A(n549), .Z(n14) );
  IVP U133 ( .A(n549), .Z(n15) );
  IVP U134 ( .A(n158), .Z(n156) );
  IVP U135 ( .A(n549), .Z(n11) );
  IVP U136 ( .A(n298), .Z(n297) );
  IVP U137 ( .A(n158), .Z(n157) );
  IVP U138 ( .A(n158), .Z(n155) );
  IVP U139 ( .A(n158), .Z(n154) );
  IVP U140 ( .A(n147), .Z(n145) );
  IVP U141 ( .A(n147), .Z(n146) );
  IVP U142 ( .A(n147), .Z(n144) );
  IVP U143 ( .A(n136), .Z(n134) );
  IVP U144 ( .A(n158), .Z(n153) );
  IVP U145 ( .A(n136), .Z(n135) );
  IVP U146 ( .A(n147), .Z(n143) );
  IVP U147 ( .A(n136), .Z(n133) );
  IVP U148 ( .A(n125), .Z(n123) );
  IVP U149 ( .A(n136), .Z(n132) );
  IVP U150 ( .A(n147), .Z(n142) );
  IVP U151 ( .A(n125), .Z(n124) );
  IVP U152 ( .A(n125), .Z(n122) );
  IVP U153 ( .A(n125), .Z(n121) );
  IVP U154 ( .A(n114), .Z(n112) );
  IVP U155 ( .A(n136), .Z(n131) );
  IVP U156 ( .A(n114), .Z(n113) );
  IVP U157 ( .A(n114), .Z(n111) );
  IVP U158 ( .A(n125), .Z(n120) );
  IVP U159 ( .A(n103), .Z(n101) );
  IVP U160 ( .A(n114), .Z(n110) );
  IVP U161 ( .A(n103), .Z(n102) );
  IVP U162 ( .A(n103), .Z(n100) );
  IVP U163 ( .A(n114), .Z(n109) );
  IVP U164 ( .A(n103), .Z(n99) );
  IVP U165 ( .A(n103), .Z(n98) );
  IVP U166 ( .A(n87), .Z(n85) );
  IVP U167 ( .A(n87), .Z(n86) );
  IVP U168 ( .A(n87), .Z(n84) );
  IVP U169 ( .A(n76), .Z(n74) );
  IVP U170 ( .A(n76), .Z(n75) );
  IVP U171 ( .A(n87), .Z(n83) );
  IVP U172 ( .A(n76), .Z(n73) );
  IVP U173 ( .A(n65), .Z(n63) );
  IVP U174 ( .A(n87), .Z(n82) );
  IVP U175 ( .A(n76), .Z(n72) );
  IVP U176 ( .A(n65), .Z(n64) );
  IVP U177 ( .A(n65), .Z(n62) );
  IVP U178 ( .A(n54), .Z(n52) );
  IVP U179 ( .A(n65), .Z(n61) );
  IVP U180 ( .A(n76), .Z(n71) );
  IVP U181 ( .A(n54), .Z(n53) );
  IVP U182 ( .A(n54), .Z(n51) );
  IVP U183 ( .A(n65), .Z(n60) );
  IVP U184 ( .A(n43), .Z(n41) );
  IVP U185 ( .A(n54), .Z(n50) );
  IVP U186 ( .A(n43), .Z(n42) );
  IVP U187 ( .A(n43), .Z(n40) );
  IVP U188 ( .A(n32), .Z(n30) );
  IVP U189 ( .A(n54), .Z(n49) );
  IVP U190 ( .A(n32), .Z(n31) );
  IVP U191 ( .A(n32), .Z(n29) );
  IVP U192 ( .A(n43), .Z(n39) );
  IVP U193 ( .A(n21), .Z(n19) );
  IVP U194 ( .A(n43), .Z(n38) );
  IVP U195 ( .A(n32), .Z(n28) );
  IVP U196 ( .A(n21), .Z(n20) );
  IVP U197 ( .A(n21), .Z(n18) );
  IVP U198 ( .A(n32), .Z(n27) );
  IVP U199 ( .A(n21), .Z(n17) );
  IVP U200 ( .A(n21), .Z(n16) );
  IVP U201 ( .A(A[1]), .Z(n181) );
  IVP U202 ( .A(A[0]), .Z(n172) );
  IVP U203 ( .A(A[2]), .Z(n190) );
  IVP U204 ( .A(A[3]), .Z(n199) );
  IVP U205 ( .A(A[4]), .Z(n208) );
  IVP U206 ( .A(A[5]), .Z(n217) );
  IVP U207 ( .A(A[6]), .Z(n226) );
  IVP U208 ( .A(A[7]), .Z(n235) );
  IVP U209 ( .A(A[8]), .Z(n244) );
  IVP U210 ( .A(A[9]), .Z(n253) );
  IVP U211 ( .A(A[10]), .Z(n262) );
  IVP U212 ( .A(A[11]), .Z(n271) );
  IVP U213 ( .A(A[12]), .Z(n280) );
  IVP U214 ( .A(A[13]), .Z(n289) );
  IVP U215 ( .A(A[14]), .Z(n298) );
  IVP U216 ( .A(A[15]), .Z(n549) );
  IVP U217 ( .A(n563), .Z(n158) );
  IVP U218 ( .A(n563), .Z(n161) );
  IVP U219 ( .A(n563), .Z(n162) );
  IVP U220 ( .A(n563), .Z(n160) );
  IVP U221 ( .A(n563), .Z(n159) );
  IVP U222 ( .A(n563), .Z(n163) );
  IVP U223 ( .A(n562), .Z(n147) );
  IVP U224 ( .A(n562), .Z(n150) );
  IVP U225 ( .A(n562), .Z(n151) );
  IVP U226 ( .A(n562), .Z(n149) );
  IVP U227 ( .A(n562), .Z(n148) );
  IVP U228 ( .A(n562), .Z(n152) );
  IVP U229 ( .A(n561), .Z(n136) );
  IVP U230 ( .A(n561), .Z(n139) );
  IVP U231 ( .A(n561), .Z(n140) );
  IVP U232 ( .A(n561), .Z(n138) );
  IVP U233 ( .A(n561), .Z(n137) );
  IVP U234 ( .A(n561), .Z(n141) );
  IVP U235 ( .A(n560), .Z(n125) );
  IVP U236 ( .A(n560), .Z(n129) );
  IVP U237 ( .A(n560), .Z(n128) );
  IVP U238 ( .A(n560), .Z(n127) );
  IVP U239 ( .A(n560), .Z(n126) );
  IVP U240 ( .A(n560), .Z(n130) );
  IVP U241 ( .A(n559), .Z(n114) );
  IVP U242 ( .A(n559), .Z(n118) );
  IVP U243 ( .A(n559), .Z(n117) );
  IVP U244 ( .A(n559), .Z(n116) );
  IVP U245 ( .A(n559), .Z(n115) );
  IVP U246 ( .A(n559), .Z(n119) );
  IVP U247 ( .A(n558), .Z(n103) );
  IVP U248 ( .A(n558), .Z(n107) );
  IVP U249 ( .A(n558), .Z(n106) );
  IVP U250 ( .A(n558), .Z(n105) );
  IVP U251 ( .A(n558), .Z(n104) );
  IVP U252 ( .A(n557), .Z(n96) );
  IVP U253 ( .A(n557), .Z(n95) );
  IVP U254 ( .A(n558), .Z(n108) );
  IVP U255 ( .A(n557), .Z(n94) );
  IVP U256 ( .A(n557), .Z(n93) );
  IVP U257 ( .A(n557), .Z(n97) );
  IVP U258 ( .A(n556), .Z(n87) );
  IVP U259 ( .A(n556), .Z(n91) );
  IVP U260 ( .A(n556), .Z(n90) );
  IVP U261 ( .A(n556), .Z(n89) );
  IVP U262 ( .A(n556), .Z(n88) );
  IVP U263 ( .A(n556), .Z(n92) );
  IVP U264 ( .A(n555), .Z(n76) );
  IVP U265 ( .A(n555), .Z(n80) );
  IVP U266 ( .A(n555), .Z(n79) );
  IVP U267 ( .A(n555), .Z(n78) );
  IVP U268 ( .A(n555), .Z(n77) );
  IVP U269 ( .A(n555), .Z(n81) );
  IVP U270 ( .A(n554), .Z(n65) );
  IVP U271 ( .A(n554), .Z(n68) );
  IVP U272 ( .A(n554), .Z(n69) );
  IVP U273 ( .A(n554), .Z(n70) );
  IVP U274 ( .A(n554), .Z(n67) );
  IVP U275 ( .A(n554), .Z(n66) );
  IVP U276 ( .A(n553), .Z(n54) );
  IVP U277 ( .A(n553), .Z(n57) );
  IVP U278 ( .A(n553), .Z(n56) );
  IVP U279 ( .A(n553), .Z(n58) );
  IVP U280 ( .A(n553), .Z(n59) );
  IVP U281 ( .A(n553), .Z(n55) );
  IVP U282 ( .A(n552), .Z(n43) );
  IVP U283 ( .A(n552), .Z(n47) );
  IVP U284 ( .A(n552), .Z(n46) );
  IVP U285 ( .A(n552), .Z(n45) );
  IVP U286 ( .A(n552), .Z(n44) );
  IVP U287 ( .A(n552), .Z(n48) );
  IVP U288 ( .A(n551), .Z(n32) );
  IVP U289 ( .A(n551), .Z(n36) );
  IVP U290 ( .A(n551), .Z(n35) );
  IVP U291 ( .A(n551), .Z(n34) );
  IVP U292 ( .A(n551), .Z(n33) );
  IVP U293 ( .A(n551), .Z(n37) );
  IVP U294 ( .A(n550), .Z(n21) );
  IVP U295 ( .A(n550), .Z(n24) );
  IVP U296 ( .A(n550), .Z(n25) );
  IVP U297 ( .A(n550), .Z(n23) );
  IVP U298 ( .A(n550), .Z(n22) );
  IVP U299 ( .A(n550), .Z(n26) );
  EO U300 ( .A(\CARRYB[29][19] ), .B(\SUMB[29][20] ), .Z(\A1[47] ) );
  EO U301 ( .A(\CARRYB[29][10] ), .B(\SUMB[29][11] ), .Z(\A1[38] ) );
  EO U302 ( .A(\CARRYB[29][15] ), .B(\SUMB[29][16] ), .Z(\A1[43] ) );
  EO U303 ( .A(\CARRYB[29][14] ), .B(\SUMB[29][15] ), .Z(\A1[42] ) );
  EO U304 ( .A(\CARRYB[29][5] ), .B(\SUMB[29][6] ), .Z(\A1[33] ) );
  EO U305 ( .A(\CARRYB[29][13] ), .B(\SUMB[29][14] ), .Z(\A1[41] ) );
  EO U306 ( .A(\CARRYB[29][9] ), .B(\SUMB[29][10] ), .Z(\A1[37] ) );
  EO U307 ( .A(\CARRYB[29][17] ), .B(\SUMB[29][18] ), .Z(\A1[45] ) );
  EO U308 ( .A(\CARRYB[29][18] ), .B(\SUMB[29][19] ), .Z(\A1[46] ) );
  EO U309 ( .A(\CARRYB[29][11] ), .B(\SUMB[29][12] ), .Z(\A1[39] ) );
  EO U310 ( .A(\CARRYB[29][16] ), .B(\SUMB[29][17] ), .Z(\A1[44] ) );
  EO U311 ( .A(\CARRYB[29][22] ), .B(\SUMB[29][23] ), .Z(\A1[50] ) );
  EO U312 ( .A(\CARRYB[29][23] ), .B(\SUMB[29][24] ), .Z(\A1[51] ) );
  EO U313 ( .A(\CARRYB[29][7] ), .B(\SUMB[29][8] ), .Z(\A1[35] ) );
  EO U314 ( .A(\CARRYB[29][25] ), .B(\SUMB[29][26] ), .Z(\A1[53] ) );
  EO U315 ( .A(\CARRYB[29][6] ), .B(\SUMB[29][7] ), .Z(\A1[34] ) );
  EO U316 ( .A(\CARRYB[29][21] ), .B(\SUMB[29][22] ), .Z(\A1[49] ) );
  EO U317 ( .A(\CARRYB[29][27] ), .B(\SUMB[29][28] ), .Z(\A1[55] ) );
  EO U318 ( .A(\CARRYB[29][26] ), .B(\SUMB[29][27] ), .Z(\A1[54] ) );
  EO U319 ( .A(\CARRYB[29][2] ), .B(\SUMB[29][3] ), .Z(\A1[30] ) );
  EO U320 ( .A(\CARRYB[29][37] ), .B(\SUMB[29][38] ), .Z(\A1[65] ) );
  EO U321 ( .A(\CARRYB[29][31] ), .B(\SUMB[29][32] ), .Z(\A1[59] ) );
  EO U322 ( .A(\CARRYB[29][34] ), .B(\SUMB[29][35] ), .Z(\A1[62] ) );
  EO U323 ( .A(\CARRYB[29][33] ), .B(\SUMB[29][34] ), .Z(\A1[61] ) );
  EO U324 ( .A(\CARRYB[29][35] ), .B(\SUMB[29][36] ), .Z(\A1[63] ) );
  EO U325 ( .A(\CARRYB[29][8] ), .B(\SUMB[29][9] ), .Z(\A1[36] ) );
  EO U326 ( .A(\CARRYB[29][4] ), .B(\SUMB[29][5] ), .Z(\A1[32] ) );
  EO U327 ( .A(\CARRYB[29][24] ), .B(\SUMB[29][25] ), .Z(\A1[52] ) );
  EO U328 ( .A(\CARRYB[29][12] ), .B(\SUMB[29][13] ), .Z(\A1[40] ) );
  EO U329 ( .A(\CARRYB[29][29] ), .B(\SUMB[29][30] ), .Z(\A1[57] ) );
  EO U330 ( .A(\CARRYB[29][30] ), .B(\SUMB[29][31] ), .Z(\A1[58] ) );
  EO U331 ( .A(\CARRYB[29][20] ), .B(\SUMB[29][21] ), .Z(\A1[48] ) );
  EO U332 ( .A(\CARRYB[29][3] ), .B(\SUMB[29][4] ), .Z(\A1[31] ) );
  EO U333 ( .A(\CARRYB[29][28] ), .B(\SUMB[29][29] ), .Z(\A1[56] ) );
  EO U334 ( .A(\CARRYB[29][36] ), .B(\SUMB[29][37] ), .Z(\A1[64] ) );
  EO U335 ( .A(\CARRYB[29][32] ), .B(\SUMB[29][33] ), .Z(\A1[60] ) );
  EO U336 ( .A(\CARRYB[29][1] ), .B(\SUMB[29][2] ), .Z(\A1[29] ) );
  EO U337 ( .A(\ab[0][2] ), .B(n3), .Z(\SUMB[1][1] ) );
  IVP U338 ( .A(A[16]), .Z(n563) );
  IVP U339 ( .A(A[17]), .Z(n562) );
  IVP U340 ( .A(A[18]), .Z(n561) );
  IVP U341 ( .A(A[19]), .Z(n560) );
  IVP U342 ( .A(A[20]), .Z(n559) );
  IVP U343 ( .A(A[21]), .Z(n558) );
  IVP U344 ( .A(A[23]), .Z(n556) );
  IVP U345 ( .A(A[24]), .Z(n555) );
  IVP U346 ( .A(A[25]), .Z(n554) );
  IVP U347 ( .A(A[26]), .Z(n553) );
  IVP U348 ( .A(A[27]), .Z(n552) );
  IVP U349 ( .A(A[28]), .Z(n551) );
  IVP U350 ( .A(A[29]), .Z(n550) );
  EO U351 ( .A(\CARRYB[29][0] ), .B(\SUMB[29][1] ), .Z(\A1[28] ) );
  EO U352 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Z(\SUMB[1][20] ) );
  EO U353 ( .A(\CARRYB[29][46] ), .B(\SUMB[29][47] ), .Z(\A1[74] ) );
  EO U354 ( .A(\CARRYB[29][50] ), .B(\SUMB[29][51] ), .Z(\A1[78] ) );
  EO U355 ( .A(\CARRYB[29][49] ), .B(\SUMB[29][50] ), .Z(\A1[77] ) );
  EO U356 ( .A(\CARRYB[29][45] ), .B(\SUMB[29][46] ), .Z(\A1[73] ) );
  EO U357 ( .A(\CARRYB[29][47] ), .B(\SUMB[29][48] ), .Z(\A1[75] ) );
  EO U358 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U359 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U360 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U361 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U362 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U363 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U364 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Z(\SUMB[1][16] ) );
  EO U365 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Z(\SUMB[1][17] ) );
  EO U366 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Z(\SUMB[1][18] ) );
  EO U367 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Z(\SUMB[1][19] ) );
  EO U368 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Z(\SUMB[1][21] ) );
  EO U369 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U370 ( .A(\CARRYB[29][39] ), .B(\SUMB[29][40] ), .Z(\A1[67] ) );
  EO U371 ( .A(\CARRYB[29][41] ), .B(\SUMB[29][42] ), .Z(\A1[69] ) );
  EO U372 ( .A(\CARRYB[29][42] ), .B(\SUMB[29][43] ), .Z(\A1[70] ) );
  EO U373 ( .A(\CARRYB[29][62] ), .B(\SUMB[29][63] ), .Z(\A1[90] ) );
  EO U374 ( .A(\CARRYB[29][61] ), .B(\SUMB[29][62] ), .Z(\A1[89] ) );
  EO U375 ( .A(\CARRYB[29][40] ), .B(\SUMB[29][41] ), .Z(\A1[68] ) );
  EO U376 ( .A(\CARRYB[29][51] ), .B(\SUMB[29][52] ), .Z(\A1[79] ) );
  EO U377 ( .A(\CARRYB[29][38] ), .B(\SUMB[29][39] ), .Z(\A1[66] ) );
  EO U378 ( .A(\CARRYB[29][43] ), .B(\SUMB[29][44] ), .Z(\A1[71] ) );
  EO U379 ( .A(\CARRYB[29][44] ), .B(\SUMB[29][45] ), .Z(\A1[72] ) );
  EO U380 ( .A(\CARRYB[29][48] ), .B(\SUMB[29][49] ), .Z(\A1[76] ) );
  EO U381 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Z(\SUMB[1][22] ) );
  EO U382 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Z(\SUMB[1][23] ) );
  EO U383 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Z(\SUMB[1][24] ) );
  EO U384 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Z(\SUMB[1][25] ) );
  EO U385 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Z(\SUMB[1][26] ) );
  EO U386 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Z(\SUMB[1][27] ) );
  EO U387 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Z(\SUMB[1][28] ) );
  EO U388 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Z(\SUMB[1][29] ) );
  EO U389 ( .A(\ab[0][33] ), .B(\ab[1][32] ), .Z(\SUMB[1][32] ) );
  EO U390 ( .A(\ab[0][34] ), .B(\ab[1][33] ), .Z(\SUMB[1][33] ) );
  EO U391 ( .A(\ab[0][35] ), .B(\ab[1][34] ), .Z(\SUMB[1][34] ) );
  EO U392 ( .A(\ab[0][36] ), .B(\ab[1][35] ), .Z(\SUMB[1][35] ) );
  EO U393 ( .A(\ab[0][37] ), .B(\ab[1][36] ), .Z(\SUMB[1][36] ) );
  EO U394 ( .A(\ab[0][38] ), .B(\ab[1][37] ), .Z(\SUMB[1][37] ) );
  EO U395 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U396 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U397 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U398 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U399 ( .A(\ab[0][63] ), .B(\ab[1][62] ), .Z(\SUMB[1][62] ) );
  EO U400 ( .A(\ab[0][64] ), .B(\ab[1][63] ), .Z(\SUMB[1][63] ) );
  EO U401 ( .A(\ab[0][65] ), .B(\ab[1][64] ), .Z(\SUMB[1][64] ) );
  EO U402 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U403 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U404 ( .A(\CARRYB[29][59] ), .B(\SUMB[29][60] ), .Z(\A1[87] ) );
  EO U405 ( .A(\CARRYB[29][66] ), .B(\SUMB[29][67] ), .Z(\A1[94] ) );
  EO U406 ( .A(\CARRYB[29][67] ), .B(\SUMB[29][68] ), .Z(\A1[95] ) );
  EO U407 ( .A(\CARRYB[29][65] ), .B(\SUMB[29][66] ), .Z(\A1[93] ) );
  EO U408 ( .A(\CARRYB[29][64] ), .B(\SUMB[29][65] ), .Z(\A1[92] ) );
  EO U409 ( .A(\CARRYB[29][63] ), .B(\SUMB[29][64] ), .Z(\A1[91] ) );
  EO U410 ( .A(\CARRYB[29][60] ), .B(\SUMB[29][61] ), .Z(\A1[88] ) );
  EO U411 ( .A(\CARRYB[29][53] ), .B(\SUMB[29][54] ), .Z(\A1[81] ) );
  EO U412 ( .A(\CARRYB[29][55] ), .B(\SUMB[29][56] ), .Z(\A1[83] ) );
  EO U413 ( .A(\CARRYB[29][58] ), .B(\SUMB[29][59] ), .Z(\A1[86] ) );
  EO U414 ( .A(\CARRYB[29][54] ), .B(\SUMB[29][55] ), .Z(\A1[82] ) );
  EO U415 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Z(\SUMB[1][30] ) );
  EO U416 ( .A(\ab[0][32] ), .B(\ab[1][31] ), .Z(\SUMB[1][31] ) );
  EO U417 ( .A(\ab[0][62] ), .B(\ab[1][61] ), .Z(\SUMB[1][61] ) );
  EO U418 ( .A(\ab[0][66] ), .B(\ab[1][65] ), .Z(\SUMB[1][65] ) );
  EO U419 ( .A(\ab[0][67] ), .B(\ab[1][66] ), .Z(\SUMB[1][66] ) );
  EO U420 ( .A(\ab[0][68] ), .B(\ab[1][67] ), .Z(\SUMB[1][67] ) );
  EO U421 ( .A(\ab[0][69] ), .B(\ab[1][68] ), .Z(\SUMB[1][68] ) );
  EO U422 ( .A(\ab[0][70] ), .B(\ab[1][69] ), .Z(\SUMB[1][69] ) );
  EO U423 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U424 ( .A(\CARRYB[29][71] ), .B(\SUMB[29][72] ), .Z(\A1[99] ) );
  EO U425 ( .A(\CARRYB[29][56] ), .B(\SUMB[29][57] ), .Z(\A1[84] ) );
  EO U426 ( .A(\CARRYB[29][69] ), .B(\SUMB[29][70] ), .Z(\A1[97] ) );
  EO U427 ( .A(\CARRYB[29][70] ), .B(\SUMB[29][71] ), .Z(\A1[98] ) );
  EO U428 ( .A(\CARRYB[29][75] ), .B(\SUMB[29][76] ), .Z(\A1[103] ) );
  EO U429 ( .A(\CARRYB[29][77] ), .B(\SUMB[29][78] ), .Z(\A1[105] ) );
  EO U430 ( .A(\CARRYB[29][78] ), .B(\SUMB[29][79] ), .Z(\A1[106] ) );
  EO U431 ( .A(\CARRYB[29][73] ), .B(\SUMB[29][74] ), .Z(\A1[101] ) );
  EO U432 ( .A(\CARRYB[29][74] ), .B(\SUMB[29][75] ), .Z(\A1[102] ) );
  EO U433 ( .A(\CARRYB[29][52] ), .B(\SUMB[29][53] ), .Z(\A1[80] ) );
  EO U434 ( .A(\CARRYB[29][68] ), .B(\SUMB[29][69] ), .Z(\A1[96] ) );
  EO U435 ( .A(\CARRYB[29][72] ), .B(\SUMB[29][73] ), .Z(\A1[100] ) );
  EO U436 ( .A(\CARRYB[29][57] ), .B(\SUMB[29][58] ), .Z(\A1[85] ) );
  EO U437 ( .A(\ab[0][71] ), .B(\ab[1][70] ), .Z(\SUMB[1][70] ) );
  EO U438 ( .A(\ab[0][72] ), .B(\ab[1][71] ), .Z(\SUMB[1][71] ) );
  EO U439 ( .A(\ab[0][73] ), .B(\ab[1][72] ), .Z(\SUMB[1][72] ) );
  EO U440 ( .A(\ab[0][74] ), .B(\ab[1][73] ), .Z(\SUMB[1][73] ) );
  EO U441 ( .A(\ab[0][75] ), .B(\ab[1][74] ), .Z(\SUMB[1][74] ) );
  EO U442 ( .A(\ab[0][76] ), .B(\ab[1][75] ), .Z(\SUMB[1][75] ) );
  EO U443 ( .A(\ab[0][77] ), .B(\ab[1][76] ), .Z(\SUMB[1][76] ) );
  EO U444 ( .A(\ab[0][78] ), .B(\ab[1][77] ), .Z(\SUMB[1][77] ) );
  EO U445 ( .A(\ab[0][79] ), .B(\ab[1][78] ), .Z(\SUMB[1][78] ) );
  EO U446 ( .A(\ab[0][80] ), .B(\ab[1][79] ), .Z(\SUMB[1][79] ) );
  EO U447 ( .A(\ab[0][81] ), .B(\ab[1][80] ), .Z(\SUMB[1][80] ) );
  EO U448 ( .A(\CARRYB[29][83] ), .B(\SUMB[29][84] ), .Z(\A1[111] ) );
  EO U449 ( .A(\CARRYB[29][76] ), .B(\SUMB[29][77] ), .Z(\A1[104] ) );
  EO U450 ( .A(\CARRYB[29][82] ), .B(\SUMB[29][83] ), .Z(\A1[110] ) );
  EO U451 ( .A(\ab[0][82] ), .B(\ab[1][81] ), .Z(\SUMB[1][81] ) );
  EO U452 ( .A(\ab[0][84] ), .B(\ab[1][83] ), .Z(\SUMB[1][83] ) );
  EO U453 ( .A(\ab[0][85] ), .B(\ab[1][84] ), .Z(\SUMB[1][84] ) );
  EO U454 ( .A(\ab[0][86] ), .B(\ab[1][85] ), .Z(\SUMB[1][85] ) );
  EO U455 ( .A(\CARRYB[29][81] ), .B(\SUMB[29][82] ), .Z(\A1[109] ) );
  EO U456 ( .A(\CARRYB[29][79] ), .B(\SUMB[29][80] ), .Z(\A1[107] ) );
  EO U457 ( .A(\CARRYB[29][80] ), .B(\SUMB[29][81] ), .Z(\A1[108] ) );
  EO U458 ( .A(\ab[0][83] ), .B(\ab[1][82] ), .Z(\SUMB[1][82] ) );
  EO U459 ( .A(\ab[0][87] ), .B(\ab[1][86] ), .Z(\SUMB[1][86] ) );
  EO U460 ( .A(\ab[0][88] ), .B(\ab[1][87] ), .Z(\SUMB[1][87] ) );
  EO U461 ( .A(\CARRYB[29][84] ), .B(\SUMB[29][85] ), .Z(\A1[112] ) );
  EO U462 ( .A(\ab[0][89] ), .B(\ab[1][88] ), .Z(\SUMB[1][88] ) );
  EO U463 ( .A(\CARRYB[29][85] ), .B(\SUMB[29][86] ), .Z(\A1[113] ) );
  EO U464 ( .A(\ab[0][90] ), .B(\ab[1][89] ), .Z(\SUMB[1][89] ) );
  EO U465 ( .A(\CARRYB[29][86] ), .B(\SUMB[29][87] ), .Z(\A1[114] ) );
  EO U466 ( .A(\CARRYB[29][87] ), .B(\SUMB[29][88] ), .Z(\A1[115] ) );
  EO U467 ( .A(\ab[0][91] ), .B(\ab[1][90] ), .Z(\SUMB[1][90] ) );
  EO U468 ( .A(\ab[0][92] ), .B(\ab[1][91] ), .Z(\SUMB[1][91] ) );
  EO U469 ( .A(\CARRYB[29][88] ), .B(\SUMB[29][89] ), .Z(\A1[116] ) );
  EO U470 ( .A(\ab[0][93] ), .B(\ab[1][92] ), .Z(\SUMB[1][92] ) );
  EO U471 ( .A(\ab[0][94] ), .B(\ab[1][93] ), .Z(\SUMB[1][93] ) );
  EO U472 ( .A(\ab[0][95] ), .B(\ab[1][94] ), .Z(\SUMB[1][94] ) );
  EO U473 ( .A(\CARRYB[29][89] ), .B(\SUMB[29][90] ), .Z(\A1[117] ) );
  EO U474 ( .A(\CARRYB[29][90] ), .B(\SUMB[29][91] ), .Z(\A1[118] ) );
  EO U475 ( .A(\CARRYB[29][91] ), .B(\SUMB[29][92] ), .Z(\A1[119] ) );
  EO U476 ( .A(\CARRYB[29][92] ), .B(\SUMB[29][93] ), .Z(\A1[120] ) );
  EO U477 ( .A(\CARRYB[29][93] ), .B(\SUMB[29][94] ), .Z(\A1[121] ) );
  EO U478 ( .A(\CARRYB[29][94] ), .B(\ab[29][95] ), .Z(\A1[122] ) );
  EO U479 ( .A(\ab[0][39] ), .B(\ab[1][38] ), .Z(\SUMB[1][38] ) );
  EO U480 ( .A(\ab[0][40] ), .B(\ab[1][39] ), .Z(\SUMB[1][39] ) );
  EO U481 ( .A(\ab[0][57] ), .B(\ab[1][56] ), .Z(\SUMB[1][56] ) );
  IVP U482 ( .A(n526), .Z(n488) );
  IVP U483 ( .A(n523), .Z(n485) );
  IVP U484 ( .A(n532), .Z(n490) );
  IVP U485 ( .A(n527), .Z(n489) );
  IVP U486 ( .A(n525), .Z(n487) );
  IVP U487 ( .A(n524), .Z(n486) );
  IVP U488 ( .A(n522), .Z(n484) );
  IVP U489 ( .A(n521), .Z(n483) );
  IVP U490 ( .A(n520), .Z(n482) );
  IVP U491 ( .A(n519), .Z(n481) );
  IVP U492 ( .A(n518), .Z(n480) );
  IVP U493 ( .A(n517), .Z(n479) );
  IVP U494 ( .A(n516), .Z(n478) );
  IVP U495 ( .A(n515), .Z(n477) );
  IVP U496 ( .A(n514), .Z(n476) );
  IVP U497 ( .A(n513), .Z(n475) );
  IVP U498 ( .A(n512), .Z(n474) );
  IVP U499 ( .A(n510), .Z(n472) );
  IVP U500 ( .A(n509), .Z(n471) );
  IVP U501 ( .A(n508), .Z(n470) );
  IVP U502 ( .A(n507), .Z(n469) );
  IVP U503 ( .A(n511), .Z(n473) );
  IVP U504 ( .A(n506), .Z(n468) );
  IVP U505 ( .A(n504), .Z(n466) );
  IVP U506 ( .A(n503), .Z(n465) );
  IVP U507 ( .A(n502), .Z(n464) );
  IVP U508 ( .A(n505), .Z(n467) );
  IVP U509 ( .A(n501), .Z(n463) );
  IVP U510 ( .A(n500), .Z(n462) );
  IVP U511 ( .A(n499), .Z(n461) );
  IVP U512 ( .A(n498), .Z(n460) );
  IVP U513 ( .A(n338), .Z(n336) );
  IVP U514 ( .A(n342), .Z(n340) );
  IVP U515 ( .A(n346), .Z(n344) );
  IVP U516 ( .A(n350), .Z(n348) );
  IVP U517 ( .A(n354), .Z(n352) );
  IVP U518 ( .A(n358), .Z(n356) );
  IVP U519 ( .A(n362), .Z(n360) );
  IVP U520 ( .A(n366), .Z(n364) );
  IVP U521 ( .A(n370), .Z(n368) );
  IVP U522 ( .A(n374), .Z(n372) );
  IVP U523 ( .A(n378), .Z(n376) );
  IVP U524 ( .A(n382), .Z(n380) );
  IVP U525 ( .A(n497), .Z(n459) );
  IVP U526 ( .A(n386), .Z(n384) );
  IVP U527 ( .A(n390), .Z(n388) );
  IVP U528 ( .A(n394), .Z(n392) );
  IVP U529 ( .A(n398), .Z(n396) );
  IVP U530 ( .A(n402), .Z(n400) );
  IVP U531 ( .A(n406), .Z(n404) );
  IVP U532 ( .A(n438), .Z(n436) );
  IVP U533 ( .A(n450), .Z(n448) );
  IVP U534 ( .A(n454), .Z(n452) );
  IVP U535 ( .A(n326), .Z(n324) );
  IVP U536 ( .A(n330), .Z(n328) );
  IVP U537 ( .A(n334), .Z(n332) );
  IVP U538 ( .A(n322), .Z(n320) );
  IVP U539 ( .A(n310), .Z(n308) );
  IVP U540 ( .A(n314), .Z(n312) );
  IVP U541 ( .A(n496), .Z(n458) );
  IVP U542 ( .A(n410), .Z(n408) );
  IVP U543 ( .A(n414), .Z(n412) );
  IVP U544 ( .A(n418), .Z(n416) );
  IVP U545 ( .A(n422), .Z(n420) );
  IVP U546 ( .A(n426), .Z(n424) );
  IVP U547 ( .A(n430), .Z(n428) );
  IVP U548 ( .A(n434), .Z(n432) );
  IVP U549 ( .A(n442), .Z(n440) );
  IVP U550 ( .A(n446), .Z(n444) );
  IVP U551 ( .A(n318), .Z(n316) );
  IVP U552 ( .A(n306), .Z(n304) );
  IVP U553 ( .A(n495), .Z(n457) );
  IVP U554 ( .A(n302), .Z(n300) );
  IVP U555 ( .A(n494), .Z(n456) );
  IVP U556 ( .A(n493), .Z(n455) );
  IVP U557 ( .A(n492), .Z(n491) );
  IVP U558 ( .A(n338), .Z(n335) );
  IVP U559 ( .A(n342), .Z(n339) );
  IVP U560 ( .A(n346), .Z(n343) );
  IVP U561 ( .A(n350), .Z(n347) );
  IVP U562 ( .A(n354), .Z(n351) );
  IVP U563 ( .A(n358), .Z(n355) );
  IVP U564 ( .A(n362), .Z(n359) );
  IVP U565 ( .A(n366), .Z(n363) );
  IVP U566 ( .A(n370), .Z(n367) );
  IVP U567 ( .A(n374), .Z(n371) );
  IVP U568 ( .A(n378), .Z(n375) );
  IVP U569 ( .A(n382), .Z(n379) );
  IVP U570 ( .A(n386), .Z(n383) );
  IVP U571 ( .A(n390), .Z(n387) );
  IVP U572 ( .A(n394), .Z(n391) );
  IVP U573 ( .A(n398), .Z(n395) );
  IVP U574 ( .A(n402), .Z(n399) );
  IVP U575 ( .A(n406), .Z(n403) );
  IVP U576 ( .A(n438), .Z(n435) );
  IVP U577 ( .A(n326), .Z(n323) );
  IVP U578 ( .A(n330), .Z(n327) );
  IVP U579 ( .A(n334), .Z(n331) );
  IVP U580 ( .A(n322), .Z(n319) );
  IVP U581 ( .A(n454), .Z(n451) );
  IVP U582 ( .A(n310), .Z(n307) );
  IVP U583 ( .A(n314), .Z(n311) );
  IVP U584 ( .A(n450), .Z(n447) );
  IVP U585 ( .A(n410), .Z(n407) );
  IVP U586 ( .A(n414), .Z(n411) );
  IVP U587 ( .A(n418), .Z(n415) );
  IVP U588 ( .A(n422), .Z(n419) );
  IVP U589 ( .A(n426), .Z(n423) );
  IVP U590 ( .A(n430), .Z(n427) );
  IVP U591 ( .A(n434), .Z(n431) );
  IVP U592 ( .A(n446), .Z(n443) );
  IVP U593 ( .A(n318), .Z(n315) );
  IVP U594 ( .A(n442), .Z(n439) );
  IVP U595 ( .A(n306), .Z(n303) );
  IVP U596 ( .A(n302), .Z(n299) );
  EO U597 ( .A(\ab[0][47] ), .B(\ab[1][46] ), .Z(\SUMB[1][46] ) );
  EO U598 ( .A(\ab[0][48] ), .B(\ab[1][47] ), .Z(\SUMB[1][47] ) );
  EO U599 ( .A(\ab[0][49] ), .B(\ab[1][48] ), .Z(\SUMB[1][48] ) );
  EO U600 ( .A(\ab[0][50] ), .B(\ab[1][49] ), .Z(\SUMB[1][49] ) );
  EO U601 ( .A(\ab[0][51] ), .B(\ab[1][50] ), .Z(\SUMB[1][50] ) );
  EO U602 ( .A(\ab[0][52] ), .B(\ab[1][51] ), .Z(\SUMB[1][51] ) );
  EO U603 ( .A(\ab[0][53] ), .B(\ab[1][52] ), .Z(\SUMB[1][52] ) );
  EO U604 ( .A(\ab[0][41] ), .B(\ab[1][40] ), .Z(\SUMB[1][40] ) );
  EO U605 ( .A(\ab[0][42] ), .B(\ab[1][41] ), .Z(\SUMB[1][41] ) );
  EO U606 ( .A(\ab[0][43] ), .B(\ab[1][42] ), .Z(\SUMB[1][42] ) );
  EO U607 ( .A(\ab[0][44] ), .B(\ab[1][43] ), .Z(\SUMB[1][43] ) );
  EO U608 ( .A(\ab[0][45] ), .B(\ab[1][44] ), .Z(\SUMB[1][44] ) );
  EO U609 ( .A(\ab[0][46] ), .B(\ab[1][45] ), .Z(\SUMB[1][45] ) );
  EO U610 ( .A(\ab[0][54] ), .B(\ab[1][53] ), .Z(\SUMB[1][53] ) );
  EO U611 ( .A(\ab[0][55] ), .B(\ab[1][54] ), .Z(\SUMB[1][54] ) );
  EO U612 ( .A(\ab[0][56] ), .B(\ab[1][55] ), .Z(\SUMB[1][55] ) );
  EO U613 ( .A(\ab[0][58] ), .B(\ab[1][57] ), .Z(\SUMB[1][57] ) );
  EO U614 ( .A(\ab[0][60] ), .B(\ab[1][59] ), .Z(\SUMB[1][59] ) );
  EO U615 ( .A(\ab[0][61] ), .B(\ab[1][60] ), .Z(\SUMB[1][60] ) );
  EO U616 ( .A(\ab[0][59] ), .B(\ab[1][58] ), .Z(\SUMB[1][58] ) );
  IVP U617 ( .A(B[61]), .Z(n526) );
  IVP U618 ( .A(B[64]), .Z(n523) );
  IVP U619 ( .A(B[55]), .Z(n532) );
  IVP U620 ( .A(B[60]), .Z(n527) );
  IVP U621 ( .A(B[62]), .Z(n525) );
  IVP U622 ( .A(B[63]), .Z(n524) );
  IVP U623 ( .A(B[65]), .Z(n522) );
  IVP U624 ( .A(B[66]), .Z(n521) );
  IVP U625 ( .A(B[67]), .Z(n520) );
  IVP U626 ( .A(B[68]), .Z(n519) );
  IVP U627 ( .A(B[69]), .Z(n518) );
  IVP U628 ( .A(B[70]), .Z(n517) );
  IVP U629 ( .A(B[71]), .Z(n516) );
  IVP U630 ( .A(B[73]), .Z(n514) );
  IVP U631 ( .A(B[74]), .Z(n513) );
  IVP U632 ( .A(B[75]), .Z(n512) );
  IVP U633 ( .A(B[77]), .Z(n510) );
  IVP U634 ( .A(B[78]), .Z(n509) );
  IVP U635 ( .A(B[79]), .Z(n508) );
  IVP U636 ( .A(B[80]), .Z(n507) );
  IVP U637 ( .A(B[76]), .Z(n511) );
  IVP U638 ( .A(B[81]), .Z(n506) );
  IVP U639 ( .A(B[83]), .Z(n504) );
  IVP U640 ( .A(B[84]), .Z(n503) );
  IVP U641 ( .A(B[85]), .Z(n502) );
  IVP U642 ( .A(B[82]), .Z(n505) );
  IVP U643 ( .A(B[86]), .Z(n501) );
  IVP U644 ( .A(B[87]), .Z(n500) );
  IVP U645 ( .A(B[88]), .Z(n499) );
  IVP U646 ( .A(B[89]), .Z(n498) );
  IVP U647 ( .A(B[90]), .Z(n497) );
  IVP U648 ( .A(B[91]), .Z(n496) );
  IVP U649 ( .A(B[92]), .Z(n495) );
  IVP U650 ( .A(B[93]), .Z(n494) );
  IVP U651 ( .A(B[94]), .Z(n493) );
  IVP U652 ( .A(B[95]), .Z(n492) );
  IVP U653 ( .A(B[45]), .Z(n542) );
  IVP U654 ( .A(B[46]), .Z(n541) );
  IVP U655 ( .A(B[47]), .Z(n540) );
  IVP U656 ( .A(B[48]), .Z(n539) );
  IVP U657 ( .A(B[49]), .Z(n538) );
  IVP U658 ( .A(B[50]), .Z(n537) );
  IVP U659 ( .A(B[51]), .Z(n536) );
  IVP U660 ( .A(B[39]), .Z(n548) );
  IVP U661 ( .A(B[58]), .Z(n529) );
  IVP U662 ( .A(B[40]), .Z(n547) );
  IVP U663 ( .A(B[41]), .Z(n546) );
  IVP U664 ( .A(B[42]), .Z(n545) );
  IVP U665 ( .A(B[43]), .Z(n544) );
  IVP U666 ( .A(B[44]), .Z(n543) );
  IVP U667 ( .A(B[52]), .Z(n535) );
  IVP U668 ( .A(B[53]), .Z(n534) );
  IVP U669 ( .A(B[57]), .Z(n530) );
  IVP U670 ( .A(B[59]), .Z(n528) );
  IVP U671 ( .A(B[54]), .Z(n533) );
  IVP U672 ( .A(B[56]), .Z(n531) );
  IVP U673 ( .A(B[72]), .Z(n515) );
  AN2P U674 ( .A(\CARRYB[29][0] ), .B(\SUMB[29][1] ), .Z(\A2[29] ) );
  AN2P U675 ( .A(\CARRYB[29][1] ), .B(\SUMB[29][2] ), .Z(\A2[30] ) );
  AN2P U676 ( .A(\CARRYB[29][2] ), .B(\SUMB[29][3] ), .Z(\A2[31] ) );
  AN2P U677 ( .A(\CARRYB[29][3] ), .B(\SUMB[29][4] ), .Z(\A2[32] ) );
  AN2P U678 ( .A(\CARRYB[29][4] ), .B(\SUMB[29][5] ), .Z(\A2[33] ) );
  AN2P U679 ( .A(\CARRYB[29][5] ), .B(\SUMB[29][6] ), .Z(\A2[34] ) );
  AN2P U680 ( .A(\CARRYB[29][6] ), .B(\SUMB[29][7] ), .Z(\A2[35] ) );
  AN2P U681 ( .A(\CARRYB[29][7] ), .B(\SUMB[29][8] ), .Z(\A2[36] ) );
  AN2P U682 ( .A(\CARRYB[29][8] ), .B(\SUMB[29][9] ), .Z(\A2[37] ) );
  AN2P U683 ( .A(\CARRYB[29][9] ), .B(\SUMB[29][10] ), .Z(\A2[38] ) );
  AN2P U684 ( .A(\CARRYB[29][10] ), .B(\SUMB[29][11] ), .Z(\A2[39] ) );
  AN2P U685 ( .A(\CARRYB[29][11] ), .B(\SUMB[29][12] ), .Z(\A2[40] ) );
  AN2P U686 ( .A(\CARRYB[29][12] ), .B(\SUMB[29][13] ), .Z(\A2[41] ) );
  AN2P U687 ( .A(\CARRYB[29][13] ), .B(\SUMB[29][14] ), .Z(\A2[42] ) );
  AN2P U688 ( .A(\CARRYB[29][14] ), .B(\SUMB[29][15] ), .Z(\A2[43] ) );
  AN2P U689 ( .A(\CARRYB[29][15] ), .B(\SUMB[29][16] ), .Z(\A2[44] ) );
  AN2P U690 ( .A(\CARRYB[29][16] ), .B(\SUMB[29][17] ), .Z(\A2[45] ) );
  AN2P U691 ( .A(\CARRYB[29][17] ), .B(\SUMB[29][18] ), .Z(\A2[46] ) );
  AN2P U692 ( .A(\CARRYB[29][18] ), .B(\SUMB[29][19] ), .Z(\A2[47] ) );
  AN2P U693 ( .A(\CARRYB[29][19] ), .B(\SUMB[29][20] ), .Z(\A2[48] ) );
  AN2P U694 ( .A(\CARRYB[29][20] ), .B(\SUMB[29][21] ), .Z(\A2[49] ) );
  AN2P U695 ( .A(\CARRYB[29][21] ), .B(\SUMB[29][22] ), .Z(\A2[50] ) );
  AN2P U696 ( .A(\CARRYB[29][22] ), .B(\SUMB[29][23] ), .Z(\A2[51] ) );
  AN2P U697 ( .A(\CARRYB[29][23] ), .B(\SUMB[29][24] ), .Z(\A2[52] ) );
  AN2P U698 ( .A(\CARRYB[29][24] ), .B(\SUMB[29][25] ), .Z(\A2[53] ) );
  AN2P U699 ( .A(\CARRYB[29][25] ), .B(\SUMB[29][26] ), .Z(\A2[54] ) );
  AN2P U700 ( .A(\CARRYB[29][26] ), .B(\SUMB[29][27] ), .Z(\A2[55] ) );
  AN2P U701 ( .A(\CARRYB[29][27] ), .B(\SUMB[29][28] ), .Z(\A2[56] ) );
  AN2P U702 ( .A(\CARRYB[29][28] ), .B(\SUMB[29][29] ), .Z(\A2[57] ) );
  AN2P U703 ( .A(\CARRYB[29][29] ), .B(\SUMB[29][30] ), .Z(\A2[58] ) );
  AN2P U704 ( .A(\CARRYB[29][30] ), .B(\SUMB[29][31] ), .Z(\A2[59] ) );
  AN2P U705 ( .A(\CARRYB[29][31] ), .B(\SUMB[29][32] ), .Z(\A2[60] ) );
  AN2P U706 ( .A(\CARRYB[29][32] ), .B(\SUMB[29][33] ), .Z(\A2[61] ) );
  AN2P U707 ( .A(\CARRYB[29][33] ), .B(\SUMB[29][34] ), .Z(\A2[62] ) );
  AN2P U708 ( .A(\CARRYB[29][34] ), .B(\SUMB[29][35] ), .Z(\A2[63] ) );
  AN2P U709 ( .A(\CARRYB[29][35] ), .B(\SUMB[29][36] ), .Z(\A2[64] ) );
  AN2P U710 ( .A(\CARRYB[29][36] ), .B(\SUMB[29][37] ), .Z(\A2[65] ) );
  AN2P U711 ( .A(\CARRYB[29][37] ), .B(\SUMB[29][38] ), .Z(\A2[66] ) );
  AN2P U712 ( .A(\CARRYB[29][38] ), .B(\SUMB[29][39] ), .Z(\A2[67] ) );
  AN2P U713 ( .A(\CARRYB[29][39] ), .B(\SUMB[29][40] ), .Z(\A2[68] ) );
  AN2P U714 ( .A(\CARRYB[29][40] ), .B(\SUMB[29][41] ), .Z(\A2[69] ) );
  AN2P U715 ( .A(\CARRYB[29][41] ), .B(\SUMB[29][42] ), .Z(\A2[70] ) );
  AN2P U716 ( .A(\CARRYB[29][42] ), .B(\SUMB[29][43] ), .Z(\A2[71] ) );
  AN2P U717 ( .A(\CARRYB[29][43] ), .B(\SUMB[29][44] ), .Z(\A2[72] ) );
  AN2P U718 ( .A(\CARRYB[29][44] ), .B(\SUMB[29][45] ), .Z(\A2[73] ) );
  AN2P U719 ( .A(\CARRYB[29][45] ), .B(\SUMB[29][46] ), .Z(\A2[74] ) );
  AN2P U720 ( .A(\CARRYB[29][46] ), .B(\SUMB[29][47] ), .Z(\A2[75] ) );
  AN2P U721 ( .A(\CARRYB[29][47] ), .B(\SUMB[29][48] ), .Z(\A2[76] ) );
  AN2P U722 ( .A(\CARRYB[29][48] ), .B(\SUMB[29][49] ), .Z(\A2[77] ) );
  AN2P U723 ( .A(\CARRYB[29][49] ), .B(\SUMB[29][50] ), .Z(\A2[78] ) );
  AN2P U724 ( .A(\CARRYB[29][50] ), .B(\SUMB[29][51] ), .Z(\A2[79] ) );
  AN2P U725 ( .A(\CARRYB[29][51] ), .B(\SUMB[29][52] ), .Z(\A2[80] ) );
  AN2P U726 ( .A(\CARRYB[29][52] ), .B(\SUMB[29][53] ), .Z(\A2[81] ) );
  AN2P U727 ( .A(\CARRYB[29][53] ), .B(\SUMB[29][54] ), .Z(\A2[82] ) );
  AN2P U728 ( .A(\CARRYB[29][54] ), .B(\SUMB[29][55] ), .Z(\A2[83] ) );
  AN2P U729 ( .A(\CARRYB[29][55] ), .B(\SUMB[29][56] ), .Z(\A2[84] ) );
  AN2P U730 ( .A(\CARRYB[29][56] ), .B(\SUMB[29][57] ), .Z(\A2[85] ) );
  AN2P U731 ( .A(\CARRYB[29][57] ), .B(\SUMB[29][58] ), .Z(\A2[86] ) );
  AN2P U732 ( .A(\CARRYB[29][58] ), .B(\SUMB[29][59] ), .Z(\A2[87] ) );
  AN2P U733 ( .A(\CARRYB[29][59] ), .B(\SUMB[29][60] ), .Z(\A2[88] ) );
  AN2P U734 ( .A(\CARRYB[29][60] ), .B(\SUMB[29][61] ), .Z(\A2[89] ) );
  AN2P U735 ( .A(\CARRYB[29][61] ), .B(\SUMB[29][62] ), .Z(\A2[90] ) );
  AN2P U736 ( .A(\CARRYB[29][62] ), .B(\SUMB[29][63] ), .Z(\A2[91] ) );
  AN2P U737 ( .A(\CARRYB[29][63] ), .B(\SUMB[29][64] ), .Z(\A2[92] ) );
  AN2P U738 ( .A(\CARRYB[29][64] ), .B(\SUMB[29][65] ), .Z(\A2[93] ) );
  AN2P U739 ( .A(\CARRYB[29][66] ), .B(\SUMB[29][67] ), .Z(\A2[95] ) );
  AN2P U740 ( .A(\CARRYB[29][67] ), .B(\SUMB[29][68] ), .Z(\A2[96] ) );
  AN2P U741 ( .A(\CARRYB[29][68] ), .B(\SUMB[29][69] ), .Z(\A2[97] ) );
  AN2P U742 ( .A(\CARRYB[29][69] ), .B(\SUMB[29][70] ), .Z(\A2[98] ) );
  AN2P U743 ( .A(\CARRYB[29][70] ), .B(\SUMB[29][71] ), .Z(\A2[99] ) );
  AN2P U744 ( .A(\CARRYB[29][71] ), .B(\SUMB[29][72] ), .Z(\A2[100] ) );
  AN2P U745 ( .A(\CARRYB[29][72] ), .B(\SUMB[29][73] ), .Z(\A2[101] ) );
  AN2P U746 ( .A(\CARRYB[29][73] ), .B(\SUMB[29][74] ), .Z(\A2[102] ) );
  AN2P U747 ( .A(\CARRYB[29][74] ), .B(\SUMB[29][75] ), .Z(\A2[103] ) );
  AN2P U748 ( .A(\CARRYB[29][75] ), .B(\SUMB[29][76] ), .Z(\A2[104] ) );
  AN2P U749 ( .A(\CARRYB[29][76] ), .B(\SUMB[29][77] ), .Z(\A2[105] ) );
  AN2P U750 ( .A(\CARRYB[29][77] ), .B(\SUMB[29][78] ), .Z(\A2[106] ) );
  AN2P U751 ( .A(\CARRYB[29][78] ), .B(\SUMB[29][79] ), .Z(\A2[107] ) );
  AN2P U752 ( .A(\CARRYB[29][79] ), .B(\SUMB[29][80] ), .Z(\A2[108] ) );
  AN2P U753 ( .A(\CARRYB[29][80] ), .B(\SUMB[29][81] ), .Z(\A2[109] ) );
  AN2P U754 ( .A(\CARRYB[29][81] ), .B(\SUMB[29][82] ), .Z(\A2[110] ) );
  AN2P U755 ( .A(\CARRYB[29][82] ), .B(\SUMB[29][83] ), .Z(\A2[111] ) );
  AN2P U756 ( .A(\CARRYB[29][83] ), .B(\SUMB[29][84] ), .Z(\A2[112] ) );
  AN2P U757 ( .A(\CARRYB[29][84] ), .B(\SUMB[29][85] ), .Z(\A2[113] ) );
  AN2P U758 ( .A(\CARRYB[29][85] ), .B(\SUMB[29][86] ), .Z(\A2[114] ) );
  AN2P U759 ( .A(\CARRYB[29][86] ), .B(\SUMB[29][87] ), .Z(\A2[115] ) );
  AN2P U760 ( .A(\CARRYB[29][87] ), .B(\SUMB[29][88] ), .Z(\A2[116] ) );
  AN2P U761 ( .A(\CARRYB[29][88] ), .B(\SUMB[29][89] ), .Z(\A2[117] ) );
  AN2P U762 ( .A(\CARRYB[29][89] ), .B(\SUMB[29][90] ), .Z(\A2[118] ) );
  AN2P U763 ( .A(\CARRYB[29][90] ), .B(\SUMB[29][91] ), .Z(\A2[119] ) );
  AN2P U764 ( .A(\CARRYB[29][91] ), .B(\SUMB[29][92] ), .Z(\A2[120] ) );
  AN2P U765 ( .A(\CARRYB[29][92] ), .B(\SUMB[29][93] ), .Z(\A2[121] ) );
  AN2P U766 ( .A(\CARRYB[29][93] ), .B(\SUMB[29][94] ), .Z(\A2[122] ) );
  AN2P U767 ( .A(\CARRYB[29][94] ), .B(\ab[29][95] ), .Z(\A2[123] ) );
  AN2P U768 ( .A(n3), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U769 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U770 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U771 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U772 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U773 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U774 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U775 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U776 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U777 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U778 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U779 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U780 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U781 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U782 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U783 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\CARRYB[1][16] ) );
  AN2P U784 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\CARRYB[1][17] ) );
  AN2P U785 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\CARRYB[1][18] ) );
  AN2P U786 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\CARRYB[1][19] ) );
  AN2P U787 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\CARRYB[1][20] ) );
  AN2P U788 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\CARRYB[1][21] ) );
  AN2P U789 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(\CARRYB[1][22] ) );
  AN2P U790 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(\CARRYB[1][23] ) );
  AN2P U791 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(\CARRYB[1][24] ) );
  AN2P U792 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(\CARRYB[1][25] ) );
  AN2P U793 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\CARRYB[1][26] ) );
  AN2P U794 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(\CARRYB[1][27] ) );
  AN2P U795 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(\CARRYB[1][28] ) );
  AN2P U796 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(\CARRYB[1][29] ) );
  AN2P U797 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(\CARRYB[1][30] ) );
  AN2P U798 ( .A(\ab[1][31] ), .B(\ab[0][32] ), .Z(\CARRYB[1][31] ) );
  AN2P U799 ( .A(\ab[1][32] ), .B(\ab[0][33] ), .Z(\CARRYB[1][32] ) );
  AN2P U800 ( .A(\ab[1][33] ), .B(\ab[0][34] ), .Z(\CARRYB[1][33] ) );
  AN2P U801 ( .A(\ab[1][34] ), .B(\ab[0][35] ), .Z(\CARRYB[1][34] ) );
  AN2P U802 ( .A(\ab[1][35] ), .B(\ab[0][36] ), .Z(\CARRYB[1][35] ) );
  AN2P U803 ( .A(\ab[1][36] ), .B(\ab[0][37] ), .Z(\CARRYB[1][36] ) );
  AN2P U804 ( .A(\ab[1][37] ), .B(\ab[0][38] ), .Z(\CARRYB[1][37] ) );
  AN2P U805 ( .A(\ab[1][38] ), .B(\ab[0][39] ), .Z(\CARRYB[1][38] ) );
  AN2P U806 ( .A(\ab[1][39] ), .B(\ab[0][40] ), .Z(\CARRYB[1][39] ) );
  AN2P U807 ( .A(\ab[1][40] ), .B(\ab[0][41] ), .Z(\CARRYB[1][40] ) );
  AN2P U808 ( .A(\ab[1][41] ), .B(\ab[0][42] ), .Z(\CARRYB[1][41] ) );
  AN2P U809 ( .A(\ab[1][42] ), .B(\ab[0][43] ), .Z(\CARRYB[1][42] ) );
  AN2P U810 ( .A(\ab[1][43] ), .B(\ab[0][44] ), .Z(\CARRYB[1][43] ) );
  AN2P U811 ( .A(\ab[1][44] ), .B(\ab[0][45] ), .Z(\CARRYB[1][44] ) );
  AN2P U812 ( .A(\ab[1][45] ), .B(\ab[0][46] ), .Z(\CARRYB[1][45] ) );
  AN2P U813 ( .A(\ab[1][46] ), .B(\ab[0][47] ), .Z(\CARRYB[1][46] ) );
  AN2P U814 ( .A(\ab[1][47] ), .B(\ab[0][48] ), .Z(\CARRYB[1][47] ) );
  AN2P U815 ( .A(\ab[1][48] ), .B(\ab[0][49] ), .Z(\CARRYB[1][48] ) );
  AN2P U816 ( .A(\ab[1][49] ), .B(\ab[0][50] ), .Z(\CARRYB[1][49] ) );
  AN2P U817 ( .A(\ab[1][50] ), .B(\ab[0][51] ), .Z(\CARRYB[1][50] ) );
  AN2P U818 ( .A(\ab[1][51] ), .B(\ab[0][52] ), .Z(\CARRYB[1][51] ) );
  AN2P U819 ( .A(\ab[1][52] ), .B(\ab[0][53] ), .Z(\CARRYB[1][52] ) );
  AN2P U820 ( .A(\ab[1][53] ), .B(\ab[0][54] ), .Z(\CARRYB[1][53] ) );
  AN2P U821 ( .A(\ab[1][54] ), .B(\ab[0][55] ), .Z(\CARRYB[1][54] ) );
  AN2P U822 ( .A(\ab[1][55] ), .B(\ab[0][56] ), .Z(\CARRYB[1][55] ) );
  AN2P U823 ( .A(\ab[1][56] ), .B(\ab[0][57] ), .Z(\CARRYB[1][56] ) );
  AN2P U824 ( .A(\ab[1][57] ), .B(\ab[0][58] ), .Z(\CARRYB[1][57] ) );
  AN2P U825 ( .A(\ab[1][58] ), .B(\ab[0][59] ), .Z(\CARRYB[1][58] ) );
  AN2P U826 ( .A(\ab[1][59] ), .B(\ab[0][60] ), .Z(\CARRYB[1][59] ) );
  AN2P U827 ( .A(\ab[1][60] ), .B(\ab[0][61] ), .Z(\CARRYB[1][60] ) );
  AN2P U828 ( .A(\ab[1][61] ), .B(\ab[0][62] ), .Z(\CARRYB[1][61] ) );
  AN2P U829 ( .A(\ab[1][62] ), .B(\ab[0][63] ), .Z(\CARRYB[1][62] ) );
  AN2P U830 ( .A(\ab[1][63] ), .B(\ab[0][64] ), .Z(\CARRYB[1][63] ) );
  AN2P U831 ( .A(\ab[1][64] ), .B(\ab[0][65] ), .Z(\CARRYB[1][64] ) );
  AN2P U832 ( .A(\ab[1][65] ), .B(\ab[0][66] ), .Z(\CARRYB[1][65] ) );
  AN2P U833 ( .A(\ab[1][66] ), .B(\ab[0][67] ), .Z(\CARRYB[1][66] ) );
  AN2P U834 ( .A(\ab[1][67] ), .B(\ab[0][68] ), .Z(\CARRYB[1][67] ) );
  AN2P U835 ( .A(\ab[1][68] ), .B(\ab[0][69] ), .Z(\CARRYB[1][68] ) );
  AN2P U836 ( .A(\ab[1][69] ), .B(\ab[0][70] ), .Z(\CARRYB[1][69] ) );
  AN2P U837 ( .A(\ab[1][70] ), .B(\ab[0][71] ), .Z(\CARRYB[1][70] ) );
  AN2P U838 ( .A(\ab[1][71] ), .B(\ab[0][72] ), .Z(\CARRYB[1][71] ) );
  AN2P U839 ( .A(\ab[1][72] ), .B(\ab[0][73] ), .Z(\CARRYB[1][72] ) );
  AN2P U840 ( .A(\ab[1][73] ), .B(\ab[0][74] ), .Z(\CARRYB[1][73] ) );
  AN2P U841 ( .A(\ab[1][74] ), .B(\ab[0][75] ), .Z(\CARRYB[1][74] ) );
  AN2P U842 ( .A(\ab[1][75] ), .B(\ab[0][76] ), .Z(\CARRYB[1][75] ) );
  AN2P U843 ( .A(\ab[1][76] ), .B(\ab[0][77] ), .Z(\CARRYB[1][76] ) );
  AN2P U844 ( .A(\ab[1][77] ), .B(\ab[0][78] ), .Z(\CARRYB[1][77] ) );
  AN2P U845 ( .A(\ab[1][78] ), .B(\ab[0][79] ), .Z(\CARRYB[1][78] ) );
  AN2P U846 ( .A(\ab[1][79] ), .B(\ab[0][80] ), .Z(\CARRYB[1][79] ) );
  AN2P U847 ( .A(\ab[1][80] ), .B(\ab[0][81] ), .Z(\CARRYB[1][80] ) );
  AN2P U848 ( .A(\ab[1][81] ), .B(\ab[0][82] ), .Z(\CARRYB[1][81] ) );
  AN2P U849 ( .A(\ab[1][82] ), .B(\ab[0][83] ), .Z(\CARRYB[1][82] ) );
  AN2P U850 ( .A(\ab[1][83] ), .B(\ab[0][84] ), .Z(\CARRYB[1][83] ) );
  AN2P U851 ( .A(\ab[1][84] ), .B(\ab[0][85] ), .Z(\CARRYB[1][84] ) );
  AN2P U852 ( .A(\ab[1][85] ), .B(\ab[0][86] ), .Z(\CARRYB[1][85] ) );
  AN2P U853 ( .A(\ab[1][86] ), .B(\ab[0][87] ), .Z(\CARRYB[1][86] ) );
  AN2P U854 ( .A(\ab[1][87] ), .B(\ab[0][88] ), .Z(\CARRYB[1][87] ) );
  AN2P U855 ( .A(\ab[1][88] ), .B(\ab[0][89] ), .Z(\CARRYB[1][88] ) );
  AN2P U856 ( .A(\ab[1][89] ), .B(\ab[0][90] ), .Z(\CARRYB[1][89] ) );
  AN2P U857 ( .A(\ab[1][90] ), .B(\ab[0][91] ), .Z(\CARRYB[1][90] ) );
  AN2P U858 ( .A(\ab[1][91] ), .B(\ab[0][92] ), .Z(\CARRYB[1][91] ) );
  AN2P U859 ( .A(\ab[1][92] ), .B(\ab[0][93] ), .Z(\CARRYB[1][92] ) );
  AN2P U860 ( .A(\ab[1][93] ), .B(\ab[0][94] ), .Z(\CARRYB[1][93] ) );
  AN2P U861 ( .A(\ab[1][94] ), .B(\ab[0][95] ), .Z(\CARRYB[1][94] ) );
  AN2P U862 ( .A(\CARRYB[29][65] ), .B(\SUMB[29][66] ), .Z(\A2[94] ) );
  IVA U863 ( .A(n302), .Z(n301) );
  IVA U864 ( .A(B[0]), .Z(n302) );
  IVA U865 ( .A(n306), .Z(n305) );
  IVA U866 ( .A(B[1]), .Z(n306) );
  IVA U867 ( .A(n310), .Z(n309) );
  IVA U868 ( .A(B[2]), .Z(n310) );
  IVA U869 ( .A(n314), .Z(n313) );
  IVA U870 ( .A(B[3]), .Z(n314) );
  IVA U871 ( .A(n318), .Z(n317) );
  IVA U872 ( .A(B[4]), .Z(n318) );
  IVA U873 ( .A(n322), .Z(n321) );
  IVA U874 ( .A(B[5]), .Z(n322) );
  IVA U875 ( .A(n326), .Z(n325) );
  IVA U876 ( .A(B[6]), .Z(n326) );
  IVA U877 ( .A(n330), .Z(n329) );
  IVA U878 ( .A(B[7]), .Z(n330) );
  IVA U879 ( .A(n334), .Z(n333) );
  IVA U880 ( .A(B[8]), .Z(n334) );
  IVA U881 ( .A(n338), .Z(n337) );
  IVA U882 ( .A(B[9]), .Z(n338) );
  IVA U883 ( .A(n342), .Z(n341) );
  IVA U884 ( .A(B[10]), .Z(n342) );
  IVA U885 ( .A(n346), .Z(n345) );
  IVA U886 ( .A(B[11]), .Z(n346) );
  IVA U887 ( .A(n350), .Z(n349) );
  IVA U888 ( .A(B[12]), .Z(n350) );
  IVA U889 ( .A(n354), .Z(n353) );
  IVA U890 ( .A(B[13]), .Z(n354) );
  IVA U891 ( .A(n358), .Z(n357) );
  IVA U892 ( .A(B[14]), .Z(n358) );
  IVA U893 ( .A(n362), .Z(n361) );
  IVA U894 ( .A(B[15]), .Z(n362) );
  IVA U895 ( .A(n366), .Z(n365) );
  IVA U896 ( .A(B[16]), .Z(n366) );
  IVA U897 ( .A(n370), .Z(n369) );
  IVA U898 ( .A(B[17]), .Z(n370) );
  IVA U899 ( .A(n374), .Z(n373) );
  IVA U900 ( .A(B[18]), .Z(n374) );
  IVA U901 ( .A(n378), .Z(n377) );
  IVA U902 ( .A(B[19]), .Z(n378) );
  IVA U903 ( .A(n382), .Z(n381) );
  IVA U904 ( .A(B[20]), .Z(n382) );
  IVA U905 ( .A(n386), .Z(n385) );
  IVA U906 ( .A(B[21]), .Z(n386) );
  IVA U907 ( .A(n390), .Z(n389) );
  IVA U908 ( .A(B[22]), .Z(n390) );
  IVA U909 ( .A(n394), .Z(n393) );
  IVA U910 ( .A(B[23]), .Z(n394) );
  IVA U911 ( .A(n398), .Z(n397) );
  IVA U912 ( .A(B[24]), .Z(n398) );
  IVA U913 ( .A(n402), .Z(n401) );
  IVA U914 ( .A(B[25]), .Z(n402) );
  IVA U915 ( .A(n406), .Z(n405) );
  IVA U916 ( .A(B[26]), .Z(n406) );
  IVA U917 ( .A(n410), .Z(n409) );
  IVA U918 ( .A(B[27]), .Z(n410) );
  IVA U919 ( .A(n414), .Z(n413) );
  IVA U920 ( .A(B[28]), .Z(n414) );
  IVA U921 ( .A(n418), .Z(n417) );
  IVA U922 ( .A(B[29]), .Z(n418) );
  IVA U923 ( .A(n422), .Z(n421) );
  IVA U924 ( .A(B[30]), .Z(n422) );
  IVA U925 ( .A(n426), .Z(n425) );
  IVA U926 ( .A(B[31]), .Z(n426) );
  IVA U927 ( .A(n430), .Z(n429) );
  IVA U928 ( .A(B[32]), .Z(n430) );
  IVA U929 ( .A(n434), .Z(n433) );
  IVA U930 ( .A(B[33]), .Z(n434) );
  IVA U931 ( .A(n438), .Z(n437) );
  IVA U932 ( .A(B[34]), .Z(n438) );
  IVA U933 ( .A(n442), .Z(n441) );
  IVA U934 ( .A(B[35]), .Z(n442) );
  IVA U935 ( .A(n446), .Z(n445) );
  IVA U936 ( .A(B[36]), .Z(n446) );
  IVA U937 ( .A(n450), .Z(n449) );
  IVA U938 ( .A(B[37]), .Z(n450) );
  IVA U939 ( .A(n454), .Z(n453) );
  IVA U940 ( .A(B[38]), .Z(n454) );
  AN2P U941 ( .A(n171), .B(n491), .Z(\ab[0][95] ) );
  AN2P U942 ( .A(n180), .B(n455), .Z(\ab[1][94] ) );
  AN2P U943 ( .A(n171), .B(n455), .Z(\ab[0][94] ) );
  AN2P U944 ( .A(n180), .B(n456), .Z(\ab[1][93] ) );
  AN2P U945 ( .A(n171), .B(n456), .Z(\ab[0][93] ) );
  AN2P U946 ( .A(n180), .B(n457), .Z(\ab[1][92] ) );
  AN2P U947 ( .A(n171), .B(n457), .Z(\ab[0][92] ) );
  AN2P U948 ( .A(n180), .B(n458), .Z(\ab[1][91] ) );
  AN2P U949 ( .A(n171), .B(n458), .Z(\ab[0][91] ) );
  AN2P U950 ( .A(n180), .B(n459), .Z(\ab[1][90] ) );
  AN2P U951 ( .A(n171), .B(n459), .Z(\ab[0][90] ) );
  AN2P U952 ( .A(n180), .B(n460), .Z(\ab[1][89] ) );
  AN2P U953 ( .A(n171), .B(n460), .Z(\ab[0][89] ) );
  AN2P U954 ( .A(n180), .B(n461), .Z(\ab[1][88] ) );
  AN2P U955 ( .A(n171), .B(n461), .Z(\ab[0][88] ) );
  AN2P U956 ( .A(n180), .B(n462), .Z(\ab[1][87] ) );
  AN2P U957 ( .A(n171), .B(n462), .Z(\ab[0][87] ) );
  AN2P U958 ( .A(n180), .B(n463), .Z(\ab[1][86] ) );
  AN2P U959 ( .A(n171), .B(n463), .Z(\ab[0][86] ) );
  AN2P U960 ( .A(n180), .B(n464), .Z(\ab[1][85] ) );
  AN2P U961 ( .A(n171), .B(n464), .Z(\ab[0][85] ) );
  AN2P U962 ( .A(n180), .B(n465), .Z(\ab[1][84] ) );
  AN2P U963 ( .A(n170), .B(n465), .Z(\ab[0][84] ) );
  AN2P U964 ( .A(n179), .B(n466), .Z(\ab[1][83] ) );
  AN2P U965 ( .A(n170), .B(n466), .Z(\ab[0][83] ) );
  AN2P U966 ( .A(n179), .B(n467), .Z(\ab[1][82] ) );
  AN2P U967 ( .A(n170), .B(n467), .Z(\ab[0][82] ) );
  AN2P U968 ( .A(n179), .B(n468), .Z(\ab[1][81] ) );
  AN2P U969 ( .A(n170), .B(n468), .Z(\ab[0][81] ) );
  AN2P U970 ( .A(n179), .B(n469), .Z(\ab[1][80] ) );
  AN2P U971 ( .A(n170), .B(n469), .Z(\ab[0][80] ) );
  AN2P U972 ( .A(n179), .B(n470), .Z(\ab[1][79] ) );
  AN2P U973 ( .A(n170), .B(n470), .Z(\ab[0][79] ) );
  AN2P U974 ( .A(n179), .B(n471), .Z(\ab[1][78] ) );
  AN2P U975 ( .A(n170), .B(n471), .Z(\ab[0][78] ) );
  AN2P U976 ( .A(n179), .B(n472), .Z(\ab[1][77] ) );
  AN2P U977 ( .A(n170), .B(n472), .Z(\ab[0][77] ) );
  AN2P U978 ( .A(n179), .B(n473), .Z(\ab[1][76] ) );
  AN2P U979 ( .A(n170), .B(n473), .Z(\ab[0][76] ) );
  AN2P U980 ( .A(n179), .B(n474), .Z(\ab[1][75] ) );
  AN2P U981 ( .A(n170), .B(n474), .Z(\ab[0][75] ) );
  AN2P U982 ( .A(n179), .B(n475), .Z(\ab[1][74] ) );
  AN2P U983 ( .A(n170), .B(n475), .Z(\ab[0][74] ) );
  AN2P U984 ( .A(n179), .B(n476), .Z(\ab[1][73] ) );
  AN2P U985 ( .A(n170), .B(n476), .Z(\ab[0][73] ) );
  AN2P U986 ( .A(n179), .B(n477), .Z(\ab[1][72] ) );
  AN2P U987 ( .A(n169), .B(n477), .Z(\ab[0][72] ) );
  AN2P U988 ( .A(n178), .B(n478), .Z(\ab[1][71] ) );
  AN2P U989 ( .A(n169), .B(n478), .Z(\ab[0][71] ) );
  AN2P U990 ( .A(n178), .B(n479), .Z(\ab[1][70] ) );
  AN2P U991 ( .A(n169), .B(n479), .Z(\ab[0][70] ) );
  AN2P U992 ( .A(n178), .B(n480), .Z(\ab[1][69] ) );
  AN2P U993 ( .A(n169), .B(n480), .Z(\ab[0][69] ) );
  AN2P U994 ( .A(n178), .B(n481), .Z(\ab[1][68] ) );
  AN2P U995 ( .A(n169), .B(n481), .Z(\ab[0][68] ) );
  AN2P U996 ( .A(n178), .B(n482), .Z(\ab[1][67] ) );
  AN2P U997 ( .A(n169), .B(n482), .Z(\ab[0][67] ) );
  AN2P U998 ( .A(n178), .B(n483), .Z(\ab[1][66] ) );
  AN2P U999 ( .A(n169), .B(n483), .Z(\ab[0][66] ) );
  AN2P U1000 ( .A(n178), .B(n484), .Z(\ab[1][65] ) );
  AN2P U1001 ( .A(n169), .B(n484), .Z(\ab[0][65] ) );
  AN2P U1002 ( .A(n178), .B(n485), .Z(\ab[1][64] ) );
  AN2P U1003 ( .A(n169), .B(n485), .Z(\ab[0][64] ) );
  AN2P U1004 ( .A(n178), .B(n486), .Z(\ab[1][63] ) );
  AN2P U1005 ( .A(n169), .B(n486), .Z(\ab[0][63] ) );
  AN2P U1006 ( .A(n178), .B(n487), .Z(\ab[1][62] ) );
  AN2P U1007 ( .A(n169), .B(n487), .Z(\ab[0][62] ) );
  AN2P U1008 ( .A(n178), .B(n488), .Z(\ab[1][61] ) );
  AN2P U1009 ( .A(n169), .B(n488), .Z(\ab[0][61] ) );
  AN2P U1010 ( .A(n178), .B(n489), .Z(\ab[1][60] ) );
  AN2P U1011 ( .A(n168), .B(n489), .Z(\ab[0][60] ) );
  AN2P U1012 ( .A(n177), .B(B[59]), .Z(\ab[1][59] ) );
  AN2P U1013 ( .A(n168), .B(B[59]), .Z(\ab[0][59] ) );
  AN2P U1014 ( .A(n177), .B(B[58]), .Z(\ab[1][58] ) );
  AN2P U1015 ( .A(n168), .B(B[58]), .Z(\ab[0][58] ) );
  AN2P U1016 ( .A(n177), .B(B[57]), .Z(\ab[1][57] ) );
  AN2P U1017 ( .A(n168), .B(B[57]), .Z(\ab[0][57] ) );
  AN2P U1018 ( .A(n177), .B(B[56]), .Z(\ab[1][56] ) );
  AN2P U1019 ( .A(n168), .B(B[56]), .Z(\ab[0][56] ) );
  AN2P U1020 ( .A(n177), .B(n490), .Z(\ab[1][55] ) );
  AN2P U1021 ( .A(n168), .B(n490), .Z(\ab[0][55] ) );
  AN2P U1022 ( .A(n177), .B(B[54]), .Z(\ab[1][54] ) );
  AN2P U1023 ( .A(n168), .B(B[54]), .Z(\ab[0][54] ) );
  AN2P U1024 ( .A(n177), .B(B[53]), .Z(\ab[1][53] ) );
  AN2P U1025 ( .A(n168), .B(B[53]), .Z(\ab[0][53] ) );
  AN2P U1026 ( .A(n177), .B(B[52]), .Z(\ab[1][52] ) );
  AN2P U1027 ( .A(n168), .B(B[52]), .Z(\ab[0][52] ) );
  AN2P U1028 ( .A(n177), .B(B[51]), .Z(\ab[1][51] ) );
  AN2P U1029 ( .A(n168), .B(B[51]), .Z(\ab[0][51] ) );
  AN2P U1030 ( .A(n177), .B(B[50]), .Z(\ab[1][50] ) );
  AN2P U1031 ( .A(n168), .B(B[50]), .Z(\ab[0][50] ) );
  AN2P U1032 ( .A(n177), .B(B[49]), .Z(\ab[1][49] ) );
  AN2P U1033 ( .A(n168), .B(B[49]), .Z(\ab[0][49] ) );
  AN2P U1034 ( .A(n177), .B(B[48]), .Z(\ab[1][48] ) );
  AN2P U1035 ( .A(n167), .B(B[48]), .Z(\ab[0][48] ) );
  AN2P U1036 ( .A(n176), .B(B[47]), .Z(\ab[1][47] ) );
  AN2P U1037 ( .A(n167), .B(B[47]), .Z(\ab[0][47] ) );
  AN2P U1038 ( .A(n176), .B(B[46]), .Z(\ab[1][46] ) );
  AN2P U1039 ( .A(n167), .B(B[46]), .Z(\ab[0][46] ) );
  AN2P U1040 ( .A(n176), .B(B[45]), .Z(\ab[1][45] ) );
  AN2P U1041 ( .A(n167), .B(B[45]), .Z(\ab[0][45] ) );
  AN2P U1042 ( .A(n176), .B(B[44]), .Z(\ab[1][44] ) );
  AN2P U1043 ( .A(n167), .B(B[44]), .Z(\ab[0][44] ) );
  AN2P U1044 ( .A(n176), .B(B[43]), .Z(\ab[1][43] ) );
  AN2P U1045 ( .A(n167), .B(B[43]), .Z(\ab[0][43] ) );
  AN2P U1046 ( .A(n176), .B(B[42]), .Z(\ab[1][42] ) );
  AN2P U1047 ( .A(n167), .B(B[42]), .Z(\ab[0][42] ) );
  AN2P U1048 ( .A(n176), .B(B[41]), .Z(\ab[1][41] ) );
  AN2P U1049 ( .A(n167), .B(B[41]), .Z(\ab[0][41] ) );
  AN2P U1050 ( .A(n176), .B(B[40]), .Z(\ab[1][40] ) );
  AN2P U1051 ( .A(n167), .B(B[40]), .Z(\ab[0][40] ) );
  AN2P U1052 ( .A(n176), .B(B[39]), .Z(\ab[1][39] ) );
  AN2P U1053 ( .A(n167), .B(B[39]), .Z(\ab[0][39] ) );
  AN2P U1054 ( .A(n176), .B(n453), .Z(\ab[1][38] ) );
  AN2P U1055 ( .A(n167), .B(n453), .Z(\ab[0][38] ) );
  AN2P U1056 ( .A(n176), .B(n449), .Z(\ab[1][37] ) );
  AN2P U1057 ( .A(n167), .B(n449), .Z(\ab[0][37] ) );
  AN2P U1058 ( .A(n176), .B(n445), .Z(\ab[1][36] ) );
  AN2P U1059 ( .A(n166), .B(n445), .Z(\ab[0][36] ) );
  AN2P U1060 ( .A(n175), .B(n441), .Z(\ab[1][35] ) );
  AN2P U1061 ( .A(n166), .B(n441), .Z(\ab[0][35] ) );
  AN2P U1062 ( .A(n175), .B(n437), .Z(\ab[1][34] ) );
  AN2P U1063 ( .A(n166), .B(n437), .Z(\ab[0][34] ) );
  AN2P U1064 ( .A(n175), .B(n433), .Z(\ab[1][33] ) );
  AN2P U1065 ( .A(n166), .B(n433), .Z(\ab[0][33] ) );
  AN2P U1066 ( .A(n175), .B(n429), .Z(\ab[1][32] ) );
  AN2P U1067 ( .A(n166), .B(n429), .Z(\ab[0][32] ) );
  AN2P U1068 ( .A(n175), .B(n425), .Z(\ab[1][31] ) );
  AN2P U1069 ( .A(n166), .B(n425), .Z(\ab[0][31] ) );
  AN2P U1070 ( .A(n175), .B(n421), .Z(\ab[1][30] ) );
  AN2P U1071 ( .A(n166), .B(n421), .Z(\ab[0][30] ) );
  AN2P U1072 ( .A(n175), .B(n417), .Z(\ab[1][29] ) );
  AN2P U1073 ( .A(n166), .B(n417), .Z(\ab[0][29] ) );
  AN2P U1074 ( .A(n175), .B(n413), .Z(\ab[1][28] ) );
  AN2P U1075 ( .A(n166), .B(n413), .Z(\ab[0][28] ) );
  AN2P U1076 ( .A(n175), .B(n409), .Z(\ab[1][27] ) );
  AN2P U1077 ( .A(n166), .B(n409), .Z(\ab[0][27] ) );
  AN2P U1078 ( .A(n175), .B(n405), .Z(\ab[1][26] ) );
  AN2P U1079 ( .A(n166), .B(n405), .Z(\ab[0][26] ) );
  AN2P U1080 ( .A(n175), .B(n401), .Z(\ab[1][25] ) );
  AN2P U1081 ( .A(n166), .B(n401), .Z(\ab[0][25] ) );
  AN2P U1082 ( .A(n175), .B(n397), .Z(\ab[1][24] ) );
  AN2P U1083 ( .A(n165), .B(n397), .Z(\ab[0][24] ) );
  AN2P U1084 ( .A(n174), .B(n393), .Z(\ab[1][23] ) );
  AN2P U1085 ( .A(n165), .B(n393), .Z(\ab[0][23] ) );
  AN2P U1086 ( .A(n174), .B(n389), .Z(\ab[1][22] ) );
  AN2P U1087 ( .A(n165), .B(n389), .Z(\ab[0][22] ) );
  AN2P U1088 ( .A(n174), .B(n385), .Z(\ab[1][21] ) );
  AN2P U1089 ( .A(n165), .B(n385), .Z(\ab[0][21] ) );
  AN2P U1090 ( .A(n174), .B(n381), .Z(\ab[1][20] ) );
  AN2P U1091 ( .A(n165), .B(n381), .Z(\ab[0][20] ) );
  AN2P U1092 ( .A(n174), .B(n377), .Z(\ab[1][19] ) );
  AN2P U1093 ( .A(n165), .B(n377), .Z(\ab[0][19] ) );
  AN2P U1094 ( .A(n174), .B(n373), .Z(\ab[1][18] ) );
  AN2P U1095 ( .A(n165), .B(n373), .Z(\ab[0][18] ) );
  AN2P U1096 ( .A(n174), .B(n369), .Z(\ab[1][17] ) );
  AN2P U1097 ( .A(n165), .B(n369), .Z(\ab[0][17] ) );
  AN2P U1098 ( .A(n174), .B(n365), .Z(\ab[1][16] ) );
  AN2P U1099 ( .A(n165), .B(n365), .Z(\ab[0][16] ) );
  AN2P U1100 ( .A(n174), .B(n361), .Z(\ab[1][15] ) );
  AN2P U1101 ( .A(n165), .B(n361), .Z(\ab[0][15] ) );
  AN2P U1102 ( .A(n174), .B(n357), .Z(\ab[1][14] ) );
  AN2P U1103 ( .A(n165), .B(n357), .Z(\ab[0][14] ) );
  AN2P U1104 ( .A(n174), .B(n353), .Z(\ab[1][13] ) );
  AN2P U1105 ( .A(n165), .B(n353), .Z(\ab[0][13] ) );
  AN2P U1106 ( .A(n174), .B(n349), .Z(\ab[1][12] ) );
  AN2P U1107 ( .A(n164), .B(n349), .Z(\ab[0][12] ) );
  AN2P U1108 ( .A(n173), .B(n345), .Z(\ab[1][11] ) );
  AN2P U1109 ( .A(n164), .B(n345), .Z(\ab[0][11] ) );
  AN2P U1110 ( .A(n173), .B(n341), .Z(\ab[1][10] ) );
  AN2P U1111 ( .A(n164), .B(n341), .Z(\ab[0][10] ) );
  AN2P U1112 ( .A(n173), .B(n337), .Z(\ab[1][9] ) );
  AN2P U1113 ( .A(n164), .B(n337), .Z(\ab[0][9] ) );
  AN2P U1114 ( .A(n173), .B(n333), .Z(\ab[1][8] ) );
  AN2P U1115 ( .A(n164), .B(n333), .Z(\ab[0][8] ) );
  AN2P U1116 ( .A(n173), .B(n329), .Z(\ab[1][7] ) );
  AN2P U1117 ( .A(n164), .B(n329), .Z(\ab[0][7] ) );
  AN2P U1118 ( .A(n173), .B(n325), .Z(\ab[1][6] ) );
  AN2P U1119 ( .A(n164), .B(n325), .Z(\ab[0][6] ) );
  AN2P U1120 ( .A(n173), .B(n321), .Z(\ab[1][5] ) );
  AN2P U1121 ( .A(n164), .B(n321), .Z(\ab[0][5] ) );
  AN2P U1122 ( .A(n173), .B(n317), .Z(\ab[1][4] ) );
  AN2P U1123 ( .A(n164), .B(n317), .Z(\ab[0][4] ) );
  AN2P U1124 ( .A(n173), .B(n313), .Z(\ab[1][3] ) );
  AN2P U1125 ( .A(n164), .B(n313), .Z(\ab[0][3] ) );
  AN2P U1126 ( .A(n173), .B(n309), .Z(\ab[1][2] ) );
  AN2P U1127 ( .A(n164), .B(n309), .Z(\ab[0][2] ) );
  AN2P U1128 ( .A(n189), .B(n455), .Z(\ab[2][94] ) );
  AN2P U1129 ( .A(n173), .B(n491), .Z(\ab[1][95] ) );
  AN2P U1130 ( .A(n189), .B(n456), .Z(\ab[2][93] ) );
  AN2P U1131 ( .A(n189), .B(n457), .Z(\ab[2][92] ) );
  AN2P U1132 ( .A(n189), .B(n458), .Z(\ab[2][91] ) );
  AN2P U1133 ( .A(n189), .B(n459), .Z(\ab[2][90] ) );
  AN2P U1134 ( .A(n189), .B(n460), .Z(\ab[2][89] ) );
  AN2P U1135 ( .A(n189), .B(n461), .Z(\ab[2][88] ) );
  AN2P U1136 ( .A(n189), .B(n462), .Z(\ab[2][87] ) );
  AN2P U1137 ( .A(n189), .B(n463), .Z(\ab[2][86] ) );
  AN2P U1138 ( .A(n189), .B(n464), .Z(\ab[2][85] ) );
  AN2P U1139 ( .A(n189), .B(n465), .Z(\ab[2][84] ) );
  AN2P U1140 ( .A(n189), .B(n466), .Z(\ab[2][83] ) );
  AN2P U1141 ( .A(n188), .B(n467), .Z(\ab[2][82] ) );
  AN2P U1142 ( .A(n188), .B(n468), .Z(\ab[2][81] ) );
  AN2P U1143 ( .A(n188), .B(n469), .Z(\ab[2][80] ) );
  AN2P U1144 ( .A(n188), .B(n470), .Z(\ab[2][79] ) );
  AN2P U1145 ( .A(n188), .B(n471), .Z(\ab[2][78] ) );
  AN2P U1146 ( .A(n188), .B(n472), .Z(\ab[2][77] ) );
  AN2P U1147 ( .A(n188), .B(n473), .Z(\ab[2][76] ) );
  AN2P U1148 ( .A(n188), .B(n474), .Z(\ab[2][75] ) );
  AN2P U1149 ( .A(n188), .B(n475), .Z(\ab[2][74] ) );
  AN2P U1150 ( .A(n188), .B(n476), .Z(\ab[2][73] ) );
  AN2P U1151 ( .A(n188), .B(n477), .Z(\ab[2][72] ) );
  AN2P U1152 ( .A(n188), .B(n478), .Z(\ab[2][71] ) );
  AN2P U1153 ( .A(n187), .B(n479), .Z(\ab[2][70] ) );
  AN2P U1154 ( .A(n187), .B(n480), .Z(\ab[2][69] ) );
  AN2P U1155 ( .A(n187), .B(n481), .Z(\ab[2][68] ) );
  AN2P U1156 ( .A(n187), .B(n482), .Z(\ab[2][67] ) );
  AN2P U1157 ( .A(n187), .B(n483), .Z(\ab[2][66] ) );
  AN2P U1158 ( .A(n187), .B(n484), .Z(\ab[2][65] ) );
  AN2P U1159 ( .A(n187), .B(n485), .Z(\ab[2][64] ) );
  AN2P U1160 ( .A(n187), .B(n486), .Z(\ab[2][63] ) );
  AN2P U1161 ( .A(n187), .B(n487), .Z(\ab[2][62] ) );
  AN2P U1162 ( .A(n187), .B(n488), .Z(\ab[2][61] ) );
  AN2P U1163 ( .A(n187), .B(n489), .Z(\ab[2][60] ) );
  AN2P U1164 ( .A(n187), .B(B[59]), .Z(\ab[2][59] ) );
  AN2P U1165 ( .A(n186), .B(B[58]), .Z(\ab[2][58] ) );
  AN2P U1166 ( .A(n186), .B(B[57]), .Z(\ab[2][57] ) );
  AN2P U1167 ( .A(n186), .B(B[56]), .Z(\ab[2][56] ) );
  AN2P U1168 ( .A(n186), .B(n490), .Z(\ab[2][55] ) );
  AN2P U1169 ( .A(n186), .B(B[54]), .Z(\ab[2][54] ) );
  AN2P U1170 ( .A(n186), .B(B[53]), .Z(\ab[2][53] ) );
  AN2P U1171 ( .A(n186), .B(B[52]), .Z(\ab[2][52] ) );
  AN2P U1172 ( .A(n186), .B(B[51]), .Z(\ab[2][51] ) );
  AN2P U1173 ( .A(n186), .B(B[50]), .Z(\ab[2][50] ) );
  AN2P U1174 ( .A(n186), .B(B[49]), .Z(\ab[2][49] ) );
  AN2P U1175 ( .A(n186), .B(B[48]), .Z(\ab[2][48] ) );
  AN2P U1176 ( .A(n186), .B(B[47]), .Z(\ab[2][47] ) );
  AN2P U1177 ( .A(n185), .B(B[46]), .Z(\ab[2][46] ) );
  AN2P U1178 ( .A(n185), .B(B[45]), .Z(\ab[2][45] ) );
  AN2P U1179 ( .A(n185), .B(B[44]), .Z(\ab[2][44] ) );
  AN2P U1180 ( .A(n185), .B(B[43]), .Z(\ab[2][43] ) );
  AN2P U1181 ( .A(n185), .B(B[42]), .Z(\ab[2][42] ) );
  AN2P U1182 ( .A(n185), .B(B[41]), .Z(\ab[2][41] ) );
  AN2P U1183 ( .A(n185), .B(B[40]), .Z(\ab[2][40] ) );
  AN2P U1184 ( .A(n185), .B(B[39]), .Z(\ab[2][39] ) );
  AN2P U1185 ( .A(n185), .B(n453), .Z(\ab[2][38] ) );
  AN2P U1186 ( .A(n185), .B(n449), .Z(\ab[2][37] ) );
  AN2P U1187 ( .A(n185), .B(n445), .Z(\ab[2][36] ) );
  AN2P U1188 ( .A(n185), .B(n441), .Z(\ab[2][35] ) );
  AN2P U1189 ( .A(n184), .B(n437), .Z(\ab[2][34] ) );
  AN2P U1190 ( .A(n184), .B(n433), .Z(\ab[2][33] ) );
  AN2P U1191 ( .A(n184), .B(n429), .Z(\ab[2][32] ) );
  AN2P U1192 ( .A(n184), .B(n425), .Z(\ab[2][31] ) );
  AN2P U1193 ( .A(n184), .B(n421), .Z(\ab[2][30] ) );
  AN2P U1194 ( .A(n184), .B(n417), .Z(\ab[2][29] ) );
  AN2P U1195 ( .A(n184), .B(n413), .Z(\ab[2][28] ) );
  AN2P U1196 ( .A(n184), .B(n409), .Z(\ab[2][27] ) );
  AN2P U1197 ( .A(n184), .B(n405), .Z(\ab[2][26] ) );
  AN2P U1198 ( .A(n184), .B(n401), .Z(\ab[2][25] ) );
  AN2P U1199 ( .A(n184), .B(n397), .Z(\ab[2][24] ) );
  AN2P U1200 ( .A(n184), .B(n393), .Z(\ab[2][23] ) );
  AN2P U1201 ( .A(n183), .B(n389), .Z(\ab[2][22] ) );
  AN2P U1202 ( .A(n183), .B(n385), .Z(\ab[2][21] ) );
  AN2P U1203 ( .A(n183), .B(n381), .Z(\ab[2][20] ) );
  AN2P U1204 ( .A(n183), .B(n377), .Z(\ab[2][19] ) );
  AN2P U1205 ( .A(n183), .B(n373), .Z(\ab[2][18] ) );
  AN2P U1206 ( .A(n183), .B(n369), .Z(\ab[2][17] ) );
  AN2P U1207 ( .A(n183), .B(n365), .Z(\ab[2][16] ) );
  AN2P U1208 ( .A(n183), .B(n361), .Z(\ab[2][15] ) );
  AN2P U1209 ( .A(n183), .B(n357), .Z(\ab[2][14] ) );
  AN2P U1210 ( .A(n183), .B(n353), .Z(\ab[2][13] ) );
  AN2P U1211 ( .A(n183), .B(n349), .Z(\ab[2][12] ) );
  AN2P U1212 ( .A(n183), .B(n345), .Z(\ab[2][11] ) );
  AN2P U1213 ( .A(n182), .B(n341), .Z(\ab[2][10] ) );
  AN2P U1214 ( .A(n182), .B(n337), .Z(\ab[2][9] ) );
  AN2P U1215 ( .A(n182), .B(n333), .Z(\ab[2][8] ) );
  AN2P U1216 ( .A(n182), .B(n329), .Z(\ab[2][7] ) );
  AN2P U1217 ( .A(n182), .B(n325), .Z(\ab[2][6] ) );
  AN2P U1218 ( .A(n182), .B(n321), .Z(\ab[2][5] ) );
  AN2P U1219 ( .A(n182), .B(n317), .Z(\ab[2][4] ) );
  AN2P U1220 ( .A(n182), .B(n313), .Z(\ab[2][3] ) );
  AN2P U1221 ( .A(n182), .B(n309), .Z(\ab[2][2] ) );
  AN2P U1222 ( .A(n182), .B(n305), .Z(\ab[2][1] ) );
  AN2P U1223 ( .A(n182), .B(n301), .Z(\ab[2][0] ) );
  AN3 U1224 ( .A(n164), .B(n301), .C(n3), .Z(\CARRYB[1][0] ) );
  AN2P U1225 ( .A(n198), .B(n455), .Z(\ab[3][94] ) );
  AN2P U1226 ( .A(n182), .B(n491), .Z(\ab[2][95] ) );
  AN2P U1227 ( .A(n198), .B(n456), .Z(\ab[3][93] ) );
  AN2P U1228 ( .A(n198), .B(n457), .Z(\ab[3][92] ) );
  AN2P U1229 ( .A(n198), .B(n458), .Z(\ab[3][91] ) );
  AN2P U1230 ( .A(n198), .B(n459), .Z(\ab[3][90] ) );
  AN2P U1231 ( .A(n198), .B(n460), .Z(\ab[3][89] ) );
  AN2P U1232 ( .A(n198), .B(n461), .Z(\ab[3][88] ) );
  AN2P U1233 ( .A(n198), .B(n462), .Z(\ab[3][87] ) );
  AN2P U1234 ( .A(n198), .B(n463), .Z(\ab[3][86] ) );
  AN2P U1235 ( .A(n198), .B(n464), .Z(\ab[3][85] ) );
  AN2P U1236 ( .A(n198), .B(n465), .Z(\ab[3][84] ) );
  AN2P U1237 ( .A(n198), .B(n466), .Z(\ab[3][83] ) );
  AN2P U1238 ( .A(n197), .B(n467), .Z(\ab[3][82] ) );
  AN2P U1239 ( .A(n197), .B(n468), .Z(\ab[3][81] ) );
  AN2P U1240 ( .A(n197), .B(n469), .Z(\ab[3][80] ) );
  AN2P U1241 ( .A(n197), .B(n470), .Z(\ab[3][79] ) );
  AN2P U1242 ( .A(n197), .B(n471), .Z(\ab[3][78] ) );
  AN2P U1243 ( .A(n197), .B(n472), .Z(\ab[3][77] ) );
  AN2P U1244 ( .A(n197), .B(n473), .Z(\ab[3][76] ) );
  AN2P U1245 ( .A(n197), .B(n474), .Z(\ab[3][75] ) );
  AN2P U1246 ( .A(n197), .B(n475), .Z(\ab[3][74] ) );
  AN2P U1247 ( .A(n197), .B(n476), .Z(\ab[3][73] ) );
  AN2P U1248 ( .A(n197), .B(n477), .Z(\ab[3][72] ) );
  AN2P U1249 ( .A(n197), .B(n478), .Z(\ab[3][71] ) );
  AN2P U1250 ( .A(n196), .B(n479), .Z(\ab[3][70] ) );
  AN2P U1251 ( .A(n196), .B(n480), .Z(\ab[3][69] ) );
  AN2P U1252 ( .A(n196), .B(n481), .Z(\ab[3][68] ) );
  AN2P U1253 ( .A(n196), .B(n482), .Z(\ab[3][67] ) );
  AN2P U1254 ( .A(n196), .B(n483), .Z(\ab[3][66] ) );
  AN2P U1255 ( .A(n196), .B(n484), .Z(\ab[3][65] ) );
  AN2P U1256 ( .A(n196), .B(n485), .Z(\ab[3][64] ) );
  AN2P U1257 ( .A(n196), .B(n486), .Z(\ab[3][63] ) );
  AN2P U1258 ( .A(n196), .B(n487), .Z(\ab[3][62] ) );
  AN2P U1259 ( .A(n196), .B(n488), .Z(\ab[3][61] ) );
  AN2P U1260 ( .A(n196), .B(n489), .Z(\ab[3][60] ) );
  AN2P U1261 ( .A(n196), .B(B[59]), .Z(\ab[3][59] ) );
  AN2P U1262 ( .A(n195), .B(B[58]), .Z(\ab[3][58] ) );
  AN2P U1263 ( .A(n195), .B(B[57]), .Z(\ab[3][57] ) );
  AN2P U1264 ( .A(n195), .B(B[56]), .Z(\ab[3][56] ) );
  AN2P U1265 ( .A(n195), .B(n490), .Z(\ab[3][55] ) );
  AN2P U1266 ( .A(n195), .B(B[54]), .Z(\ab[3][54] ) );
  AN2P U1267 ( .A(n195), .B(B[53]), .Z(\ab[3][53] ) );
  AN2P U1268 ( .A(n195), .B(B[52]), .Z(\ab[3][52] ) );
  AN2P U1269 ( .A(n195), .B(B[51]), .Z(\ab[3][51] ) );
  AN2P U1270 ( .A(n195), .B(B[50]), .Z(\ab[3][50] ) );
  AN2P U1271 ( .A(n195), .B(B[49]), .Z(\ab[3][49] ) );
  AN2P U1272 ( .A(n195), .B(B[48]), .Z(\ab[3][48] ) );
  AN2P U1273 ( .A(n195), .B(B[47]), .Z(\ab[3][47] ) );
  AN2P U1274 ( .A(n194), .B(B[46]), .Z(\ab[3][46] ) );
  AN2P U1275 ( .A(n194), .B(B[45]), .Z(\ab[3][45] ) );
  AN2P U1276 ( .A(n194), .B(B[44]), .Z(\ab[3][44] ) );
  AN2P U1277 ( .A(n194), .B(B[43]), .Z(\ab[3][43] ) );
  AN2P U1278 ( .A(n194), .B(B[42]), .Z(\ab[3][42] ) );
  AN2P U1279 ( .A(n194), .B(B[41]), .Z(\ab[3][41] ) );
  AN2P U1280 ( .A(n194), .B(B[40]), .Z(\ab[3][40] ) );
  AN2P U1281 ( .A(n194), .B(B[39]), .Z(\ab[3][39] ) );
  AN2P U1282 ( .A(n194), .B(n453), .Z(\ab[3][38] ) );
  AN2P U1283 ( .A(n194), .B(n449), .Z(\ab[3][37] ) );
  AN2P U1284 ( .A(n194), .B(n445), .Z(\ab[3][36] ) );
  AN2P U1285 ( .A(n194), .B(n441), .Z(\ab[3][35] ) );
  AN2P U1286 ( .A(n193), .B(n437), .Z(\ab[3][34] ) );
  AN2P U1287 ( .A(n193), .B(n433), .Z(\ab[3][33] ) );
  AN2P U1288 ( .A(n193), .B(n429), .Z(\ab[3][32] ) );
  AN2P U1289 ( .A(n193), .B(n425), .Z(\ab[3][31] ) );
  AN2P U1290 ( .A(n193), .B(n421), .Z(\ab[3][30] ) );
  AN2P U1291 ( .A(n193), .B(n417), .Z(\ab[3][29] ) );
  AN2P U1292 ( .A(n193), .B(n413), .Z(\ab[3][28] ) );
  AN2P U1293 ( .A(n193), .B(n409), .Z(\ab[3][27] ) );
  AN2P U1294 ( .A(n193), .B(n405), .Z(\ab[3][26] ) );
  AN2P U1295 ( .A(n193), .B(n401), .Z(\ab[3][25] ) );
  AN2P U1296 ( .A(n193), .B(n397), .Z(\ab[3][24] ) );
  AN2P U1297 ( .A(n193), .B(n393), .Z(\ab[3][23] ) );
  AN2P U1298 ( .A(n192), .B(n389), .Z(\ab[3][22] ) );
  AN2P U1299 ( .A(n192), .B(n385), .Z(\ab[3][21] ) );
  AN2P U1300 ( .A(n192), .B(n381), .Z(\ab[3][20] ) );
  AN2P U1301 ( .A(n192), .B(n377), .Z(\ab[3][19] ) );
  AN2P U1302 ( .A(n192), .B(n373), .Z(\ab[3][18] ) );
  AN2P U1303 ( .A(n192), .B(n369), .Z(\ab[3][17] ) );
  AN2P U1304 ( .A(n192), .B(n365), .Z(\ab[3][16] ) );
  AN2P U1305 ( .A(n192), .B(n361), .Z(\ab[3][15] ) );
  AN2P U1306 ( .A(n192), .B(n357), .Z(\ab[3][14] ) );
  AN2P U1307 ( .A(n192), .B(n353), .Z(\ab[3][13] ) );
  AN2P U1308 ( .A(n192), .B(n349), .Z(\ab[3][12] ) );
  AN2P U1309 ( .A(n192), .B(n345), .Z(\ab[3][11] ) );
  AN2P U1310 ( .A(n191), .B(n341), .Z(\ab[3][10] ) );
  AN2P U1311 ( .A(n191), .B(n337), .Z(\ab[3][9] ) );
  AN2P U1312 ( .A(n191), .B(n333), .Z(\ab[3][8] ) );
  AN2P U1313 ( .A(n191), .B(n329), .Z(\ab[3][7] ) );
  AN2P U1314 ( .A(n191), .B(n325), .Z(\ab[3][6] ) );
  AN2P U1315 ( .A(n191), .B(n321), .Z(\ab[3][5] ) );
  AN2P U1316 ( .A(n191), .B(n317), .Z(\ab[3][4] ) );
  AN2P U1317 ( .A(n191), .B(n313), .Z(\ab[3][3] ) );
  AN2P U1318 ( .A(n191), .B(n309), .Z(\ab[3][2] ) );
  AN2P U1319 ( .A(n191), .B(n305), .Z(\ab[3][1] ) );
  AN2P U1320 ( .A(n191), .B(n301), .Z(\ab[3][0] ) );
  AN2P U1321 ( .A(n207), .B(n455), .Z(\ab[4][94] ) );
  AN2P U1322 ( .A(n191), .B(n491), .Z(\ab[3][95] ) );
  AN2P U1323 ( .A(n207), .B(n456), .Z(\ab[4][93] ) );
  AN2P U1324 ( .A(n207), .B(n457), .Z(\ab[4][92] ) );
  AN2P U1325 ( .A(n207), .B(n458), .Z(\ab[4][91] ) );
  AN2P U1326 ( .A(n207), .B(n459), .Z(\ab[4][90] ) );
  AN2P U1327 ( .A(n207), .B(n460), .Z(\ab[4][89] ) );
  AN2P U1328 ( .A(n207), .B(n461), .Z(\ab[4][88] ) );
  AN2P U1329 ( .A(n207), .B(n462), .Z(\ab[4][87] ) );
  AN2P U1330 ( .A(n207), .B(n463), .Z(\ab[4][86] ) );
  AN2P U1331 ( .A(n207), .B(n464), .Z(\ab[4][85] ) );
  AN2P U1332 ( .A(n207), .B(n465), .Z(\ab[4][84] ) );
  AN2P U1333 ( .A(n207), .B(n466), .Z(\ab[4][83] ) );
  AN2P U1334 ( .A(n206), .B(n467), .Z(\ab[4][82] ) );
  AN2P U1335 ( .A(n206), .B(n468), .Z(\ab[4][81] ) );
  AN2P U1336 ( .A(n206), .B(n469), .Z(\ab[4][80] ) );
  AN2P U1337 ( .A(n206), .B(n470), .Z(\ab[4][79] ) );
  AN2P U1338 ( .A(n206), .B(n471), .Z(\ab[4][78] ) );
  AN2P U1339 ( .A(n206), .B(n472), .Z(\ab[4][77] ) );
  AN2P U1340 ( .A(n206), .B(n473), .Z(\ab[4][76] ) );
  AN2P U1341 ( .A(n206), .B(n474), .Z(\ab[4][75] ) );
  AN2P U1342 ( .A(n206), .B(n475), .Z(\ab[4][74] ) );
  AN2P U1343 ( .A(n206), .B(n476), .Z(\ab[4][73] ) );
  AN2P U1344 ( .A(n206), .B(n477), .Z(\ab[4][72] ) );
  AN2P U1345 ( .A(n206), .B(n478), .Z(\ab[4][71] ) );
  AN2P U1346 ( .A(n205), .B(n479), .Z(\ab[4][70] ) );
  AN2P U1347 ( .A(n205), .B(n480), .Z(\ab[4][69] ) );
  AN2P U1348 ( .A(n205), .B(n481), .Z(\ab[4][68] ) );
  AN2P U1349 ( .A(n205), .B(n482), .Z(\ab[4][67] ) );
  AN2P U1350 ( .A(n205), .B(n483), .Z(\ab[4][66] ) );
  AN2P U1351 ( .A(n205), .B(n484), .Z(\ab[4][65] ) );
  AN2P U1352 ( .A(n205), .B(n485), .Z(\ab[4][64] ) );
  AN2P U1353 ( .A(n205), .B(n486), .Z(\ab[4][63] ) );
  AN2P U1354 ( .A(n205), .B(n487), .Z(\ab[4][62] ) );
  AN2P U1355 ( .A(n205), .B(n488), .Z(\ab[4][61] ) );
  AN2P U1356 ( .A(n205), .B(n489), .Z(\ab[4][60] ) );
  AN2P U1357 ( .A(n205), .B(B[59]), .Z(\ab[4][59] ) );
  AN2P U1358 ( .A(n204), .B(B[58]), .Z(\ab[4][58] ) );
  AN2P U1359 ( .A(n204), .B(B[57]), .Z(\ab[4][57] ) );
  AN2P U1360 ( .A(n204), .B(B[56]), .Z(\ab[4][56] ) );
  AN2P U1361 ( .A(n204), .B(n490), .Z(\ab[4][55] ) );
  AN2P U1362 ( .A(n204), .B(B[54]), .Z(\ab[4][54] ) );
  AN2P U1363 ( .A(n204), .B(B[53]), .Z(\ab[4][53] ) );
  AN2P U1364 ( .A(n204), .B(B[52]), .Z(\ab[4][52] ) );
  AN2P U1365 ( .A(n204), .B(B[51]), .Z(\ab[4][51] ) );
  AN2P U1366 ( .A(n204), .B(B[50]), .Z(\ab[4][50] ) );
  AN2P U1367 ( .A(n204), .B(B[49]), .Z(\ab[4][49] ) );
  AN2P U1368 ( .A(n204), .B(B[48]), .Z(\ab[4][48] ) );
  AN2P U1369 ( .A(n204), .B(B[47]), .Z(\ab[4][47] ) );
  AN2P U1370 ( .A(n203), .B(B[46]), .Z(\ab[4][46] ) );
  AN2P U1371 ( .A(n203), .B(B[45]), .Z(\ab[4][45] ) );
  AN2P U1372 ( .A(n203), .B(B[44]), .Z(\ab[4][44] ) );
  AN2P U1373 ( .A(n203), .B(B[43]), .Z(\ab[4][43] ) );
  AN2P U1374 ( .A(n203), .B(B[42]), .Z(\ab[4][42] ) );
  AN2P U1375 ( .A(n203), .B(B[41]), .Z(\ab[4][41] ) );
  AN2P U1376 ( .A(n203), .B(B[40]), .Z(\ab[4][40] ) );
  AN2P U1377 ( .A(n203), .B(B[39]), .Z(\ab[4][39] ) );
  AN2P U1378 ( .A(n203), .B(n453), .Z(\ab[4][38] ) );
  AN2P U1379 ( .A(n203), .B(n449), .Z(\ab[4][37] ) );
  AN2P U1380 ( .A(n203), .B(n445), .Z(\ab[4][36] ) );
  AN2P U1381 ( .A(n203), .B(n441), .Z(\ab[4][35] ) );
  AN2P U1382 ( .A(n202), .B(n437), .Z(\ab[4][34] ) );
  AN2P U1383 ( .A(n202), .B(n433), .Z(\ab[4][33] ) );
  AN2P U1384 ( .A(n202), .B(n429), .Z(\ab[4][32] ) );
  AN2P U1385 ( .A(n202), .B(n425), .Z(\ab[4][31] ) );
  AN2P U1386 ( .A(n202), .B(n421), .Z(\ab[4][30] ) );
  AN2P U1387 ( .A(n202), .B(n417), .Z(\ab[4][29] ) );
  AN2P U1388 ( .A(n202), .B(n413), .Z(\ab[4][28] ) );
  AN2P U1389 ( .A(n202), .B(n409), .Z(\ab[4][27] ) );
  AN2P U1390 ( .A(n202), .B(n405), .Z(\ab[4][26] ) );
  AN2P U1391 ( .A(n202), .B(n401), .Z(\ab[4][25] ) );
  AN2P U1392 ( .A(n202), .B(n397), .Z(\ab[4][24] ) );
  AN2P U1393 ( .A(n202), .B(n393), .Z(\ab[4][23] ) );
  AN2P U1394 ( .A(n201), .B(n389), .Z(\ab[4][22] ) );
  AN2P U1395 ( .A(n201), .B(n385), .Z(\ab[4][21] ) );
  AN2P U1396 ( .A(n201), .B(n381), .Z(\ab[4][20] ) );
  AN2P U1397 ( .A(n201), .B(n377), .Z(\ab[4][19] ) );
  AN2P U1398 ( .A(n201), .B(n373), .Z(\ab[4][18] ) );
  AN2P U1399 ( .A(n201), .B(n369), .Z(\ab[4][17] ) );
  AN2P U1400 ( .A(n201), .B(n365), .Z(\ab[4][16] ) );
  AN2P U1401 ( .A(n201), .B(n361), .Z(\ab[4][15] ) );
  AN2P U1402 ( .A(n201), .B(n357), .Z(\ab[4][14] ) );
  AN2P U1403 ( .A(n201), .B(n353), .Z(\ab[4][13] ) );
  AN2P U1404 ( .A(n201), .B(n349), .Z(\ab[4][12] ) );
  AN2P U1405 ( .A(n201), .B(n345), .Z(\ab[4][11] ) );
  AN2P U1406 ( .A(n200), .B(n341), .Z(\ab[4][10] ) );
  AN2P U1407 ( .A(n200), .B(n337), .Z(\ab[4][9] ) );
  AN2P U1408 ( .A(n200), .B(n333), .Z(\ab[4][8] ) );
  AN2P U1409 ( .A(n200), .B(n329), .Z(\ab[4][7] ) );
  AN2P U1410 ( .A(n200), .B(n325), .Z(\ab[4][6] ) );
  AN2P U1411 ( .A(n200), .B(n321), .Z(\ab[4][5] ) );
  AN2P U1412 ( .A(n200), .B(n317), .Z(\ab[4][4] ) );
  AN2P U1413 ( .A(n200), .B(n313), .Z(\ab[4][3] ) );
  AN2P U1414 ( .A(n200), .B(n309), .Z(\ab[4][2] ) );
  AN2P U1415 ( .A(n200), .B(n305), .Z(\ab[4][1] ) );
  AN2P U1416 ( .A(n200), .B(n301), .Z(\ab[4][0] ) );
  AN2P U1417 ( .A(n216), .B(n455), .Z(\ab[5][94] ) );
  AN2P U1418 ( .A(n200), .B(n491), .Z(\ab[4][95] ) );
  AN2P U1419 ( .A(n216), .B(n456), .Z(\ab[5][93] ) );
  AN2P U1420 ( .A(n216), .B(n457), .Z(\ab[5][92] ) );
  AN2P U1421 ( .A(n216), .B(n458), .Z(\ab[5][91] ) );
  AN2P U1422 ( .A(n216), .B(n459), .Z(\ab[5][90] ) );
  AN2P U1423 ( .A(n216), .B(n460), .Z(\ab[5][89] ) );
  AN2P U1424 ( .A(n216), .B(n461), .Z(\ab[5][88] ) );
  AN2P U1425 ( .A(n216), .B(n462), .Z(\ab[5][87] ) );
  AN2P U1426 ( .A(n216), .B(n463), .Z(\ab[5][86] ) );
  AN2P U1427 ( .A(n216), .B(n464), .Z(\ab[5][85] ) );
  AN2P U1428 ( .A(n216), .B(n465), .Z(\ab[5][84] ) );
  AN2P U1429 ( .A(n216), .B(n466), .Z(\ab[5][83] ) );
  AN2P U1430 ( .A(n215), .B(n467), .Z(\ab[5][82] ) );
  AN2P U1431 ( .A(n215), .B(n468), .Z(\ab[5][81] ) );
  AN2P U1432 ( .A(n215), .B(n469), .Z(\ab[5][80] ) );
  AN2P U1433 ( .A(n215), .B(n470), .Z(\ab[5][79] ) );
  AN2P U1434 ( .A(n215), .B(n471), .Z(\ab[5][78] ) );
  AN2P U1435 ( .A(n215), .B(n472), .Z(\ab[5][77] ) );
  AN2P U1436 ( .A(n215), .B(n473), .Z(\ab[5][76] ) );
  AN2P U1437 ( .A(n215), .B(n474), .Z(\ab[5][75] ) );
  AN2P U1438 ( .A(n215), .B(n475), .Z(\ab[5][74] ) );
  AN2P U1439 ( .A(n215), .B(n476), .Z(\ab[5][73] ) );
  AN2P U1440 ( .A(n215), .B(n477), .Z(\ab[5][72] ) );
  AN2P U1441 ( .A(n215), .B(n478), .Z(\ab[5][71] ) );
  AN2P U1442 ( .A(n214), .B(n479), .Z(\ab[5][70] ) );
  AN2P U1443 ( .A(n214), .B(n480), .Z(\ab[5][69] ) );
  AN2P U1444 ( .A(n214), .B(n481), .Z(\ab[5][68] ) );
  AN2P U1445 ( .A(n214), .B(n482), .Z(\ab[5][67] ) );
  AN2P U1446 ( .A(n214), .B(n483), .Z(\ab[5][66] ) );
  AN2P U1447 ( .A(n214), .B(n484), .Z(\ab[5][65] ) );
  AN2P U1448 ( .A(n214), .B(n485), .Z(\ab[5][64] ) );
  AN2P U1449 ( .A(n214), .B(n486), .Z(\ab[5][63] ) );
  AN2P U1450 ( .A(n214), .B(n487), .Z(\ab[5][62] ) );
  AN2P U1451 ( .A(n214), .B(n488), .Z(\ab[5][61] ) );
  AN2P U1452 ( .A(n214), .B(n489), .Z(\ab[5][60] ) );
  AN2P U1453 ( .A(n214), .B(B[59]), .Z(\ab[5][59] ) );
  AN2P U1454 ( .A(n213), .B(B[58]), .Z(\ab[5][58] ) );
  AN2P U1455 ( .A(n213), .B(B[57]), .Z(\ab[5][57] ) );
  AN2P U1456 ( .A(n213), .B(B[56]), .Z(\ab[5][56] ) );
  AN2P U1457 ( .A(n213), .B(n490), .Z(\ab[5][55] ) );
  AN2P U1458 ( .A(n213), .B(B[54]), .Z(\ab[5][54] ) );
  AN2P U1459 ( .A(n213), .B(B[53]), .Z(\ab[5][53] ) );
  AN2P U1460 ( .A(n213), .B(B[52]), .Z(\ab[5][52] ) );
  AN2P U1461 ( .A(n213), .B(B[51]), .Z(\ab[5][51] ) );
  AN2P U1462 ( .A(n213), .B(B[50]), .Z(\ab[5][50] ) );
  AN2P U1463 ( .A(n213), .B(B[49]), .Z(\ab[5][49] ) );
  AN2P U1464 ( .A(n213), .B(B[48]), .Z(\ab[5][48] ) );
  AN2P U1465 ( .A(n213), .B(B[47]), .Z(\ab[5][47] ) );
  AN2P U1466 ( .A(n212), .B(B[46]), .Z(\ab[5][46] ) );
  AN2P U1467 ( .A(n212), .B(B[45]), .Z(\ab[5][45] ) );
  AN2P U1468 ( .A(n212), .B(B[44]), .Z(\ab[5][44] ) );
  AN2P U1469 ( .A(n212), .B(B[43]), .Z(\ab[5][43] ) );
  AN2P U1470 ( .A(n212), .B(B[42]), .Z(\ab[5][42] ) );
  AN2P U1471 ( .A(n212), .B(B[41]), .Z(\ab[5][41] ) );
  AN2P U1472 ( .A(n212), .B(B[40]), .Z(\ab[5][40] ) );
  AN2P U1473 ( .A(n212), .B(B[39]), .Z(\ab[5][39] ) );
  AN2P U1474 ( .A(n212), .B(n453), .Z(\ab[5][38] ) );
  AN2P U1475 ( .A(n212), .B(n449), .Z(\ab[5][37] ) );
  AN2P U1476 ( .A(n212), .B(n445), .Z(\ab[5][36] ) );
  AN2P U1477 ( .A(n212), .B(n441), .Z(\ab[5][35] ) );
  AN2P U1478 ( .A(n211), .B(n437), .Z(\ab[5][34] ) );
  AN2P U1479 ( .A(n211), .B(n433), .Z(\ab[5][33] ) );
  AN2P U1480 ( .A(n211), .B(n429), .Z(\ab[5][32] ) );
  AN2P U1481 ( .A(n211), .B(n425), .Z(\ab[5][31] ) );
  AN2P U1482 ( .A(n211), .B(n421), .Z(\ab[5][30] ) );
  AN2P U1483 ( .A(n211), .B(n417), .Z(\ab[5][29] ) );
  AN2P U1484 ( .A(n211), .B(n413), .Z(\ab[5][28] ) );
  AN2P U1485 ( .A(n211), .B(n409), .Z(\ab[5][27] ) );
  AN2P U1486 ( .A(n211), .B(n405), .Z(\ab[5][26] ) );
  AN2P U1487 ( .A(n211), .B(n401), .Z(\ab[5][25] ) );
  AN2P U1488 ( .A(n211), .B(n397), .Z(\ab[5][24] ) );
  AN2P U1489 ( .A(n211), .B(n393), .Z(\ab[5][23] ) );
  AN2P U1490 ( .A(n210), .B(n389), .Z(\ab[5][22] ) );
  AN2P U1491 ( .A(n210), .B(n385), .Z(\ab[5][21] ) );
  AN2P U1492 ( .A(n210), .B(n381), .Z(\ab[5][20] ) );
  AN2P U1493 ( .A(n210), .B(n377), .Z(\ab[5][19] ) );
  AN2P U1494 ( .A(n210), .B(n373), .Z(\ab[5][18] ) );
  AN2P U1495 ( .A(n210), .B(n369), .Z(\ab[5][17] ) );
  AN2P U1496 ( .A(n210), .B(n365), .Z(\ab[5][16] ) );
  AN2P U1497 ( .A(n210), .B(n361), .Z(\ab[5][15] ) );
  AN2P U1498 ( .A(n210), .B(n357), .Z(\ab[5][14] ) );
  AN2P U1499 ( .A(n210), .B(n353), .Z(\ab[5][13] ) );
  AN2P U1500 ( .A(n210), .B(n349), .Z(\ab[5][12] ) );
  AN2P U1501 ( .A(n210), .B(n345), .Z(\ab[5][11] ) );
  AN2P U1502 ( .A(n209), .B(n341), .Z(\ab[5][10] ) );
  AN2P U1503 ( .A(n209), .B(n337), .Z(\ab[5][9] ) );
  AN2P U1504 ( .A(n209), .B(n333), .Z(\ab[5][8] ) );
  AN2P U1505 ( .A(n209), .B(n329), .Z(\ab[5][7] ) );
  AN2P U1506 ( .A(n209), .B(n325), .Z(\ab[5][6] ) );
  AN2P U1507 ( .A(n209), .B(n321), .Z(\ab[5][5] ) );
  AN2P U1508 ( .A(n209), .B(n317), .Z(\ab[5][4] ) );
  AN2P U1509 ( .A(n209), .B(n313), .Z(\ab[5][3] ) );
  AN2P U1510 ( .A(n209), .B(n309), .Z(\ab[5][2] ) );
  AN2P U1511 ( .A(n209), .B(n305), .Z(\ab[5][1] ) );
  AN2P U1512 ( .A(n209), .B(n301), .Z(\ab[5][0] ) );
  AN2P U1513 ( .A(n225), .B(n455), .Z(\ab[6][94] ) );
  AN2P U1514 ( .A(n209), .B(n491), .Z(\ab[5][95] ) );
  AN2P U1515 ( .A(n225), .B(n456), .Z(\ab[6][93] ) );
  AN2P U1516 ( .A(n225), .B(n457), .Z(\ab[6][92] ) );
  AN2P U1517 ( .A(n225), .B(n458), .Z(\ab[6][91] ) );
  AN2P U1518 ( .A(n225), .B(n459), .Z(\ab[6][90] ) );
  AN2P U1519 ( .A(n225), .B(n460), .Z(\ab[6][89] ) );
  AN2P U1520 ( .A(n225), .B(n461), .Z(\ab[6][88] ) );
  AN2P U1521 ( .A(n225), .B(n462), .Z(\ab[6][87] ) );
  AN2P U1522 ( .A(n225), .B(n463), .Z(\ab[6][86] ) );
  AN2P U1523 ( .A(n225), .B(n464), .Z(\ab[6][85] ) );
  AN2P U1524 ( .A(n225), .B(n465), .Z(\ab[6][84] ) );
  AN2P U1525 ( .A(n225), .B(n466), .Z(\ab[6][83] ) );
  AN2P U1526 ( .A(n224), .B(n467), .Z(\ab[6][82] ) );
  AN2P U1527 ( .A(n224), .B(n468), .Z(\ab[6][81] ) );
  AN2P U1528 ( .A(n224), .B(n469), .Z(\ab[6][80] ) );
  AN2P U1529 ( .A(n224), .B(n470), .Z(\ab[6][79] ) );
  AN2P U1530 ( .A(n224), .B(n471), .Z(\ab[6][78] ) );
  AN2P U1531 ( .A(n224), .B(n472), .Z(\ab[6][77] ) );
  AN2P U1532 ( .A(n224), .B(n473), .Z(\ab[6][76] ) );
  AN2P U1533 ( .A(n224), .B(n474), .Z(\ab[6][75] ) );
  AN2P U1534 ( .A(n224), .B(n475), .Z(\ab[6][74] ) );
  AN2P U1535 ( .A(n224), .B(n476), .Z(\ab[6][73] ) );
  AN2P U1536 ( .A(n224), .B(n477), .Z(\ab[6][72] ) );
  AN2P U1537 ( .A(n224), .B(n478), .Z(\ab[6][71] ) );
  AN2P U1538 ( .A(n223), .B(n479), .Z(\ab[6][70] ) );
  AN2P U1539 ( .A(n223), .B(n480), .Z(\ab[6][69] ) );
  AN2P U1540 ( .A(n223), .B(n481), .Z(\ab[6][68] ) );
  AN2P U1541 ( .A(n223), .B(n482), .Z(\ab[6][67] ) );
  AN2P U1542 ( .A(n223), .B(n483), .Z(\ab[6][66] ) );
  AN2P U1543 ( .A(n223), .B(n484), .Z(\ab[6][65] ) );
  AN2P U1544 ( .A(n223), .B(n485), .Z(\ab[6][64] ) );
  AN2P U1545 ( .A(n223), .B(n486), .Z(\ab[6][63] ) );
  AN2P U1546 ( .A(n223), .B(n487), .Z(\ab[6][62] ) );
  AN2P U1547 ( .A(n223), .B(n488), .Z(\ab[6][61] ) );
  AN2P U1548 ( .A(n223), .B(n489), .Z(\ab[6][60] ) );
  AN2P U1549 ( .A(n223), .B(B[59]), .Z(\ab[6][59] ) );
  AN2P U1550 ( .A(n222), .B(B[58]), .Z(\ab[6][58] ) );
  AN2P U1551 ( .A(n222), .B(B[57]), .Z(\ab[6][57] ) );
  AN2P U1552 ( .A(n222), .B(B[56]), .Z(\ab[6][56] ) );
  AN2P U1553 ( .A(n222), .B(n490), .Z(\ab[6][55] ) );
  AN2P U1554 ( .A(n222), .B(B[54]), .Z(\ab[6][54] ) );
  AN2P U1555 ( .A(n222), .B(B[53]), .Z(\ab[6][53] ) );
  AN2P U1556 ( .A(n222), .B(B[52]), .Z(\ab[6][52] ) );
  AN2P U1557 ( .A(n222), .B(B[51]), .Z(\ab[6][51] ) );
  AN2P U1558 ( .A(n222), .B(B[50]), .Z(\ab[6][50] ) );
  AN2P U1559 ( .A(n222), .B(B[49]), .Z(\ab[6][49] ) );
  AN2P U1560 ( .A(n222), .B(B[48]), .Z(\ab[6][48] ) );
  AN2P U1561 ( .A(n222), .B(B[47]), .Z(\ab[6][47] ) );
  AN2P U1562 ( .A(n221), .B(B[46]), .Z(\ab[6][46] ) );
  AN2P U1563 ( .A(n221), .B(B[45]), .Z(\ab[6][45] ) );
  AN2P U1564 ( .A(n221), .B(B[44]), .Z(\ab[6][44] ) );
  AN2P U1565 ( .A(n221), .B(B[43]), .Z(\ab[6][43] ) );
  AN2P U1566 ( .A(n221), .B(B[42]), .Z(\ab[6][42] ) );
  AN2P U1567 ( .A(n221), .B(B[41]), .Z(\ab[6][41] ) );
  AN2P U1568 ( .A(n221), .B(B[40]), .Z(\ab[6][40] ) );
  AN2P U1569 ( .A(n221), .B(B[39]), .Z(\ab[6][39] ) );
  AN2P U1570 ( .A(n221), .B(n452), .Z(\ab[6][38] ) );
  AN2P U1571 ( .A(n221), .B(n448), .Z(\ab[6][37] ) );
  AN2P U1572 ( .A(n221), .B(n444), .Z(\ab[6][36] ) );
  AN2P U1573 ( .A(n221), .B(n440), .Z(\ab[6][35] ) );
  AN2P U1574 ( .A(n220), .B(n436), .Z(\ab[6][34] ) );
  AN2P U1575 ( .A(n220), .B(n432), .Z(\ab[6][33] ) );
  AN2P U1576 ( .A(n220), .B(n428), .Z(\ab[6][32] ) );
  AN2P U1577 ( .A(n220), .B(n424), .Z(\ab[6][31] ) );
  AN2P U1578 ( .A(n220), .B(n420), .Z(\ab[6][30] ) );
  AN2P U1579 ( .A(n220), .B(n416), .Z(\ab[6][29] ) );
  AN2P U1580 ( .A(n220), .B(n412), .Z(\ab[6][28] ) );
  AN2P U1581 ( .A(n220), .B(n408), .Z(\ab[6][27] ) );
  AN2P U1582 ( .A(n220), .B(n404), .Z(\ab[6][26] ) );
  AN2P U1583 ( .A(n220), .B(n400), .Z(\ab[6][25] ) );
  AN2P U1584 ( .A(n220), .B(n396), .Z(\ab[6][24] ) );
  AN2P U1585 ( .A(n220), .B(n392), .Z(\ab[6][23] ) );
  AN2P U1586 ( .A(n219), .B(n388), .Z(\ab[6][22] ) );
  AN2P U1587 ( .A(n219), .B(n384), .Z(\ab[6][21] ) );
  AN2P U1588 ( .A(n219), .B(n380), .Z(\ab[6][20] ) );
  AN2P U1589 ( .A(n219), .B(n376), .Z(\ab[6][19] ) );
  AN2P U1590 ( .A(n219), .B(n372), .Z(\ab[6][18] ) );
  AN2P U1591 ( .A(n219), .B(n368), .Z(\ab[6][17] ) );
  AN2P U1592 ( .A(n219), .B(n364), .Z(\ab[6][16] ) );
  AN2P U1593 ( .A(n219), .B(n360), .Z(\ab[6][15] ) );
  AN2P U1594 ( .A(n219), .B(n356), .Z(\ab[6][14] ) );
  AN2P U1595 ( .A(n219), .B(n352), .Z(\ab[6][13] ) );
  AN2P U1596 ( .A(n219), .B(n348), .Z(\ab[6][12] ) );
  AN2P U1597 ( .A(n219), .B(n344), .Z(\ab[6][11] ) );
  AN2P U1598 ( .A(n218), .B(n340), .Z(\ab[6][10] ) );
  AN2P U1599 ( .A(n218), .B(n336), .Z(\ab[6][9] ) );
  AN2P U1600 ( .A(n218), .B(n332), .Z(\ab[6][8] ) );
  AN2P U1601 ( .A(n218), .B(n328), .Z(\ab[6][7] ) );
  AN2P U1602 ( .A(n218), .B(n324), .Z(\ab[6][6] ) );
  AN2P U1603 ( .A(n218), .B(n320), .Z(\ab[6][5] ) );
  AN2P U1604 ( .A(n218), .B(n316), .Z(\ab[6][4] ) );
  AN2P U1605 ( .A(n218), .B(n312), .Z(\ab[6][3] ) );
  AN2P U1606 ( .A(n218), .B(n308), .Z(\ab[6][2] ) );
  AN2P U1607 ( .A(n218), .B(n304), .Z(\ab[6][1] ) );
  AN2P U1608 ( .A(n218), .B(n300), .Z(\ab[6][0] ) );
  AN2P U1609 ( .A(n234), .B(n455), .Z(\ab[7][94] ) );
  AN2P U1610 ( .A(n218), .B(n491), .Z(\ab[6][95] ) );
  AN2P U1611 ( .A(n234), .B(n456), .Z(\ab[7][93] ) );
  AN2P U1612 ( .A(n234), .B(n457), .Z(\ab[7][92] ) );
  AN2P U1613 ( .A(n234), .B(n458), .Z(\ab[7][91] ) );
  AN2P U1614 ( .A(n234), .B(n459), .Z(\ab[7][90] ) );
  AN2P U1615 ( .A(n234), .B(n460), .Z(\ab[7][89] ) );
  AN2P U1616 ( .A(n234), .B(n461), .Z(\ab[7][88] ) );
  AN2P U1617 ( .A(n234), .B(n462), .Z(\ab[7][87] ) );
  AN2P U1618 ( .A(n234), .B(n463), .Z(\ab[7][86] ) );
  AN2P U1619 ( .A(n234), .B(n464), .Z(\ab[7][85] ) );
  AN2P U1620 ( .A(n234), .B(n465), .Z(\ab[7][84] ) );
  AN2P U1621 ( .A(n234), .B(n466), .Z(\ab[7][83] ) );
  AN2P U1622 ( .A(n233), .B(n467), .Z(\ab[7][82] ) );
  AN2P U1623 ( .A(n233), .B(n468), .Z(\ab[7][81] ) );
  AN2P U1624 ( .A(n233), .B(n469), .Z(\ab[7][80] ) );
  AN2P U1625 ( .A(n233), .B(n470), .Z(\ab[7][79] ) );
  AN2P U1626 ( .A(n233), .B(n471), .Z(\ab[7][78] ) );
  AN2P U1627 ( .A(n233), .B(n472), .Z(\ab[7][77] ) );
  AN2P U1628 ( .A(n233), .B(n473), .Z(\ab[7][76] ) );
  AN2P U1629 ( .A(n233), .B(n474), .Z(\ab[7][75] ) );
  AN2P U1630 ( .A(n233), .B(n475), .Z(\ab[7][74] ) );
  AN2P U1631 ( .A(n233), .B(n476), .Z(\ab[7][73] ) );
  AN2P U1632 ( .A(n233), .B(n477), .Z(\ab[7][72] ) );
  AN2P U1633 ( .A(n233), .B(n478), .Z(\ab[7][71] ) );
  AN2P U1634 ( .A(n232), .B(n479), .Z(\ab[7][70] ) );
  AN2P U1635 ( .A(n232), .B(n480), .Z(\ab[7][69] ) );
  AN2P U1636 ( .A(n232), .B(n481), .Z(\ab[7][68] ) );
  AN2P U1637 ( .A(n232), .B(n482), .Z(\ab[7][67] ) );
  AN2P U1638 ( .A(n232), .B(n483), .Z(\ab[7][66] ) );
  AN2P U1639 ( .A(n232), .B(n484), .Z(\ab[7][65] ) );
  AN2P U1640 ( .A(n232), .B(n485), .Z(\ab[7][64] ) );
  AN2P U1641 ( .A(n232), .B(n486), .Z(\ab[7][63] ) );
  AN2P U1642 ( .A(n232), .B(n487), .Z(\ab[7][62] ) );
  AN2P U1643 ( .A(n232), .B(n488), .Z(\ab[7][61] ) );
  AN2P U1644 ( .A(n232), .B(n489), .Z(\ab[7][60] ) );
  AN2P U1645 ( .A(n232), .B(B[59]), .Z(\ab[7][59] ) );
  AN2P U1646 ( .A(n231), .B(B[58]), .Z(\ab[7][58] ) );
  AN2P U1647 ( .A(n231), .B(B[57]), .Z(\ab[7][57] ) );
  AN2P U1648 ( .A(n231), .B(B[56]), .Z(\ab[7][56] ) );
  AN2P U1649 ( .A(n231), .B(n490), .Z(\ab[7][55] ) );
  AN2P U1650 ( .A(n231), .B(B[54]), .Z(\ab[7][54] ) );
  AN2P U1651 ( .A(n231), .B(B[53]), .Z(\ab[7][53] ) );
  AN2P U1652 ( .A(n231), .B(B[52]), .Z(\ab[7][52] ) );
  AN2P U1653 ( .A(n231), .B(B[51]), .Z(\ab[7][51] ) );
  AN2P U1654 ( .A(n231), .B(B[50]), .Z(\ab[7][50] ) );
  AN2P U1655 ( .A(n231), .B(B[49]), .Z(\ab[7][49] ) );
  AN2P U1656 ( .A(n231), .B(B[48]), .Z(\ab[7][48] ) );
  AN2P U1657 ( .A(n231), .B(B[47]), .Z(\ab[7][47] ) );
  AN2P U1658 ( .A(n230), .B(B[46]), .Z(\ab[7][46] ) );
  AN2P U1659 ( .A(n230), .B(B[45]), .Z(\ab[7][45] ) );
  AN2P U1660 ( .A(n230), .B(B[44]), .Z(\ab[7][44] ) );
  AN2P U1661 ( .A(n230), .B(B[43]), .Z(\ab[7][43] ) );
  AN2P U1662 ( .A(n230), .B(B[42]), .Z(\ab[7][42] ) );
  AN2P U1663 ( .A(n230), .B(B[41]), .Z(\ab[7][41] ) );
  AN2P U1664 ( .A(n230), .B(B[40]), .Z(\ab[7][40] ) );
  AN2P U1665 ( .A(n230), .B(B[39]), .Z(\ab[7][39] ) );
  AN2P U1666 ( .A(n230), .B(n452), .Z(\ab[7][38] ) );
  AN2P U1667 ( .A(n230), .B(n448), .Z(\ab[7][37] ) );
  AN2P U1668 ( .A(n230), .B(n444), .Z(\ab[7][36] ) );
  AN2P U1669 ( .A(n230), .B(n440), .Z(\ab[7][35] ) );
  AN2P U1670 ( .A(n229), .B(n436), .Z(\ab[7][34] ) );
  AN2P U1671 ( .A(n229), .B(n432), .Z(\ab[7][33] ) );
  AN2P U1672 ( .A(n229), .B(n428), .Z(\ab[7][32] ) );
  AN2P U1673 ( .A(n229), .B(n424), .Z(\ab[7][31] ) );
  AN2P U1674 ( .A(n229), .B(n420), .Z(\ab[7][30] ) );
  AN2P U1675 ( .A(n229), .B(n416), .Z(\ab[7][29] ) );
  AN2P U1676 ( .A(n229), .B(n412), .Z(\ab[7][28] ) );
  AN2P U1677 ( .A(n229), .B(n408), .Z(\ab[7][27] ) );
  AN2P U1678 ( .A(n229), .B(n404), .Z(\ab[7][26] ) );
  AN2P U1679 ( .A(n229), .B(n400), .Z(\ab[7][25] ) );
  AN2P U1680 ( .A(n229), .B(n396), .Z(\ab[7][24] ) );
  AN2P U1681 ( .A(n229), .B(n392), .Z(\ab[7][23] ) );
  AN2P U1682 ( .A(n228), .B(n388), .Z(\ab[7][22] ) );
  AN2P U1683 ( .A(n228), .B(n384), .Z(\ab[7][21] ) );
  AN2P U1684 ( .A(n228), .B(n380), .Z(\ab[7][20] ) );
  AN2P U1685 ( .A(n228), .B(n376), .Z(\ab[7][19] ) );
  AN2P U1686 ( .A(n228), .B(n372), .Z(\ab[7][18] ) );
  AN2P U1687 ( .A(n228), .B(n368), .Z(\ab[7][17] ) );
  AN2P U1688 ( .A(n228), .B(n364), .Z(\ab[7][16] ) );
  AN2P U1689 ( .A(n228), .B(n360), .Z(\ab[7][15] ) );
  AN2P U1690 ( .A(n228), .B(n356), .Z(\ab[7][14] ) );
  AN2P U1691 ( .A(n228), .B(n352), .Z(\ab[7][13] ) );
  AN2P U1692 ( .A(n228), .B(n348), .Z(\ab[7][12] ) );
  AN2P U1693 ( .A(n228), .B(n344), .Z(\ab[7][11] ) );
  AN2P U1694 ( .A(n227), .B(n340), .Z(\ab[7][10] ) );
  AN2P U1695 ( .A(n227), .B(n336), .Z(\ab[7][9] ) );
  AN2P U1696 ( .A(n227), .B(n332), .Z(\ab[7][8] ) );
  AN2P U1697 ( .A(n227), .B(n328), .Z(\ab[7][7] ) );
  AN2P U1698 ( .A(n227), .B(n324), .Z(\ab[7][6] ) );
  AN2P U1699 ( .A(n227), .B(n320), .Z(\ab[7][5] ) );
  AN2P U1700 ( .A(n227), .B(n316), .Z(\ab[7][4] ) );
  AN2P U1701 ( .A(n227), .B(n312), .Z(\ab[7][3] ) );
  AN2P U1702 ( .A(n227), .B(n308), .Z(\ab[7][2] ) );
  AN2P U1703 ( .A(n227), .B(n304), .Z(\ab[7][1] ) );
  AN2P U1704 ( .A(n227), .B(n300), .Z(\ab[7][0] ) );
  AN2P U1705 ( .A(n243), .B(n455), .Z(\ab[8][94] ) );
  AN2P U1706 ( .A(n227), .B(n491), .Z(\ab[7][95] ) );
  AN2P U1707 ( .A(n243), .B(n456), .Z(\ab[8][93] ) );
  AN2P U1708 ( .A(n243), .B(n457), .Z(\ab[8][92] ) );
  AN2P U1709 ( .A(n243), .B(n458), .Z(\ab[8][91] ) );
  AN2P U1710 ( .A(n243), .B(n459), .Z(\ab[8][90] ) );
  AN2P U1711 ( .A(n243), .B(n460), .Z(\ab[8][89] ) );
  AN2P U1712 ( .A(n243), .B(n461), .Z(\ab[8][88] ) );
  AN2P U1713 ( .A(n243), .B(n462), .Z(\ab[8][87] ) );
  AN2P U1714 ( .A(n243), .B(n463), .Z(\ab[8][86] ) );
  AN2P U1715 ( .A(n243), .B(n464), .Z(\ab[8][85] ) );
  AN2P U1716 ( .A(n243), .B(n465), .Z(\ab[8][84] ) );
  AN2P U1717 ( .A(n243), .B(n466), .Z(\ab[8][83] ) );
  AN2P U1718 ( .A(n242), .B(n467), .Z(\ab[8][82] ) );
  AN2P U1719 ( .A(n242), .B(n468), .Z(\ab[8][81] ) );
  AN2P U1720 ( .A(n242), .B(n469), .Z(\ab[8][80] ) );
  AN2P U1721 ( .A(n242), .B(n470), .Z(\ab[8][79] ) );
  AN2P U1722 ( .A(n242), .B(n471), .Z(\ab[8][78] ) );
  AN2P U1723 ( .A(n242), .B(n472), .Z(\ab[8][77] ) );
  AN2P U1724 ( .A(n242), .B(n473), .Z(\ab[8][76] ) );
  AN2P U1725 ( .A(n242), .B(n474), .Z(\ab[8][75] ) );
  AN2P U1726 ( .A(n242), .B(n475), .Z(\ab[8][74] ) );
  AN2P U1727 ( .A(n242), .B(n476), .Z(\ab[8][73] ) );
  AN2P U1728 ( .A(n242), .B(n477), .Z(\ab[8][72] ) );
  AN2P U1729 ( .A(n242), .B(n478), .Z(\ab[8][71] ) );
  AN2P U1730 ( .A(n241), .B(n479), .Z(\ab[8][70] ) );
  AN2P U1731 ( .A(n241), .B(n480), .Z(\ab[8][69] ) );
  AN2P U1732 ( .A(n241), .B(n481), .Z(\ab[8][68] ) );
  AN2P U1733 ( .A(n241), .B(n482), .Z(\ab[8][67] ) );
  AN2P U1734 ( .A(n241), .B(n483), .Z(\ab[8][66] ) );
  AN2P U1735 ( .A(n241), .B(n484), .Z(\ab[8][65] ) );
  AN2P U1736 ( .A(n241), .B(n485), .Z(\ab[8][64] ) );
  AN2P U1737 ( .A(n241), .B(n486), .Z(\ab[8][63] ) );
  AN2P U1738 ( .A(n241), .B(n487), .Z(\ab[8][62] ) );
  AN2P U1739 ( .A(n241), .B(n488), .Z(\ab[8][61] ) );
  AN2P U1740 ( .A(n241), .B(n489), .Z(\ab[8][60] ) );
  AN2P U1741 ( .A(n241), .B(B[59]), .Z(\ab[8][59] ) );
  AN2P U1742 ( .A(n240), .B(B[58]), .Z(\ab[8][58] ) );
  AN2P U1743 ( .A(n240), .B(B[57]), .Z(\ab[8][57] ) );
  AN2P U1744 ( .A(n240), .B(B[56]), .Z(\ab[8][56] ) );
  AN2P U1745 ( .A(n240), .B(n490), .Z(\ab[8][55] ) );
  AN2P U1746 ( .A(n240), .B(B[54]), .Z(\ab[8][54] ) );
  AN2P U1747 ( .A(n240), .B(B[53]), .Z(\ab[8][53] ) );
  AN2P U1748 ( .A(n240), .B(B[52]), .Z(\ab[8][52] ) );
  AN2P U1749 ( .A(n240), .B(B[51]), .Z(\ab[8][51] ) );
  AN2P U1750 ( .A(n240), .B(B[50]), .Z(\ab[8][50] ) );
  AN2P U1751 ( .A(n240), .B(B[49]), .Z(\ab[8][49] ) );
  AN2P U1752 ( .A(n240), .B(B[48]), .Z(\ab[8][48] ) );
  AN2P U1753 ( .A(n240), .B(B[47]), .Z(\ab[8][47] ) );
  AN2P U1754 ( .A(n239), .B(B[46]), .Z(\ab[8][46] ) );
  AN2P U1755 ( .A(n239), .B(B[45]), .Z(\ab[8][45] ) );
  AN2P U1756 ( .A(n239), .B(B[44]), .Z(\ab[8][44] ) );
  AN2P U1757 ( .A(n239), .B(B[43]), .Z(\ab[8][43] ) );
  AN2P U1758 ( .A(n239), .B(B[42]), .Z(\ab[8][42] ) );
  AN2P U1759 ( .A(n239), .B(B[41]), .Z(\ab[8][41] ) );
  AN2P U1760 ( .A(n239), .B(B[40]), .Z(\ab[8][40] ) );
  AN2P U1761 ( .A(n239), .B(B[39]), .Z(\ab[8][39] ) );
  AN2P U1762 ( .A(n239), .B(n452), .Z(\ab[8][38] ) );
  AN2P U1763 ( .A(n239), .B(n448), .Z(\ab[8][37] ) );
  AN2P U1764 ( .A(n239), .B(n444), .Z(\ab[8][36] ) );
  AN2P U1765 ( .A(n239), .B(n440), .Z(\ab[8][35] ) );
  AN2P U1766 ( .A(n238), .B(n436), .Z(\ab[8][34] ) );
  AN2P U1767 ( .A(n238), .B(n432), .Z(\ab[8][33] ) );
  AN2P U1768 ( .A(n238), .B(n428), .Z(\ab[8][32] ) );
  AN2P U1769 ( .A(n238), .B(n424), .Z(\ab[8][31] ) );
  AN2P U1770 ( .A(n238), .B(n420), .Z(\ab[8][30] ) );
  AN2P U1771 ( .A(n238), .B(n416), .Z(\ab[8][29] ) );
  AN2P U1772 ( .A(n238), .B(n412), .Z(\ab[8][28] ) );
  AN2P U1773 ( .A(n238), .B(n408), .Z(\ab[8][27] ) );
  AN2P U1774 ( .A(n238), .B(n404), .Z(\ab[8][26] ) );
  AN2P U1775 ( .A(n238), .B(n400), .Z(\ab[8][25] ) );
  AN2P U1776 ( .A(n238), .B(n396), .Z(\ab[8][24] ) );
  AN2P U1777 ( .A(n238), .B(n392), .Z(\ab[8][23] ) );
  AN2P U1778 ( .A(n237), .B(n388), .Z(\ab[8][22] ) );
  AN2P U1779 ( .A(n237), .B(n384), .Z(\ab[8][21] ) );
  AN2P U1780 ( .A(n237), .B(n380), .Z(\ab[8][20] ) );
  AN2P U1781 ( .A(n237), .B(n376), .Z(\ab[8][19] ) );
  AN2P U1782 ( .A(n237), .B(n372), .Z(\ab[8][18] ) );
  AN2P U1783 ( .A(n237), .B(n368), .Z(\ab[8][17] ) );
  AN2P U1784 ( .A(n237), .B(n364), .Z(\ab[8][16] ) );
  AN2P U1785 ( .A(n237), .B(n360), .Z(\ab[8][15] ) );
  AN2P U1786 ( .A(n237), .B(n356), .Z(\ab[8][14] ) );
  AN2P U1787 ( .A(n237), .B(n352), .Z(\ab[8][13] ) );
  AN2P U1788 ( .A(n237), .B(n348), .Z(\ab[8][12] ) );
  AN2P U1789 ( .A(n237), .B(n344), .Z(\ab[8][11] ) );
  AN2P U1790 ( .A(n236), .B(n340), .Z(\ab[8][10] ) );
  AN2P U1791 ( .A(n236), .B(n336), .Z(\ab[8][9] ) );
  AN2P U1792 ( .A(n236), .B(n332), .Z(\ab[8][8] ) );
  AN2P U1793 ( .A(n236), .B(n328), .Z(\ab[8][7] ) );
  AN2P U1794 ( .A(n236), .B(n324), .Z(\ab[8][6] ) );
  AN2P U1795 ( .A(n236), .B(n320), .Z(\ab[8][5] ) );
  AN2P U1796 ( .A(n236), .B(n316), .Z(\ab[8][4] ) );
  AN2P U1797 ( .A(n236), .B(n312), .Z(\ab[8][3] ) );
  AN2P U1798 ( .A(n236), .B(n308), .Z(\ab[8][2] ) );
  AN2P U1799 ( .A(n236), .B(n304), .Z(\ab[8][1] ) );
  AN2P U1800 ( .A(n236), .B(n300), .Z(\ab[8][0] ) );
  AN2P U1801 ( .A(n252), .B(n455), .Z(\ab[9][94] ) );
  AN2P U1802 ( .A(n236), .B(n491), .Z(\ab[8][95] ) );
  AN2P U1803 ( .A(n252), .B(n456), .Z(\ab[9][93] ) );
  AN2P U1804 ( .A(n252), .B(n457), .Z(\ab[9][92] ) );
  AN2P U1805 ( .A(n252), .B(n458), .Z(\ab[9][91] ) );
  AN2P U1806 ( .A(n252), .B(n459), .Z(\ab[9][90] ) );
  AN2P U1807 ( .A(n252), .B(n460), .Z(\ab[9][89] ) );
  AN2P U1808 ( .A(n252), .B(n461), .Z(\ab[9][88] ) );
  AN2P U1809 ( .A(n252), .B(n462), .Z(\ab[9][87] ) );
  AN2P U1810 ( .A(n252), .B(n463), .Z(\ab[9][86] ) );
  AN2P U1811 ( .A(n252), .B(n464), .Z(\ab[9][85] ) );
  AN2P U1812 ( .A(n252), .B(n465), .Z(\ab[9][84] ) );
  AN2P U1813 ( .A(n252), .B(n466), .Z(\ab[9][83] ) );
  AN2P U1814 ( .A(n251), .B(n467), .Z(\ab[9][82] ) );
  AN2P U1815 ( .A(n251), .B(n468), .Z(\ab[9][81] ) );
  AN2P U1816 ( .A(n251), .B(n469), .Z(\ab[9][80] ) );
  AN2P U1817 ( .A(n251), .B(n470), .Z(\ab[9][79] ) );
  AN2P U1818 ( .A(n251), .B(n471), .Z(\ab[9][78] ) );
  AN2P U1819 ( .A(n251), .B(n472), .Z(\ab[9][77] ) );
  AN2P U1820 ( .A(n251), .B(n473), .Z(\ab[9][76] ) );
  AN2P U1821 ( .A(n251), .B(n474), .Z(\ab[9][75] ) );
  AN2P U1822 ( .A(n251), .B(n475), .Z(\ab[9][74] ) );
  AN2P U1823 ( .A(n251), .B(n476), .Z(\ab[9][73] ) );
  AN2P U1824 ( .A(n251), .B(n477), .Z(\ab[9][72] ) );
  AN2P U1825 ( .A(n251), .B(n478), .Z(\ab[9][71] ) );
  AN2P U1826 ( .A(n250), .B(n479), .Z(\ab[9][70] ) );
  AN2P U1827 ( .A(n250), .B(n480), .Z(\ab[9][69] ) );
  AN2P U1828 ( .A(n250), .B(n481), .Z(\ab[9][68] ) );
  AN2P U1829 ( .A(n250), .B(n482), .Z(\ab[9][67] ) );
  AN2P U1830 ( .A(n250), .B(n483), .Z(\ab[9][66] ) );
  AN2P U1831 ( .A(n250), .B(n484), .Z(\ab[9][65] ) );
  AN2P U1832 ( .A(n250), .B(n485), .Z(\ab[9][64] ) );
  AN2P U1833 ( .A(n250), .B(n486), .Z(\ab[9][63] ) );
  AN2P U1834 ( .A(n250), .B(n487), .Z(\ab[9][62] ) );
  AN2P U1835 ( .A(n250), .B(n488), .Z(\ab[9][61] ) );
  AN2P U1836 ( .A(n250), .B(n489), .Z(\ab[9][60] ) );
  AN2P U1837 ( .A(n250), .B(B[59]), .Z(\ab[9][59] ) );
  AN2P U1838 ( .A(n249), .B(B[58]), .Z(\ab[9][58] ) );
  AN2P U1839 ( .A(n249), .B(B[57]), .Z(\ab[9][57] ) );
  AN2P U1840 ( .A(n249), .B(B[56]), .Z(\ab[9][56] ) );
  AN2P U1841 ( .A(n249), .B(n490), .Z(\ab[9][55] ) );
  AN2P U1842 ( .A(n249), .B(B[54]), .Z(\ab[9][54] ) );
  AN2P U1843 ( .A(n249), .B(B[53]), .Z(\ab[9][53] ) );
  AN2P U1844 ( .A(n249), .B(B[52]), .Z(\ab[9][52] ) );
  AN2P U1845 ( .A(n249), .B(B[51]), .Z(\ab[9][51] ) );
  AN2P U1846 ( .A(n249), .B(B[50]), .Z(\ab[9][50] ) );
  AN2P U1847 ( .A(n249), .B(B[49]), .Z(\ab[9][49] ) );
  AN2P U1848 ( .A(n249), .B(B[48]), .Z(\ab[9][48] ) );
  AN2P U1849 ( .A(n249), .B(B[47]), .Z(\ab[9][47] ) );
  AN2P U1850 ( .A(n248), .B(B[46]), .Z(\ab[9][46] ) );
  AN2P U1851 ( .A(n248), .B(B[45]), .Z(\ab[9][45] ) );
  AN2P U1852 ( .A(n248), .B(B[44]), .Z(\ab[9][44] ) );
  AN2P U1853 ( .A(n248), .B(B[43]), .Z(\ab[9][43] ) );
  AN2P U1854 ( .A(n248), .B(B[42]), .Z(\ab[9][42] ) );
  AN2P U1855 ( .A(n248), .B(B[41]), .Z(\ab[9][41] ) );
  AN2P U1856 ( .A(n248), .B(B[40]), .Z(\ab[9][40] ) );
  AN2P U1857 ( .A(n248), .B(B[39]), .Z(\ab[9][39] ) );
  AN2P U1858 ( .A(n248), .B(n452), .Z(\ab[9][38] ) );
  AN2P U1859 ( .A(n248), .B(n448), .Z(\ab[9][37] ) );
  AN2P U1860 ( .A(n248), .B(n444), .Z(\ab[9][36] ) );
  AN2P U1861 ( .A(n248), .B(n440), .Z(\ab[9][35] ) );
  AN2P U1862 ( .A(n247), .B(n436), .Z(\ab[9][34] ) );
  AN2P U1863 ( .A(n247), .B(n432), .Z(\ab[9][33] ) );
  AN2P U1864 ( .A(n247), .B(n428), .Z(\ab[9][32] ) );
  AN2P U1865 ( .A(n247), .B(n424), .Z(\ab[9][31] ) );
  AN2P U1866 ( .A(n247), .B(n420), .Z(\ab[9][30] ) );
  AN2P U1867 ( .A(n247), .B(n416), .Z(\ab[9][29] ) );
  AN2P U1868 ( .A(n247), .B(n412), .Z(\ab[9][28] ) );
  AN2P U1869 ( .A(n247), .B(n408), .Z(\ab[9][27] ) );
  AN2P U1870 ( .A(n247), .B(n404), .Z(\ab[9][26] ) );
  AN2P U1871 ( .A(n247), .B(n400), .Z(\ab[9][25] ) );
  AN2P U1872 ( .A(n247), .B(n396), .Z(\ab[9][24] ) );
  AN2P U1873 ( .A(n247), .B(n392), .Z(\ab[9][23] ) );
  AN2P U1874 ( .A(n246), .B(n388), .Z(\ab[9][22] ) );
  AN2P U1875 ( .A(n246), .B(n384), .Z(\ab[9][21] ) );
  AN2P U1876 ( .A(n246), .B(n380), .Z(\ab[9][20] ) );
  AN2P U1877 ( .A(n246), .B(n376), .Z(\ab[9][19] ) );
  AN2P U1878 ( .A(n246), .B(n372), .Z(\ab[9][18] ) );
  AN2P U1879 ( .A(n246), .B(n368), .Z(\ab[9][17] ) );
  AN2P U1880 ( .A(n246), .B(n364), .Z(\ab[9][16] ) );
  AN2P U1881 ( .A(n246), .B(n360), .Z(\ab[9][15] ) );
  AN2P U1882 ( .A(n246), .B(n356), .Z(\ab[9][14] ) );
  AN2P U1883 ( .A(n246), .B(n352), .Z(\ab[9][13] ) );
  AN2P U1884 ( .A(n246), .B(n348), .Z(\ab[9][12] ) );
  AN2P U1885 ( .A(n246), .B(n344), .Z(\ab[9][11] ) );
  AN2P U1886 ( .A(n245), .B(n340), .Z(\ab[9][10] ) );
  AN2P U1887 ( .A(n245), .B(n336), .Z(\ab[9][9] ) );
  AN2P U1888 ( .A(n245), .B(n332), .Z(\ab[9][8] ) );
  AN2P U1889 ( .A(n245), .B(n328), .Z(\ab[9][7] ) );
  AN2P U1890 ( .A(n245), .B(n324), .Z(\ab[9][6] ) );
  AN2P U1891 ( .A(n245), .B(n320), .Z(\ab[9][5] ) );
  AN2P U1892 ( .A(n245), .B(n316), .Z(\ab[9][4] ) );
  AN2P U1893 ( .A(n245), .B(n312), .Z(\ab[9][3] ) );
  AN2P U1894 ( .A(n245), .B(n308), .Z(\ab[9][2] ) );
  AN2P U1895 ( .A(n245), .B(n304), .Z(\ab[9][1] ) );
  AN2P U1896 ( .A(n245), .B(n300), .Z(\ab[9][0] ) );
  AN2P U1897 ( .A(n261), .B(n455), .Z(\ab[10][94] ) );
  AN2P U1898 ( .A(n245), .B(n491), .Z(\ab[9][95] ) );
  AN2P U1899 ( .A(n261), .B(n456), .Z(\ab[10][93] ) );
  AN2P U1900 ( .A(n261), .B(n457), .Z(\ab[10][92] ) );
  AN2P U1901 ( .A(n261), .B(n458), .Z(\ab[10][91] ) );
  AN2P U1902 ( .A(n261), .B(n459), .Z(\ab[10][90] ) );
  AN2P U1903 ( .A(n261), .B(n460), .Z(\ab[10][89] ) );
  AN2P U1904 ( .A(n261), .B(n461), .Z(\ab[10][88] ) );
  AN2P U1905 ( .A(n261), .B(n462), .Z(\ab[10][87] ) );
  AN2P U1906 ( .A(n261), .B(n463), .Z(\ab[10][86] ) );
  AN2P U1907 ( .A(n261), .B(n464), .Z(\ab[10][85] ) );
  AN2P U1908 ( .A(n261), .B(n465), .Z(\ab[10][84] ) );
  AN2P U1909 ( .A(n261), .B(n466), .Z(\ab[10][83] ) );
  AN2P U1910 ( .A(n260), .B(n467), .Z(\ab[10][82] ) );
  AN2P U1911 ( .A(n260), .B(n468), .Z(\ab[10][81] ) );
  AN2P U1912 ( .A(n260), .B(n469), .Z(\ab[10][80] ) );
  AN2P U1913 ( .A(n260), .B(n470), .Z(\ab[10][79] ) );
  AN2P U1914 ( .A(n260), .B(n471), .Z(\ab[10][78] ) );
  AN2P U1915 ( .A(n260), .B(n472), .Z(\ab[10][77] ) );
  AN2P U1916 ( .A(n260), .B(n473), .Z(\ab[10][76] ) );
  AN2P U1917 ( .A(n260), .B(n474), .Z(\ab[10][75] ) );
  AN2P U1918 ( .A(n260), .B(n475), .Z(\ab[10][74] ) );
  AN2P U1919 ( .A(n260), .B(n476), .Z(\ab[10][73] ) );
  AN2P U1920 ( .A(n260), .B(n477), .Z(\ab[10][72] ) );
  AN2P U1921 ( .A(n260), .B(n478), .Z(\ab[10][71] ) );
  AN2P U1922 ( .A(n259), .B(n479), .Z(\ab[10][70] ) );
  AN2P U1923 ( .A(n259), .B(n480), .Z(\ab[10][69] ) );
  AN2P U1924 ( .A(n259), .B(n481), .Z(\ab[10][68] ) );
  AN2P U1925 ( .A(n259), .B(n482), .Z(\ab[10][67] ) );
  AN2P U1926 ( .A(n259), .B(n483), .Z(\ab[10][66] ) );
  AN2P U1927 ( .A(n259), .B(n484), .Z(\ab[10][65] ) );
  AN2P U1928 ( .A(n259), .B(n485), .Z(\ab[10][64] ) );
  AN2P U1929 ( .A(n259), .B(n486), .Z(\ab[10][63] ) );
  AN2P U1930 ( .A(n259), .B(n487), .Z(\ab[10][62] ) );
  AN2P U1931 ( .A(n259), .B(n488), .Z(\ab[10][61] ) );
  AN2P U1932 ( .A(n259), .B(n489), .Z(\ab[10][60] ) );
  AN2P U1933 ( .A(n259), .B(B[59]), .Z(\ab[10][59] ) );
  AN2P U1934 ( .A(n258), .B(B[58]), .Z(\ab[10][58] ) );
  AN2P U1935 ( .A(n258), .B(B[57]), .Z(\ab[10][57] ) );
  AN2P U1936 ( .A(n258), .B(B[56]), .Z(\ab[10][56] ) );
  AN2P U1937 ( .A(n258), .B(n490), .Z(\ab[10][55] ) );
  AN2P U1938 ( .A(n258), .B(B[54]), .Z(\ab[10][54] ) );
  AN2P U1939 ( .A(n258), .B(B[53]), .Z(\ab[10][53] ) );
  AN2P U1940 ( .A(n258), .B(B[52]), .Z(\ab[10][52] ) );
  AN2P U1941 ( .A(n258), .B(B[51]), .Z(\ab[10][51] ) );
  AN2P U1942 ( .A(n258), .B(B[50]), .Z(\ab[10][50] ) );
  AN2P U1943 ( .A(n258), .B(B[49]), .Z(\ab[10][49] ) );
  AN2P U1944 ( .A(n258), .B(B[48]), .Z(\ab[10][48] ) );
  AN2P U1945 ( .A(n258), .B(B[47]), .Z(\ab[10][47] ) );
  AN2P U1946 ( .A(n257), .B(B[46]), .Z(\ab[10][46] ) );
  AN2P U1947 ( .A(n257), .B(B[45]), .Z(\ab[10][45] ) );
  AN2P U1948 ( .A(n257), .B(B[44]), .Z(\ab[10][44] ) );
  AN2P U1949 ( .A(n257), .B(B[43]), .Z(\ab[10][43] ) );
  AN2P U1950 ( .A(n257), .B(B[42]), .Z(\ab[10][42] ) );
  AN2P U1951 ( .A(n257), .B(B[41]), .Z(\ab[10][41] ) );
  AN2P U1952 ( .A(n257), .B(B[40]), .Z(\ab[10][40] ) );
  AN2P U1953 ( .A(n257), .B(B[39]), .Z(\ab[10][39] ) );
  AN2P U1954 ( .A(n257), .B(n452), .Z(\ab[10][38] ) );
  AN2P U1955 ( .A(n257), .B(n448), .Z(\ab[10][37] ) );
  AN2P U1956 ( .A(n257), .B(n444), .Z(\ab[10][36] ) );
  AN2P U1957 ( .A(n257), .B(n440), .Z(\ab[10][35] ) );
  AN2P U1958 ( .A(n256), .B(n436), .Z(\ab[10][34] ) );
  AN2P U1959 ( .A(n256), .B(n432), .Z(\ab[10][33] ) );
  AN2P U1960 ( .A(n256), .B(n428), .Z(\ab[10][32] ) );
  AN2P U1961 ( .A(n256), .B(n424), .Z(\ab[10][31] ) );
  AN2P U1962 ( .A(n256), .B(n420), .Z(\ab[10][30] ) );
  AN2P U1963 ( .A(n256), .B(n416), .Z(\ab[10][29] ) );
  AN2P U1964 ( .A(n256), .B(n412), .Z(\ab[10][28] ) );
  AN2P U1965 ( .A(n256), .B(n408), .Z(\ab[10][27] ) );
  AN2P U1966 ( .A(n256), .B(n404), .Z(\ab[10][26] ) );
  AN2P U1967 ( .A(n256), .B(n400), .Z(\ab[10][25] ) );
  AN2P U1968 ( .A(n256), .B(n396), .Z(\ab[10][24] ) );
  AN2P U1969 ( .A(n256), .B(n392), .Z(\ab[10][23] ) );
  AN2P U1970 ( .A(n255), .B(n388), .Z(\ab[10][22] ) );
  AN2P U1971 ( .A(n255), .B(n384), .Z(\ab[10][21] ) );
  AN2P U1972 ( .A(n255), .B(n380), .Z(\ab[10][20] ) );
  AN2P U1973 ( .A(n255), .B(n376), .Z(\ab[10][19] ) );
  AN2P U1974 ( .A(n255), .B(n372), .Z(\ab[10][18] ) );
  AN2P U1975 ( .A(n255), .B(n368), .Z(\ab[10][17] ) );
  AN2P U1976 ( .A(n255), .B(n364), .Z(\ab[10][16] ) );
  AN2P U1977 ( .A(n255), .B(n360), .Z(\ab[10][15] ) );
  AN2P U1978 ( .A(n255), .B(n356), .Z(\ab[10][14] ) );
  AN2P U1979 ( .A(n255), .B(n352), .Z(\ab[10][13] ) );
  AN2P U1980 ( .A(n255), .B(n348), .Z(\ab[10][12] ) );
  AN2P U1981 ( .A(n255), .B(n344), .Z(\ab[10][11] ) );
  AN2P U1982 ( .A(n254), .B(n340), .Z(\ab[10][10] ) );
  AN2P U1983 ( .A(n254), .B(n336), .Z(\ab[10][9] ) );
  AN2P U1984 ( .A(n254), .B(n332), .Z(\ab[10][8] ) );
  AN2P U1985 ( .A(n254), .B(n328), .Z(\ab[10][7] ) );
  AN2P U1986 ( .A(n254), .B(n324), .Z(\ab[10][6] ) );
  AN2P U1987 ( .A(n254), .B(n320), .Z(\ab[10][5] ) );
  AN2P U1988 ( .A(n254), .B(n316), .Z(\ab[10][4] ) );
  AN2P U1989 ( .A(n254), .B(n312), .Z(\ab[10][3] ) );
  AN2P U1990 ( .A(n254), .B(n308), .Z(\ab[10][2] ) );
  AN2P U1991 ( .A(n254), .B(n304), .Z(\ab[10][1] ) );
  AN2P U1992 ( .A(n254), .B(n300), .Z(\ab[10][0] ) );
  AN2P U1993 ( .A(n270), .B(n455), .Z(\ab[11][94] ) );
  AN2P U1994 ( .A(n254), .B(n491), .Z(\ab[10][95] ) );
  AN2P U1995 ( .A(n270), .B(n456), .Z(\ab[11][93] ) );
  AN2P U1996 ( .A(n270), .B(n457), .Z(\ab[11][92] ) );
  AN2P U1997 ( .A(n270), .B(n458), .Z(\ab[11][91] ) );
  AN2P U1998 ( .A(n270), .B(n459), .Z(\ab[11][90] ) );
  AN2P U1999 ( .A(n270), .B(n460), .Z(\ab[11][89] ) );
  AN2P U2000 ( .A(n270), .B(n461), .Z(\ab[11][88] ) );
  AN2P U2001 ( .A(n270), .B(n462), .Z(\ab[11][87] ) );
  AN2P U2002 ( .A(n270), .B(n463), .Z(\ab[11][86] ) );
  AN2P U2003 ( .A(n270), .B(n464), .Z(\ab[11][85] ) );
  AN2P U2004 ( .A(n270), .B(n465), .Z(\ab[11][84] ) );
  AN2P U2005 ( .A(n270), .B(n466), .Z(\ab[11][83] ) );
  AN2P U2006 ( .A(n269), .B(n467), .Z(\ab[11][82] ) );
  AN2P U2007 ( .A(n269), .B(n468), .Z(\ab[11][81] ) );
  AN2P U2008 ( .A(n269), .B(n469), .Z(\ab[11][80] ) );
  AN2P U2009 ( .A(n269), .B(n470), .Z(\ab[11][79] ) );
  AN2P U2010 ( .A(n269), .B(n471), .Z(\ab[11][78] ) );
  AN2P U2011 ( .A(n269), .B(n472), .Z(\ab[11][77] ) );
  AN2P U2012 ( .A(n269), .B(n473), .Z(\ab[11][76] ) );
  AN2P U2013 ( .A(n269), .B(n474), .Z(\ab[11][75] ) );
  AN2P U2014 ( .A(n269), .B(n475), .Z(\ab[11][74] ) );
  AN2P U2015 ( .A(n269), .B(n476), .Z(\ab[11][73] ) );
  AN2P U2016 ( .A(n269), .B(n477), .Z(\ab[11][72] ) );
  AN2P U2017 ( .A(n269), .B(n478), .Z(\ab[11][71] ) );
  AN2P U2018 ( .A(n268), .B(n479), .Z(\ab[11][70] ) );
  AN2P U2019 ( .A(n268), .B(n480), .Z(\ab[11][69] ) );
  AN2P U2020 ( .A(n268), .B(n481), .Z(\ab[11][68] ) );
  AN2P U2021 ( .A(n268), .B(n482), .Z(\ab[11][67] ) );
  AN2P U2022 ( .A(n268), .B(n483), .Z(\ab[11][66] ) );
  AN2P U2023 ( .A(n268), .B(n484), .Z(\ab[11][65] ) );
  AN2P U2024 ( .A(n268), .B(n485), .Z(\ab[11][64] ) );
  AN2P U2025 ( .A(n268), .B(n486), .Z(\ab[11][63] ) );
  AN2P U2026 ( .A(n268), .B(n487), .Z(\ab[11][62] ) );
  AN2P U2027 ( .A(n268), .B(n488), .Z(\ab[11][61] ) );
  AN2P U2028 ( .A(n268), .B(n489), .Z(\ab[11][60] ) );
  AN2P U2029 ( .A(n268), .B(B[59]), .Z(\ab[11][59] ) );
  AN2P U2030 ( .A(n267), .B(B[58]), .Z(\ab[11][58] ) );
  AN2P U2031 ( .A(n267), .B(B[57]), .Z(\ab[11][57] ) );
  AN2P U2032 ( .A(n267), .B(B[56]), .Z(\ab[11][56] ) );
  AN2P U2033 ( .A(n267), .B(n490), .Z(\ab[11][55] ) );
  AN2P U2034 ( .A(n267), .B(B[54]), .Z(\ab[11][54] ) );
  AN2P U2035 ( .A(n267), .B(B[53]), .Z(\ab[11][53] ) );
  AN2P U2036 ( .A(n267), .B(B[52]), .Z(\ab[11][52] ) );
  AN2P U2037 ( .A(n267), .B(B[51]), .Z(\ab[11][51] ) );
  AN2P U2038 ( .A(n267), .B(B[50]), .Z(\ab[11][50] ) );
  AN2P U2039 ( .A(n267), .B(B[49]), .Z(\ab[11][49] ) );
  AN2P U2040 ( .A(n267), .B(B[48]), .Z(\ab[11][48] ) );
  AN2P U2041 ( .A(n267), .B(B[47]), .Z(\ab[11][47] ) );
  AN2P U2042 ( .A(n266), .B(B[46]), .Z(\ab[11][46] ) );
  AN2P U2043 ( .A(n266), .B(B[45]), .Z(\ab[11][45] ) );
  AN2P U2044 ( .A(n266), .B(B[44]), .Z(\ab[11][44] ) );
  AN2P U2045 ( .A(n266), .B(B[43]), .Z(\ab[11][43] ) );
  AN2P U2046 ( .A(n266), .B(B[42]), .Z(\ab[11][42] ) );
  AN2P U2047 ( .A(n266), .B(B[41]), .Z(\ab[11][41] ) );
  AN2P U2048 ( .A(n266), .B(B[40]), .Z(\ab[11][40] ) );
  AN2P U2049 ( .A(n266), .B(B[39]), .Z(\ab[11][39] ) );
  AN2P U2050 ( .A(n266), .B(n452), .Z(\ab[11][38] ) );
  AN2P U2051 ( .A(n266), .B(n448), .Z(\ab[11][37] ) );
  AN2P U2052 ( .A(n266), .B(n444), .Z(\ab[11][36] ) );
  AN2P U2053 ( .A(n266), .B(n440), .Z(\ab[11][35] ) );
  AN2P U2054 ( .A(n265), .B(n436), .Z(\ab[11][34] ) );
  AN2P U2055 ( .A(n265), .B(n432), .Z(\ab[11][33] ) );
  AN2P U2056 ( .A(n265), .B(n428), .Z(\ab[11][32] ) );
  AN2P U2057 ( .A(n265), .B(n424), .Z(\ab[11][31] ) );
  AN2P U2058 ( .A(n265), .B(n420), .Z(\ab[11][30] ) );
  AN2P U2059 ( .A(n265), .B(n416), .Z(\ab[11][29] ) );
  AN2P U2060 ( .A(n265), .B(n412), .Z(\ab[11][28] ) );
  AN2P U2061 ( .A(n265), .B(n408), .Z(\ab[11][27] ) );
  AN2P U2062 ( .A(n265), .B(n404), .Z(\ab[11][26] ) );
  AN2P U2063 ( .A(n265), .B(n400), .Z(\ab[11][25] ) );
  AN2P U2064 ( .A(n265), .B(n396), .Z(\ab[11][24] ) );
  AN2P U2065 ( .A(n265), .B(n392), .Z(\ab[11][23] ) );
  AN2P U2066 ( .A(n264), .B(n388), .Z(\ab[11][22] ) );
  AN2P U2067 ( .A(n264), .B(n384), .Z(\ab[11][21] ) );
  AN2P U2068 ( .A(n264), .B(n380), .Z(\ab[11][20] ) );
  AN2P U2069 ( .A(n264), .B(n376), .Z(\ab[11][19] ) );
  AN2P U2070 ( .A(n264), .B(n372), .Z(\ab[11][18] ) );
  AN2P U2071 ( .A(n264), .B(n368), .Z(\ab[11][17] ) );
  AN2P U2072 ( .A(n264), .B(n364), .Z(\ab[11][16] ) );
  AN2P U2073 ( .A(n264), .B(n360), .Z(\ab[11][15] ) );
  AN2P U2074 ( .A(n264), .B(n356), .Z(\ab[11][14] ) );
  AN2P U2075 ( .A(n264), .B(n352), .Z(\ab[11][13] ) );
  AN2P U2076 ( .A(n264), .B(n348), .Z(\ab[11][12] ) );
  AN2P U2077 ( .A(n264), .B(n344), .Z(\ab[11][11] ) );
  AN2P U2078 ( .A(n263), .B(n340), .Z(\ab[11][10] ) );
  AN2P U2079 ( .A(n263), .B(n336), .Z(\ab[11][9] ) );
  AN2P U2080 ( .A(n263), .B(n332), .Z(\ab[11][8] ) );
  AN2P U2081 ( .A(n263), .B(n328), .Z(\ab[11][7] ) );
  AN2P U2082 ( .A(n263), .B(n324), .Z(\ab[11][6] ) );
  AN2P U2083 ( .A(n263), .B(n320), .Z(\ab[11][5] ) );
  AN2P U2084 ( .A(n263), .B(n316), .Z(\ab[11][4] ) );
  AN2P U2085 ( .A(n263), .B(n312), .Z(\ab[11][3] ) );
  AN2P U2086 ( .A(n263), .B(n308), .Z(\ab[11][2] ) );
  AN2P U2087 ( .A(n263), .B(n304), .Z(\ab[11][1] ) );
  AN2P U2088 ( .A(n263), .B(n300), .Z(\ab[11][0] ) );
  AN2P U2089 ( .A(n279), .B(n455), .Z(\ab[12][94] ) );
  AN2P U2090 ( .A(n263), .B(n491), .Z(\ab[11][95] ) );
  AN2P U2091 ( .A(n279), .B(n456), .Z(\ab[12][93] ) );
  AN2P U2092 ( .A(n279), .B(n457), .Z(\ab[12][92] ) );
  AN2P U2093 ( .A(n279), .B(n458), .Z(\ab[12][91] ) );
  AN2P U2094 ( .A(n279), .B(n459), .Z(\ab[12][90] ) );
  AN2P U2095 ( .A(n279), .B(n460), .Z(\ab[12][89] ) );
  AN2P U2096 ( .A(n279), .B(n461), .Z(\ab[12][88] ) );
  AN2P U2097 ( .A(n279), .B(n462), .Z(\ab[12][87] ) );
  AN2P U2098 ( .A(n279), .B(n463), .Z(\ab[12][86] ) );
  AN2P U2099 ( .A(n279), .B(n464), .Z(\ab[12][85] ) );
  AN2P U2100 ( .A(n279), .B(n465), .Z(\ab[12][84] ) );
  AN2P U2101 ( .A(n279), .B(n466), .Z(\ab[12][83] ) );
  AN2P U2102 ( .A(n278), .B(n467), .Z(\ab[12][82] ) );
  AN2P U2103 ( .A(n278), .B(n468), .Z(\ab[12][81] ) );
  AN2P U2104 ( .A(n278), .B(n469), .Z(\ab[12][80] ) );
  AN2P U2105 ( .A(n278), .B(n470), .Z(\ab[12][79] ) );
  AN2P U2106 ( .A(n278), .B(n471), .Z(\ab[12][78] ) );
  AN2P U2107 ( .A(n278), .B(n472), .Z(\ab[12][77] ) );
  AN2P U2108 ( .A(n278), .B(n473), .Z(\ab[12][76] ) );
  AN2P U2109 ( .A(n278), .B(n474), .Z(\ab[12][75] ) );
  AN2P U2110 ( .A(n278), .B(n475), .Z(\ab[12][74] ) );
  AN2P U2111 ( .A(n278), .B(n476), .Z(\ab[12][73] ) );
  AN2P U2112 ( .A(n278), .B(n477), .Z(\ab[12][72] ) );
  AN2P U2113 ( .A(n278), .B(n478), .Z(\ab[12][71] ) );
  AN2P U2114 ( .A(n277), .B(n479), .Z(\ab[12][70] ) );
  AN2P U2115 ( .A(n277), .B(n480), .Z(\ab[12][69] ) );
  AN2P U2116 ( .A(n277), .B(n481), .Z(\ab[12][68] ) );
  AN2P U2117 ( .A(n277), .B(n482), .Z(\ab[12][67] ) );
  AN2P U2118 ( .A(n277), .B(n483), .Z(\ab[12][66] ) );
  AN2P U2119 ( .A(n277), .B(n484), .Z(\ab[12][65] ) );
  AN2P U2120 ( .A(n277), .B(n485), .Z(\ab[12][64] ) );
  AN2P U2121 ( .A(n277), .B(n486), .Z(\ab[12][63] ) );
  AN2P U2122 ( .A(n277), .B(n487), .Z(\ab[12][62] ) );
  AN2P U2123 ( .A(n277), .B(n488), .Z(\ab[12][61] ) );
  AN2P U2124 ( .A(n277), .B(n489), .Z(\ab[12][60] ) );
  AN2P U2125 ( .A(n277), .B(B[59]), .Z(\ab[12][59] ) );
  AN2P U2126 ( .A(n276), .B(B[58]), .Z(\ab[12][58] ) );
  AN2P U2127 ( .A(n276), .B(B[57]), .Z(\ab[12][57] ) );
  AN2P U2128 ( .A(n276), .B(B[56]), .Z(\ab[12][56] ) );
  AN2P U2129 ( .A(n276), .B(n490), .Z(\ab[12][55] ) );
  AN2P U2130 ( .A(n276), .B(B[54]), .Z(\ab[12][54] ) );
  AN2P U2131 ( .A(n276), .B(B[53]), .Z(\ab[12][53] ) );
  AN2P U2132 ( .A(n276), .B(B[52]), .Z(\ab[12][52] ) );
  AN2P U2133 ( .A(n276), .B(B[51]), .Z(\ab[12][51] ) );
  AN2P U2134 ( .A(n276), .B(B[50]), .Z(\ab[12][50] ) );
  AN2P U2135 ( .A(n276), .B(B[49]), .Z(\ab[12][49] ) );
  AN2P U2136 ( .A(n276), .B(B[48]), .Z(\ab[12][48] ) );
  AN2P U2137 ( .A(n276), .B(B[47]), .Z(\ab[12][47] ) );
  AN2P U2138 ( .A(n275), .B(B[46]), .Z(\ab[12][46] ) );
  AN2P U2139 ( .A(n275), .B(B[45]), .Z(\ab[12][45] ) );
  AN2P U2140 ( .A(n275), .B(B[44]), .Z(\ab[12][44] ) );
  AN2P U2141 ( .A(n275), .B(B[43]), .Z(\ab[12][43] ) );
  AN2P U2142 ( .A(n275), .B(B[42]), .Z(\ab[12][42] ) );
  AN2P U2143 ( .A(n275), .B(B[41]), .Z(\ab[12][41] ) );
  AN2P U2144 ( .A(n275), .B(B[40]), .Z(\ab[12][40] ) );
  AN2P U2145 ( .A(n275), .B(B[39]), .Z(\ab[12][39] ) );
  AN2P U2146 ( .A(n275), .B(n452), .Z(\ab[12][38] ) );
  AN2P U2147 ( .A(n275), .B(n448), .Z(\ab[12][37] ) );
  AN2P U2148 ( .A(n275), .B(n444), .Z(\ab[12][36] ) );
  AN2P U2149 ( .A(n275), .B(n440), .Z(\ab[12][35] ) );
  AN2P U2150 ( .A(n274), .B(n436), .Z(\ab[12][34] ) );
  AN2P U2151 ( .A(n274), .B(n432), .Z(\ab[12][33] ) );
  AN2P U2152 ( .A(n274), .B(n428), .Z(\ab[12][32] ) );
  AN2P U2153 ( .A(n274), .B(n424), .Z(\ab[12][31] ) );
  AN2P U2154 ( .A(n274), .B(n420), .Z(\ab[12][30] ) );
  AN2P U2155 ( .A(n274), .B(n416), .Z(\ab[12][29] ) );
  AN2P U2156 ( .A(n274), .B(n412), .Z(\ab[12][28] ) );
  AN2P U2157 ( .A(n274), .B(n408), .Z(\ab[12][27] ) );
  AN2P U2158 ( .A(n274), .B(n404), .Z(\ab[12][26] ) );
  AN2P U2159 ( .A(n274), .B(n400), .Z(\ab[12][25] ) );
  AN2P U2160 ( .A(n274), .B(n396), .Z(\ab[12][24] ) );
  AN2P U2161 ( .A(n274), .B(n392), .Z(\ab[12][23] ) );
  AN2P U2162 ( .A(n273), .B(n388), .Z(\ab[12][22] ) );
  AN2P U2163 ( .A(n273), .B(n384), .Z(\ab[12][21] ) );
  AN2P U2164 ( .A(n273), .B(n380), .Z(\ab[12][20] ) );
  AN2P U2165 ( .A(n273), .B(n376), .Z(\ab[12][19] ) );
  AN2P U2166 ( .A(n273), .B(n372), .Z(\ab[12][18] ) );
  AN2P U2167 ( .A(n273), .B(n368), .Z(\ab[12][17] ) );
  AN2P U2168 ( .A(n273), .B(n364), .Z(\ab[12][16] ) );
  AN2P U2169 ( .A(n273), .B(n360), .Z(\ab[12][15] ) );
  AN2P U2170 ( .A(n273), .B(n356), .Z(\ab[12][14] ) );
  AN2P U2171 ( .A(n273), .B(n352), .Z(\ab[12][13] ) );
  AN2P U2172 ( .A(n273), .B(n348), .Z(\ab[12][12] ) );
  AN2P U2173 ( .A(n273), .B(n344), .Z(\ab[12][11] ) );
  AN2P U2174 ( .A(n272), .B(n340), .Z(\ab[12][10] ) );
  AN2P U2175 ( .A(n272), .B(n336), .Z(\ab[12][9] ) );
  AN2P U2176 ( .A(n272), .B(n332), .Z(\ab[12][8] ) );
  AN2P U2177 ( .A(n272), .B(n328), .Z(\ab[12][7] ) );
  AN2P U2178 ( .A(n272), .B(n324), .Z(\ab[12][6] ) );
  AN2P U2179 ( .A(n272), .B(n320), .Z(\ab[12][5] ) );
  AN2P U2180 ( .A(n272), .B(n316), .Z(\ab[12][4] ) );
  AN2P U2181 ( .A(n272), .B(n312), .Z(\ab[12][3] ) );
  AN2P U2182 ( .A(n272), .B(n308), .Z(\ab[12][2] ) );
  AN2P U2183 ( .A(n272), .B(n304), .Z(\ab[12][1] ) );
  AN2P U2184 ( .A(n272), .B(n300), .Z(\ab[12][0] ) );
  AN2P U2185 ( .A(n288), .B(n455), .Z(\ab[13][94] ) );
  AN2P U2186 ( .A(n272), .B(n491), .Z(\ab[12][95] ) );
  AN2P U2187 ( .A(n288), .B(n456), .Z(\ab[13][93] ) );
  AN2P U2188 ( .A(n288), .B(n457), .Z(\ab[13][92] ) );
  AN2P U2189 ( .A(n288), .B(n458), .Z(\ab[13][91] ) );
  AN2P U2190 ( .A(n288), .B(n459), .Z(\ab[13][90] ) );
  AN2P U2191 ( .A(n288), .B(n460), .Z(\ab[13][89] ) );
  AN2P U2192 ( .A(n288), .B(n461), .Z(\ab[13][88] ) );
  AN2P U2193 ( .A(n288), .B(n462), .Z(\ab[13][87] ) );
  AN2P U2194 ( .A(n288), .B(n463), .Z(\ab[13][86] ) );
  AN2P U2195 ( .A(n288), .B(n464), .Z(\ab[13][85] ) );
  AN2P U2196 ( .A(n288), .B(n465), .Z(\ab[13][84] ) );
  AN2P U2197 ( .A(n288), .B(n466), .Z(\ab[13][83] ) );
  AN2P U2198 ( .A(n287), .B(n467), .Z(\ab[13][82] ) );
  AN2P U2199 ( .A(n287), .B(n468), .Z(\ab[13][81] ) );
  AN2P U2200 ( .A(n287), .B(n469), .Z(\ab[13][80] ) );
  AN2P U2201 ( .A(n287), .B(n470), .Z(\ab[13][79] ) );
  AN2P U2202 ( .A(n287), .B(n471), .Z(\ab[13][78] ) );
  AN2P U2203 ( .A(n287), .B(n472), .Z(\ab[13][77] ) );
  AN2P U2204 ( .A(n287), .B(n473), .Z(\ab[13][76] ) );
  AN2P U2205 ( .A(n287), .B(n474), .Z(\ab[13][75] ) );
  AN2P U2206 ( .A(n287), .B(n475), .Z(\ab[13][74] ) );
  AN2P U2207 ( .A(n287), .B(n476), .Z(\ab[13][73] ) );
  AN2P U2208 ( .A(n287), .B(n477), .Z(\ab[13][72] ) );
  AN2P U2209 ( .A(n287), .B(n478), .Z(\ab[13][71] ) );
  AN2P U2210 ( .A(n286), .B(n479), .Z(\ab[13][70] ) );
  AN2P U2211 ( .A(n286), .B(n480), .Z(\ab[13][69] ) );
  AN2P U2212 ( .A(n286), .B(n481), .Z(\ab[13][68] ) );
  AN2P U2213 ( .A(n286), .B(n482), .Z(\ab[13][67] ) );
  AN2P U2214 ( .A(n286), .B(n483), .Z(\ab[13][66] ) );
  AN2P U2215 ( .A(n286), .B(n484), .Z(\ab[13][65] ) );
  AN2P U2216 ( .A(n286), .B(n485), .Z(\ab[13][64] ) );
  AN2P U2217 ( .A(n286), .B(n486), .Z(\ab[13][63] ) );
  AN2P U2218 ( .A(n286), .B(n487), .Z(\ab[13][62] ) );
  AN2P U2219 ( .A(n286), .B(n488), .Z(\ab[13][61] ) );
  AN2P U2220 ( .A(n286), .B(n489), .Z(\ab[13][60] ) );
  AN2P U2221 ( .A(n286), .B(B[59]), .Z(\ab[13][59] ) );
  AN2P U2222 ( .A(n285), .B(B[58]), .Z(\ab[13][58] ) );
  AN2P U2223 ( .A(n285), .B(B[57]), .Z(\ab[13][57] ) );
  AN2P U2224 ( .A(n285), .B(B[56]), .Z(\ab[13][56] ) );
  AN2P U2225 ( .A(n285), .B(n490), .Z(\ab[13][55] ) );
  AN2P U2226 ( .A(n285), .B(B[54]), .Z(\ab[13][54] ) );
  AN2P U2227 ( .A(n285), .B(B[53]), .Z(\ab[13][53] ) );
  AN2P U2228 ( .A(n285), .B(B[52]), .Z(\ab[13][52] ) );
  AN2P U2229 ( .A(n285), .B(B[51]), .Z(\ab[13][51] ) );
  AN2P U2230 ( .A(n285), .B(B[50]), .Z(\ab[13][50] ) );
  AN2P U2231 ( .A(n285), .B(B[49]), .Z(\ab[13][49] ) );
  AN2P U2232 ( .A(n285), .B(B[48]), .Z(\ab[13][48] ) );
  AN2P U2233 ( .A(n285), .B(B[47]), .Z(\ab[13][47] ) );
  AN2P U2234 ( .A(n284), .B(B[46]), .Z(\ab[13][46] ) );
  AN2P U2235 ( .A(n284), .B(B[45]), .Z(\ab[13][45] ) );
  AN2P U2236 ( .A(n284), .B(B[44]), .Z(\ab[13][44] ) );
  AN2P U2237 ( .A(n284), .B(B[43]), .Z(\ab[13][43] ) );
  AN2P U2238 ( .A(n284), .B(B[42]), .Z(\ab[13][42] ) );
  AN2P U2239 ( .A(n284), .B(B[41]), .Z(\ab[13][41] ) );
  AN2P U2240 ( .A(n284), .B(B[40]), .Z(\ab[13][40] ) );
  AN2P U2241 ( .A(n284), .B(B[39]), .Z(\ab[13][39] ) );
  AN2P U2242 ( .A(n284), .B(n452), .Z(\ab[13][38] ) );
  AN2P U2243 ( .A(n284), .B(n448), .Z(\ab[13][37] ) );
  AN2P U2244 ( .A(n284), .B(n444), .Z(\ab[13][36] ) );
  AN2P U2245 ( .A(n284), .B(n440), .Z(\ab[13][35] ) );
  AN2P U2246 ( .A(n283), .B(n436), .Z(\ab[13][34] ) );
  AN2P U2247 ( .A(n283), .B(n432), .Z(\ab[13][33] ) );
  AN2P U2248 ( .A(n283), .B(n428), .Z(\ab[13][32] ) );
  AN2P U2249 ( .A(n283), .B(n424), .Z(\ab[13][31] ) );
  AN2P U2250 ( .A(n283), .B(n420), .Z(\ab[13][30] ) );
  AN2P U2251 ( .A(n283), .B(n416), .Z(\ab[13][29] ) );
  AN2P U2252 ( .A(n283), .B(n412), .Z(\ab[13][28] ) );
  AN2P U2253 ( .A(n283), .B(n408), .Z(\ab[13][27] ) );
  AN2P U2254 ( .A(n283), .B(n404), .Z(\ab[13][26] ) );
  AN2P U2255 ( .A(n283), .B(n400), .Z(\ab[13][25] ) );
  AN2P U2256 ( .A(n283), .B(n396), .Z(\ab[13][24] ) );
  AN2P U2257 ( .A(n283), .B(n392), .Z(\ab[13][23] ) );
  AN2P U2258 ( .A(n282), .B(n388), .Z(\ab[13][22] ) );
  AN2P U2259 ( .A(n282), .B(n384), .Z(\ab[13][21] ) );
  AN2P U2260 ( .A(n282), .B(n380), .Z(\ab[13][20] ) );
  AN2P U2261 ( .A(n282), .B(n376), .Z(\ab[13][19] ) );
  AN2P U2262 ( .A(n282), .B(n372), .Z(\ab[13][18] ) );
  AN2P U2263 ( .A(n282), .B(n368), .Z(\ab[13][17] ) );
  AN2P U2264 ( .A(n282), .B(n364), .Z(\ab[13][16] ) );
  AN2P U2265 ( .A(n282), .B(n360), .Z(\ab[13][15] ) );
  AN2P U2266 ( .A(n282), .B(n356), .Z(\ab[13][14] ) );
  AN2P U2267 ( .A(n282), .B(n352), .Z(\ab[13][13] ) );
  AN2P U2268 ( .A(n282), .B(n348), .Z(\ab[13][12] ) );
  AN2P U2269 ( .A(n282), .B(n344), .Z(\ab[13][11] ) );
  AN2P U2270 ( .A(n281), .B(n340), .Z(\ab[13][10] ) );
  AN2P U2271 ( .A(n281), .B(n336), .Z(\ab[13][9] ) );
  AN2P U2272 ( .A(n281), .B(n332), .Z(\ab[13][8] ) );
  AN2P U2273 ( .A(n281), .B(n328), .Z(\ab[13][7] ) );
  AN2P U2274 ( .A(n281), .B(n324), .Z(\ab[13][6] ) );
  AN2P U2275 ( .A(n281), .B(n320), .Z(\ab[13][5] ) );
  AN2P U2276 ( .A(n281), .B(n316), .Z(\ab[13][4] ) );
  AN2P U2277 ( .A(n281), .B(n312), .Z(\ab[13][3] ) );
  AN2P U2278 ( .A(n281), .B(n308), .Z(\ab[13][2] ) );
  AN2P U2279 ( .A(n281), .B(n304), .Z(\ab[13][1] ) );
  AN2P U2280 ( .A(n281), .B(n300), .Z(\ab[13][0] ) );
  AN2P U2281 ( .A(n297), .B(n455), .Z(\ab[14][94] ) );
  AN2P U2282 ( .A(n281), .B(n491), .Z(\ab[13][95] ) );
  AN2P U2283 ( .A(n297), .B(n456), .Z(\ab[14][93] ) );
  AN2P U2284 ( .A(n297), .B(n457), .Z(\ab[14][92] ) );
  AN2P U2285 ( .A(n297), .B(n458), .Z(\ab[14][91] ) );
  AN2P U2286 ( .A(n297), .B(n459), .Z(\ab[14][90] ) );
  AN2P U2287 ( .A(n297), .B(n460), .Z(\ab[14][89] ) );
  AN2P U2288 ( .A(n297), .B(n461), .Z(\ab[14][88] ) );
  AN2P U2289 ( .A(n297), .B(n462), .Z(\ab[14][87] ) );
  AN2P U2290 ( .A(n297), .B(n463), .Z(\ab[14][86] ) );
  AN2P U2291 ( .A(n297), .B(n464), .Z(\ab[14][85] ) );
  AN2P U2292 ( .A(n297), .B(n465), .Z(\ab[14][84] ) );
  AN2P U2293 ( .A(n297), .B(n466), .Z(\ab[14][83] ) );
  AN2P U2294 ( .A(n296), .B(n467), .Z(\ab[14][82] ) );
  AN2P U2295 ( .A(n296), .B(n468), .Z(\ab[14][81] ) );
  AN2P U2296 ( .A(n296), .B(n469), .Z(\ab[14][80] ) );
  AN2P U2297 ( .A(n296), .B(n470), .Z(\ab[14][79] ) );
  AN2P U2298 ( .A(n296), .B(n471), .Z(\ab[14][78] ) );
  AN2P U2299 ( .A(n296), .B(n472), .Z(\ab[14][77] ) );
  AN2P U2300 ( .A(n296), .B(n473), .Z(\ab[14][76] ) );
  AN2P U2301 ( .A(n296), .B(n474), .Z(\ab[14][75] ) );
  AN2P U2302 ( .A(n296), .B(n475), .Z(\ab[14][74] ) );
  AN2P U2303 ( .A(n296), .B(n476), .Z(\ab[14][73] ) );
  AN2P U2304 ( .A(n296), .B(n477), .Z(\ab[14][72] ) );
  AN2P U2305 ( .A(n296), .B(n478), .Z(\ab[14][71] ) );
  AN2P U2306 ( .A(n295), .B(n479), .Z(\ab[14][70] ) );
  AN2P U2307 ( .A(n295), .B(n480), .Z(\ab[14][69] ) );
  AN2P U2308 ( .A(n295), .B(n481), .Z(\ab[14][68] ) );
  AN2P U2309 ( .A(n295), .B(n482), .Z(\ab[14][67] ) );
  AN2P U2310 ( .A(n295), .B(n483), .Z(\ab[14][66] ) );
  AN2P U2311 ( .A(n295), .B(n484), .Z(\ab[14][65] ) );
  AN2P U2312 ( .A(n295), .B(n485), .Z(\ab[14][64] ) );
  AN2P U2313 ( .A(n295), .B(n486), .Z(\ab[14][63] ) );
  AN2P U2314 ( .A(n295), .B(n487), .Z(\ab[14][62] ) );
  AN2P U2315 ( .A(n295), .B(n488), .Z(\ab[14][61] ) );
  AN2P U2316 ( .A(n295), .B(n489), .Z(\ab[14][60] ) );
  AN2P U2317 ( .A(n295), .B(B[59]), .Z(\ab[14][59] ) );
  AN2P U2318 ( .A(n294), .B(B[58]), .Z(\ab[14][58] ) );
  AN2P U2319 ( .A(n294), .B(B[57]), .Z(\ab[14][57] ) );
  AN2P U2320 ( .A(n294), .B(B[56]), .Z(\ab[14][56] ) );
  AN2P U2321 ( .A(n294), .B(n490), .Z(\ab[14][55] ) );
  AN2P U2322 ( .A(n294), .B(B[54]), .Z(\ab[14][54] ) );
  AN2P U2323 ( .A(n294), .B(B[53]), .Z(\ab[14][53] ) );
  AN2P U2324 ( .A(n294), .B(B[52]), .Z(\ab[14][52] ) );
  AN2P U2325 ( .A(n294), .B(B[51]), .Z(\ab[14][51] ) );
  AN2P U2326 ( .A(n294), .B(B[50]), .Z(\ab[14][50] ) );
  AN2P U2327 ( .A(n294), .B(B[49]), .Z(\ab[14][49] ) );
  AN2P U2328 ( .A(n294), .B(B[48]), .Z(\ab[14][48] ) );
  AN2P U2329 ( .A(n294), .B(B[47]), .Z(\ab[14][47] ) );
  AN2P U2330 ( .A(n293), .B(B[46]), .Z(\ab[14][46] ) );
  AN2P U2331 ( .A(n293), .B(B[45]), .Z(\ab[14][45] ) );
  AN2P U2332 ( .A(n293), .B(B[44]), .Z(\ab[14][44] ) );
  AN2P U2333 ( .A(n293), .B(B[43]), .Z(\ab[14][43] ) );
  AN2P U2334 ( .A(n293), .B(B[42]), .Z(\ab[14][42] ) );
  AN2P U2335 ( .A(n293), .B(B[41]), .Z(\ab[14][41] ) );
  AN2P U2336 ( .A(n293), .B(B[40]), .Z(\ab[14][40] ) );
  AN2P U2337 ( .A(n293), .B(B[39]), .Z(\ab[14][39] ) );
  AN2P U2338 ( .A(n293), .B(n452), .Z(\ab[14][38] ) );
  AN2P U2339 ( .A(n293), .B(n448), .Z(\ab[14][37] ) );
  AN2P U2340 ( .A(n293), .B(n444), .Z(\ab[14][36] ) );
  AN2P U2341 ( .A(n293), .B(n440), .Z(\ab[14][35] ) );
  AN2P U2342 ( .A(n292), .B(n436), .Z(\ab[14][34] ) );
  AN2P U2343 ( .A(n292), .B(n432), .Z(\ab[14][33] ) );
  AN2P U2344 ( .A(n292), .B(n428), .Z(\ab[14][32] ) );
  AN2P U2345 ( .A(n292), .B(n424), .Z(\ab[14][31] ) );
  AN2P U2346 ( .A(n292), .B(n420), .Z(\ab[14][30] ) );
  AN2P U2347 ( .A(n292), .B(n416), .Z(\ab[14][29] ) );
  AN2P U2348 ( .A(n292), .B(n412), .Z(\ab[14][28] ) );
  AN2P U2349 ( .A(n292), .B(n408), .Z(\ab[14][27] ) );
  AN2P U2350 ( .A(n292), .B(n404), .Z(\ab[14][26] ) );
  AN2P U2351 ( .A(n292), .B(n400), .Z(\ab[14][25] ) );
  AN2P U2352 ( .A(n292), .B(n396), .Z(\ab[14][24] ) );
  AN2P U2353 ( .A(n292), .B(n392), .Z(\ab[14][23] ) );
  AN2P U2354 ( .A(n291), .B(n388), .Z(\ab[14][22] ) );
  AN2P U2355 ( .A(n291), .B(n384), .Z(\ab[14][21] ) );
  AN2P U2356 ( .A(n291), .B(n380), .Z(\ab[14][20] ) );
  AN2P U2357 ( .A(n291), .B(n376), .Z(\ab[14][19] ) );
  AN2P U2358 ( .A(n291), .B(n372), .Z(\ab[14][18] ) );
  AN2P U2359 ( .A(n291), .B(n368), .Z(\ab[14][17] ) );
  AN2P U2360 ( .A(n291), .B(n364), .Z(\ab[14][16] ) );
  AN2P U2361 ( .A(n291), .B(n360), .Z(\ab[14][15] ) );
  AN2P U2362 ( .A(n291), .B(n356), .Z(\ab[14][14] ) );
  AN2P U2363 ( .A(n291), .B(n352), .Z(\ab[14][13] ) );
  AN2P U2364 ( .A(n291), .B(n348), .Z(\ab[14][12] ) );
  AN2P U2365 ( .A(n291), .B(n344), .Z(\ab[14][11] ) );
  AN2P U2366 ( .A(n290), .B(n340), .Z(\ab[14][10] ) );
  AN2P U2367 ( .A(n290), .B(n336), .Z(\ab[14][9] ) );
  AN2P U2368 ( .A(n290), .B(n332), .Z(\ab[14][8] ) );
  AN2P U2369 ( .A(n290), .B(n328), .Z(\ab[14][7] ) );
  AN2P U2370 ( .A(n290), .B(n324), .Z(\ab[14][6] ) );
  AN2P U2371 ( .A(n290), .B(n320), .Z(\ab[14][5] ) );
  AN2P U2372 ( .A(n290), .B(n316), .Z(\ab[14][4] ) );
  AN2P U2373 ( .A(n290), .B(n312), .Z(\ab[14][3] ) );
  AN2P U2374 ( .A(n290), .B(n308), .Z(\ab[14][2] ) );
  AN2P U2375 ( .A(n290), .B(n304), .Z(\ab[14][1] ) );
  AN2P U2376 ( .A(n290), .B(n300), .Z(\ab[14][0] ) );
  AN2P U2377 ( .A(n290), .B(n491), .Z(\ab[14][95] ) );
  AN2P U2378 ( .A(n452), .B(n11), .Z(\ab[15][38] ) );
  AN2P U2379 ( .A(n448), .B(n11), .Z(\ab[15][37] ) );
  AN2P U2380 ( .A(n444), .B(n11), .Z(\ab[15][36] ) );
  AN2P U2381 ( .A(n440), .B(n11), .Z(\ab[15][35] ) );
  AN2P U2382 ( .A(n436), .B(n11), .Z(\ab[15][34] ) );
  AN2P U2383 ( .A(n432), .B(n11), .Z(\ab[15][33] ) );
  AN2P U2384 ( .A(n428), .B(n11), .Z(\ab[15][32] ) );
  AN2P U2385 ( .A(n424), .B(n11), .Z(\ab[15][31] ) );
  AN2P U2386 ( .A(n420), .B(n12), .Z(\ab[15][30] ) );
  AN2P U2387 ( .A(n416), .B(n12), .Z(\ab[15][29] ) );
  AN2P U2388 ( .A(n412), .B(n12), .Z(\ab[15][28] ) );
  AN2P U2389 ( .A(n408), .B(n12), .Z(\ab[15][27] ) );
  AN2P U2390 ( .A(n404), .B(n12), .Z(\ab[15][26] ) );
  AN2P U2391 ( .A(n400), .B(n12), .Z(\ab[15][25] ) );
  AN2P U2392 ( .A(n396), .B(n12), .Z(\ab[15][24] ) );
  AN2P U2393 ( .A(n392), .B(n12), .Z(\ab[15][23] ) );
  AN2P U2394 ( .A(n388), .B(n13), .Z(\ab[15][22] ) );
  AN2P U2395 ( .A(n384), .B(n13), .Z(\ab[15][21] ) );
  AN2P U2396 ( .A(n380), .B(n13), .Z(\ab[15][20] ) );
  AN2P U2397 ( .A(n376), .B(n13), .Z(\ab[15][19] ) );
  AN2P U2398 ( .A(n372), .B(n13), .Z(\ab[15][18] ) );
  AN2P U2399 ( .A(n368), .B(n13), .Z(\ab[15][17] ) );
  AN2P U2400 ( .A(n364), .B(n13), .Z(\ab[15][16] ) );
  AN2P U2401 ( .A(n360), .B(n13), .Z(\ab[15][15] ) );
  AN2P U2402 ( .A(n356), .B(n14), .Z(\ab[15][14] ) );
  AN2P U2403 ( .A(n352), .B(n14), .Z(\ab[15][13] ) );
  AN2P U2404 ( .A(n348), .B(n14), .Z(\ab[15][12] ) );
  AN2P U2405 ( .A(n344), .B(n14), .Z(\ab[15][11] ) );
  AN2P U2406 ( .A(n340), .B(n14), .Z(\ab[15][10] ) );
  AN2P U2407 ( .A(n336), .B(n14), .Z(\ab[15][9] ) );
  AN2P U2408 ( .A(n332), .B(n14), .Z(\ab[15][8] ) );
  AN2P U2409 ( .A(n328), .B(n14), .Z(\ab[15][7] ) );
  AN2P U2410 ( .A(n324), .B(n15), .Z(\ab[15][6] ) );
  AN2P U2411 ( .A(n320), .B(n15), .Z(\ab[15][5] ) );
  AN2P U2412 ( .A(n316), .B(n15), .Z(\ab[15][4] ) );
  AN2P U2413 ( .A(n312), .B(n15), .Z(\ab[15][3] ) );
  AN2P U2414 ( .A(n308), .B(n15), .Z(\ab[15][2] ) );
  AN2P U2415 ( .A(n304), .B(n15), .Z(\ab[15][1] ) );
  AN2P U2416 ( .A(n300), .B(n15), .Z(\ab[15][0] ) );
  AN2P U2417 ( .A(n452), .B(n159), .Z(\ab[16][38] ) );
  AN2P U2418 ( .A(n448), .B(n159), .Z(\ab[16][37] ) );
  AN2P U2419 ( .A(n444), .B(n159), .Z(\ab[16][36] ) );
  AN2P U2420 ( .A(n440), .B(n159), .Z(\ab[16][35] ) );
  AN2P U2421 ( .A(n436), .B(n159), .Z(\ab[16][34] ) );
  AN2P U2422 ( .A(n432), .B(n159), .Z(\ab[16][33] ) );
  AN2P U2423 ( .A(n428), .B(n159), .Z(\ab[16][32] ) );
  AN2P U2424 ( .A(n424), .B(n159), .Z(\ab[16][31] ) );
  AN2P U2425 ( .A(n420), .B(n160), .Z(\ab[16][30] ) );
  AN2P U2426 ( .A(n416), .B(n160), .Z(\ab[16][29] ) );
  AN2P U2427 ( .A(n412), .B(n160), .Z(\ab[16][28] ) );
  AN2P U2428 ( .A(n408), .B(n160), .Z(\ab[16][27] ) );
  AN2P U2429 ( .A(n404), .B(n160), .Z(\ab[16][26] ) );
  AN2P U2430 ( .A(n400), .B(n160), .Z(\ab[16][25] ) );
  AN2P U2431 ( .A(n396), .B(n160), .Z(\ab[16][24] ) );
  AN2P U2432 ( .A(n392), .B(n160), .Z(\ab[16][23] ) );
  AN2P U2433 ( .A(n388), .B(n161), .Z(\ab[16][22] ) );
  AN2P U2434 ( .A(n384), .B(n161), .Z(\ab[16][21] ) );
  AN2P U2435 ( .A(n380), .B(n161), .Z(\ab[16][20] ) );
  AN2P U2436 ( .A(n376), .B(n161), .Z(\ab[16][19] ) );
  AN2P U2437 ( .A(n372), .B(n161), .Z(\ab[16][18] ) );
  AN2P U2438 ( .A(n368), .B(n161), .Z(\ab[16][17] ) );
  AN2P U2439 ( .A(n364), .B(n161), .Z(\ab[16][16] ) );
  AN2P U2440 ( .A(n360), .B(n161), .Z(\ab[16][15] ) );
  AN2P U2441 ( .A(n356), .B(n162), .Z(\ab[16][14] ) );
  AN2P U2442 ( .A(n352), .B(n162), .Z(\ab[16][13] ) );
  AN2P U2443 ( .A(n348), .B(n162), .Z(\ab[16][12] ) );
  AN2P U2444 ( .A(n344), .B(n162), .Z(\ab[16][11] ) );
  AN2P U2445 ( .A(n340), .B(n162), .Z(\ab[16][10] ) );
  AN2P U2446 ( .A(n336), .B(n162), .Z(\ab[16][9] ) );
  AN2P U2447 ( .A(n332), .B(n162), .Z(\ab[16][8] ) );
  AN2P U2448 ( .A(n328), .B(n162), .Z(\ab[16][7] ) );
  AN2P U2449 ( .A(n324), .B(n163), .Z(\ab[16][6] ) );
  AN2P U2450 ( .A(n320), .B(n163), .Z(\ab[16][5] ) );
  AN2P U2451 ( .A(n316), .B(n163), .Z(\ab[16][4] ) );
  AN2P U2452 ( .A(n312), .B(n163), .Z(\ab[16][3] ) );
  AN2P U2453 ( .A(n308), .B(n163), .Z(\ab[16][2] ) );
  AN2P U2454 ( .A(n304), .B(n163), .Z(\ab[16][1] ) );
  AN2P U2455 ( .A(n300), .B(n163), .Z(\ab[16][0] ) );
  AN2P U2456 ( .A(n452), .B(n148), .Z(\ab[17][38] ) );
  AN2P U2457 ( .A(n448), .B(n148), .Z(\ab[17][37] ) );
  AN2P U2458 ( .A(n444), .B(n148), .Z(\ab[17][36] ) );
  AN2P U2459 ( .A(n440), .B(n148), .Z(\ab[17][35] ) );
  AN2P U2460 ( .A(n436), .B(n148), .Z(\ab[17][34] ) );
  AN2P U2461 ( .A(n432), .B(n148), .Z(\ab[17][33] ) );
  AN2P U2462 ( .A(n428), .B(n148), .Z(\ab[17][32] ) );
  AN2P U2463 ( .A(n424), .B(n148), .Z(\ab[17][31] ) );
  AN2P U2464 ( .A(n420), .B(n149), .Z(\ab[17][30] ) );
  AN2P U2465 ( .A(n416), .B(n149), .Z(\ab[17][29] ) );
  AN2P U2466 ( .A(n412), .B(n149), .Z(\ab[17][28] ) );
  AN2P U2467 ( .A(n408), .B(n149), .Z(\ab[17][27] ) );
  AN2P U2468 ( .A(n404), .B(n149), .Z(\ab[17][26] ) );
  AN2P U2469 ( .A(n400), .B(n149), .Z(\ab[17][25] ) );
  AN2P U2470 ( .A(n396), .B(n149), .Z(\ab[17][24] ) );
  AN2P U2471 ( .A(n392), .B(n149), .Z(\ab[17][23] ) );
  AN2P U2472 ( .A(n388), .B(n150), .Z(\ab[17][22] ) );
  AN2P U2473 ( .A(n384), .B(n150), .Z(\ab[17][21] ) );
  AN2P U2474 ( .A(n380), .B(n150), .Z(\ab[17][20] ) );
  AN2P U2475 ( .A(n376), .B(n150), .Z(\ab[17][19] ) );
  AN2P U2476 ( .A(n372), .B(n150), .Z(\ab[17][18] ) );
  AN2P U2477 ( .A(n368), .B(n150), .Z(\ab[17][17] ) );
  AN2P U2478 ( .A(n364), .B(n150), .Z(\ab[17][16] ) );
  AN2P U2479 ( .A(n360), .B(n150), .Z(\ab[17][15] ) );
  AN2P U2480 ( .A(n356), .B(n151), .Z(\ab[17][14] ) );
  AN2P U2481 ( .A(n352), .B(n151), .Z(\ab[17][13] ) );
  AN2P U2482 ( .A(n348), .B(n151), .Z(\ab[17][12] ) );
  AN2P U2483 ( .A(n344), .B(n151), .Z(\ab[17][11] ) );
  AN2P U2484 ( .A(n340), .B(n151), .Z(\ab[17][10] ) );
  AN2P U2485 ( .A(n336), .B(n151), .Z(\ab[17][9] ) );
  AN2P U2486 ( .A(n332), .B(n151), .Z(\ab[17][8] ) );
  AN2P U2487 ( .A(n328), .B(n151), .Z(\ab[17][7] ) );
  AN2P U2488 ( .A(n324), .B(n152), .Z(\ab[17][6] ) );
  AN2P U2489 ( .A(n320), .B(n152), .Z(\ab[17][5] ) );
  AN2P U2490 ( .A(n316), .B(n152), .Z(\ab[17][4] ) );
  AN2P U2491 ( .A(n312), .B(n152), .Z(\ab[17][3] ) );
  AN2P U2492 ( .A(n308), .B(n152), .Z(\ab[17][2] ) );
  AN2P U2493 ( .A(n304), .B(n152), .Z(\ab[17][1] ) );
  AN2P U2494 ( .A(n300), .B(n152), .Z(\ab[17][0] ) );
  AN2P U2495 ( .A(n451), .B(n137), .Z(\ab[18][38] ) );
  AN2P U2496 ( .A(n447), .B(n137), .Z(\ab[18][37] ) );
  AN2P U2497 ( .A(n443), .B(n137), .Z(\ab[18][36] ) );
  AN2P U2498 ( .A(n439), .B(n137), .Z(\ab[18][35] ) );
  AN2P U2499 ( .A(n435), .B(n137), .Z(\ab[18][34] ) );
  AN2P U2500 ( .A(n431), .B(n137), .Z(\ab[18][33] ) );
  AN2P U2501 ( .A(n427), .B(n137), .Z(\ab[18][32] ) );
  AN2P U2502 ( .A(n423), .B(n137), .Z(\ab[18][31] ) );
  AN2P U2503 ( .A(n419), .B(n138), .Z(\ab[18][30] ) );
  AN2P U2504 ( .A(n415), .B(n138), .Z(\ab[18][29] ) );
  AN2P U2505 ( .A(n411), .B(n138), .Z(\ab[18][28] ) );
  AN2P U2506 ( .A(n407), .B(n138), .Z(\ab[18][27] ) );
  AN2P U2507 ( .A(n403), .B(n138), .Z(\ab[18][26] ) );
  AN2P U2508 ( .A(n399), .B(n138), .Z(\ab[18][25] ) );
  AN2P U2509 ( .A(n395), .B(n138), .Z(\ab[18][24] ) );
  AN2P U2510 ( .A(n391), .B(n138), .Z(\ab[18][23] ) );
  AN2P U2511 ( .A(n387), .B(n139), .Z(\ab[18][22] ) );
  AN2P U2512 ( .A(n383), .B(n139), .Z(\ab[18][21] ) );
  AN2P U2513 ( .A(n379), .B(n139), .Z(\ab[18][20] ) );
  AN2P U2514 ( .A(n375), .B(n139), .Z(\ab[18][19] ) );
  AN2P U2515 ( .A(n371), .B(n139), .Z(\ab[18][18] ) );
  AN2P U2516 ( .A(n367), .B(n139), .Z(\ab[18][17] ) );
  AN2P U2517 ( .A(n363), .B(n139), .Z(\ab[18][16] ) );
  AN2P U2518 ( .A(n359), .B(n139), .Z(\ab[18][15] ) );
  AN2P U2519 ( .A(n355), .B(n140), .Z(\ab[18][14] ) );
  AN2P U2520 ( .A(n351), .B(n140), .Z(\ab[18][13] ) );
  AN2P U2521 ( .A(n347), .B(n140), .Z(\ab[18][12] ) );
  AN2P U2522 ( .A(n343), .B(n140), .Z(\ab[18][11] ) );
  AN2P U2523 ( .A(n339), .B(n140), .Z(\ab[18][10] ) );
  AN2P U2524 ( .A(n335), .B(n140), .Z(\ab[18][9] ) );
  AN2P U2525 ( .A(n331), .B(n140), .Z(\ab[18][8] ) );
  AN2P U2526 ( .A(n327), .B(n140), .Z(\ab[18][7] ) );
  AN2P U2527 ( .A(n323), .B(n141), .Z(\ab[18][6] ) );
  AN2P U2528 ( .A(n319), .B(n141), .Z(\ab[18][5] ) );
  AN2P U2529 ( .A(n315), .B(n141), .Z(\ab[18][4] ) );
  AN2P U2530 ( .A(n311), .B(n141), .Z(\ab[18][3] ) );
  AN2P U2531 ( .A(n307), .B(n141), .Z(\ab[18][2] ) );
  AN2P U2532 ( .A(n303), .B(n141), .Z(\ab[18][1] ) );
  AN2P U2533 ( .A(n299), .B(n141), .Z(\ab[18][0] ) );
  AN2P U2534 ( .A(n451), .B(n126), .Z(\ab[19][38] ) );
  AN2P U2535 ( .A(n447), .B(n126), .Z(\ab[19][37] ) );
  AN2P U2536 ( .A(n443), .B(n126), .Z(\ab[19][36] ) );
  AN2P U2537 ( .A(n439), .B(n126), .Z(\ab[19][35] ) );
  AN2P U2538 ( .A(n435), .B(n126), .Z(\ab[19][34] ) );
  AN2P U2539 ( .A(n431), .B(n126), .Z(\ab[19][33] ) );
  AN2P U2540 ( .A(n427), .B(n126), .Z(\ab[19][32] ) );
  AN2P U2541 ( .A(n423), .B(n126), .Z(\ab[19][31] ) );
  AN2P U2542 ( .A(n419), .B(n127), .Z(\ab[19][30] ) );
  AN2P U2543 ( .A(n415), .B(n127), .Z(\ab[19][29] ) );
  AN2P U2544 ( .A(n411), .B(n127), .Z(\ab[19][28] ) );
  AN2P U2545 ( .A(n407), .B(n127), .Z(\ab[19][27] ) );
  AN2P U2546 ( .A(n403), .B(n127), .Z(\ab[19][26] ) );
  AN2P U2547 ( .A(n399), .B(n127), .Z(\ab[19][25] ) );
  AN2P U2548 ( .A(n395), .B(n127), .Z(\ab[19][24] ) );
  AN2P U2549 ( .A(n391), .B(n127), .Z(\ab[19][23] ) );
  AN2P U2550 ( .A(n387), .B(n128), .Z(\ab[19][22] ) );
  AN2P U2551 ( .A(n383), .B(n128), .Z(\ab[19][21] ) );
  AN2P U2552 ( .A(n379), .B(n128), .Z(\ab[19][20] ) );
  AN2P U2553 ( .A(n375), .B(n128), .Z(\ab[19][19] ) );
  AN2P U2554 ( .A(n371), .B(n128), .Z(\ab[19][18] ) );
  AN2P U2555 ( .A(n367), .B(n128), .Z(\ab[19][17] ) );
  AN2P U2556 ( .A(n363), .B(n128), .Z(\ab[19][16] ) );
  AN2P U2557 ( .A(n359), .B(n128), .Z(\ab[19][15] ) );
  AN2P U2558 ( .A(n355), .B(n129), .Z(\ab[19][14] ) );
  AN2P U2559 ( .A(n351), .B(n129), .Z(\ab[19][13] ) );
  AN2P U2560 ( .A(n347), .B(n129), .Z(\ab[19][12] ) );
  AN2P U2561 ( .A(n343), .B(n129), .Z(\ab[19][11] ) );
  AN2P U2562 ( .A(n339), .B(n129), .Z(\ab[19][10] ) );
  AN2P U2563 ( .A(n335), .B(n129), .Z(\ab[19][9] ) );
  AN2P U2564 ( .A(n331), .B(n129), .Z(\ab[19][8] ) );
  AN2P U2565 ( .A(n327), .B(n129), .Z(\ab[19][7] ) );
  AN2P U2566 ( .A(n323), .B(n130), .Z(\ab[19][6] ) );
  AN2P U2567 ( .A(n319), .B(n130), .Z(\ab[19][5] ) );
  AN2P U2568 ( .A(n315), .B(n130), .Z(\ab[19][4] ) );
  AN2P U2569 ( .A(n311), .B(n130), .Z(\ab[19][3] ) );
  AN2P U2570 ( .A(n307), .B(n130), .Z(\ab[19][2] ) );
  AN2P U2571 ( .A(n303), .B(n130), .Z(\ab[19][1] ) );
  AN2P U2572 ( .A(n299), .B(n130), .Z(\ab[19][0] ) );
  AN2P U2573 ( .A(n451), .B(n115), .Z(\ab[20][38] ) );
  AN2P U2574 ( .A(n447), .B(n115), .Z(\ab[20][37] ) );
  AN2P U2575 ( .A(n443), .B(n115), .Z(\ab[20][36] ) );
  AN2P U2576 ( .A(n439), .B(n115), .Z(\ab[20][35] ) );
  AN2P U2577 ( .A(n435), .B(n115), .Z(\ab[20][34] ) );
  AN2P U2578 ( .A(n431), .B(n115), .Z(\ab[20][33] ) );
  AN2P U2579 ( .A(n427), .B(n115), .Z(\ab[20][32] ) );
  AN2P U2580 ( .A(n423), .B(n115), .Z(\ab[20][31] ) );
  AN2P U2581 ( .A(n419), .B(n116), .Z(\ab[20][30] ) );
  AN2P U2582 ( .A(n415), .B(n116), .Z(\ab[20][29] ) );
  AN2P U2583 ( .A(n411), .B(n116), .Z(\ab[20][28] ) );
  AN2P U2584 ( .A(n407), .B(n116), .Z(\ab[20][27] ) );
  AN2P U2585 ( .A(n403), .B(n116), .Z(\ab[20][26] ) );
  AN2P U2586 ( .A(n399), .B(n116), .Z(\ab[20][25] ) );
  AN2P U2587 ( .A(n395), .B(n116), .Z(\ab[20][24] ) );
  AN2P U2588 ( .A(n391), .B(n116), .Z(\ab[20][23] ) );
  AN2P U2589 ( .A(n387), .B(n117), .Z(\ab[20][22] ) );
  AN2P U2590 ( .A(n383), .B(n117), .Z(\ab[20][21] ) );
  AN2P U2591 ( .A(n379), .B(n117), .Z(\ab[20][20] ) );
  AN2P U2592 ( .A(n375), .B(n117), .Z(\ab[20][19] ) );
  AN2P U2593 ( .A(n371), .B(n117), .Z(\ab[20][18] ) );
  AN2P U2594 ( .A(n367), .B(n117), .Z(\ab[20][17] ) );
  AN2P U2595 ( .A(n363), .B(n117), .Z(\ab[20][16] ) );
  AN2P U2596 ( .A(n359), .B(n117), .Z(\ab[20][15] ) );
  AN2P U2597 ( .A(n355), .B(n118), .Z(\ab[20][14] ) );
  AN2P U2598 ( .A(n351), .B(n118), .Z(\ab[20][13] ) );
  AN2P U2599 ( .A(n347), .B(n118), .Z(\ab[20][12] ) );
  AN2P U2600 ( .A(n343), .B(n118), .Z(\ab[20][11] ) );
  AN2P U2601 ( .A(n339), .B(n118), .Z(\ab[20][10] ) );
  AN2P U2602 ( .A(n335), .B(n118), .Z(\ab[20][9] ) );
  AN2P U2603 ( .A(n331), .B(n118), .Z(\ab[20][8] ) );
  AN2P U2604 ( .A(n327), .B(n118), .Z(\ab[20][7] ) );
  AN2P U2605 ( .A(n323), .B(n119), .Z(\ab[20][6] ) );
  AN2P U2606 ( .A(n319), .B(n119), .Z(\ab[20][5] ) );
  AN2P U2607 ( .A(n315), .B(n119), .Z(\ab[20][4] ) );
  AN2P U2608 ( .A(n311), .B(n119), .Z(\ab[20][3] ) );
  AN2P U2609 ( .A(n307), .B(n119), .Z(\ab[20][2] ) );
  AN2P U2610 ( .A(n303), .B(n119), .Z(\ab[20][1] ) );
  AN2P U2611 ( .A(n299), .B(n119), .Z(\ab[20][0] ) );
  AN2P U2612 ( .A(n451), .B(n104), .Z(\ab[21][38] ) );
  AN2P U2613 ( .A(n447), .B(n104), .Z(\ab[21][37] ) );
  AN2P U2614 ( .A(n443), .B(n104), .Z(\ab[21][36] ) );
  AN2P U2615 ( .A(n439), .B(n104), .Z(\ab[21][35] ) );
  AN2P U2616 ( .A(n435), .B(n104), .Z(\ab[21][34] ) );
  AN2P U2617 ( .A(n431), .B(n104), .Z(\ab[21][33] ) );
  AN2P U2618 ( .A(n427), .B(n104), .Z(\ab[21][32] ) );
  AN2P U2619 ( .A(n423), .B(n104), .Z(\ab[21][31] ) );
  AN2P U2620 ( .A(n419), .B(n105), .Z(\ab[21][30] ) );
  AN2P U2621 ( .A(n415), .B(n105), .Z(\ab[21][29] ) );
  AN2P U2622 ( .A(n411), .B(n105), .Z(\ab[21][28] ) );
  AN2P U2623 ( .A(n407), .B(n105), .Z(\ab[21][27] ) );
  AN2P U2624 ( .A(n403), .B(n105), .Z(\ab[21][26] ) );
  AN2P U2625 ( .A(n399), .B(n105), .Z(\ab[21][25] ) );
  AN2P U2626 ( .A(n395), .B(n105), .Z(\ab[21][24] ) );
  AN2P U2627 ( .A(n391), .B(n105), .Z(\ab[21][23] ) );
  AN2P U2628 ( .A(n387), .B(n106), .Z(\ab[21][22] ) );
  AN2P U2629 ( .A(n383), .B(n106), .Z(\ab[21][21] ) );
  AN2P U2630 ( .A(n379), .B(n106), .Z(\ab[21][20] ) );
  AN2P U2631 ( .A(n375), .B(n106), .Z(\ab[21][19] ) );
  AN2P U2632 ( .A(n371), .B(n106), .Z(\ab[21][18] ) );
  AN2P U2633 ( .A(n367), .B(n106), .Z(\ab[21][17] ) );
  AN2P U2634 ( .A(n363), .B(n106), .Z(\ab[21][16] ) );
  AN2P U2635 ( .A(n359), .B(n106), .Z(\ab[21][15] ) );
  AN2P U2636 ( .A(n355), .B(n107), .Z(\ab[21][14] ) );
  AN2P U2637 ( .A(n351), .B(n107), .Z(\ab[21][13] ) );
  AN2P U2638 ( .A(n347), .B(n107), .Z(\ab[21][12] ) );
  AN2P U2639 ( .A(n343), .B(n107), .Z(\ab[21][11] ) );
  AN2P U2640 ( .A(n339), .B(n107), .Z(\ab[21][10] ) );
  AN2P U2641 ( .A(n335), .B(n107), .Z(\ab[21][9] ) );
  AN2P U2642 ( .A(n331), .B(n107), .Z(\ab[21][8] ) );
  AN2P U2643 ( .A(n327), .B(n107), .Z(\ab[21][7] ) );
  AN2P U2644 ( .A(n323), .B(n108), .Z(\ab[21][6] ) );
  AN2P U2645 ( .A(n319), .B(n108), .Z(\ab[21][5] ) );
  AN2P U2646 ( .A(n315), .B(n108), .Z(\ab[21][4] ) );
  AN2P U2647 ( .A(n311), .B(n108), .Z(\ab[21][3] ) );
  AN2P U2648 ( .A(n307), .B(n108), .Z(\ab[21][2] ) );
  AN2P U2649 ( .A(n303), .B(n108), .Z(\ab[21][1] ) );
  AN2P U2650 ( .A(n299), .B(n108), .Z(\ab[21][0] ) );
  AN2P U2651 ( .A(n451), .B(n93), .Z(\ab[22][38] ) );
  AN2P U2652 ( .A(n447), .B(n93), .Z(\ab[22][37] ) );
  AN2P U2653 ( .A(n443), .B(n93), .Z(\ab[22][36] ) );
  AN2P U2654 ( .A(n439), .B(n93), .Z(\ab[22][35] ) );
  AN2P U2655 ( .A(n435), .B(n93), .Z(\ab[22][34] ) );
  AN2P U2656 ( .A(n431), .B(n93), .Z(\ab[22][33] ) );
  AN2P U2657 ( .A(n427), .B(n93), .Z(\ab[22][32] ) );
  AN2P U2658 ( .A(n423), .B(n93), .Z(\ab[22][31] ) );
  AN2P U2659 ( .A(n419), .B(n94), .Z(\ab[22][30] ) );
  AN2P U2660 ( .A(n415), .B(n94), .Z(\ab[22][29] ) );
  AN2P U2661 ( .A(n411), .B(n94), .Z(\ab[22][28] ) );
  AN2P U2662 ( .A(n407), .B(n94), .Z(\ab[22][27] ) );
  AN2P U2663 ( .A(n403), .B(n94), .Z(\ab[22][26] ) );
  AN2P U2664 ( .A(n399), .B(n94), .Z(\ab[22][25] ) );
  AN2P U2665 ( .A(n395), .B(n94), .Z(\ab[22][24] ) );
  AN2P U2666 ( .A(n391), .B(n94), .Z(\ab[22][23] ) );
  AN2P U2667 ( .A(n387), .B(n95), .Z(\ab[22][22] ) );
  AN2P U2668 ( .A(n383), .B(n95), .Z(\ab[22][21] ) );
  AN2P U2669 ( .A(n379), .B(n95), .Z(\ab[22][20] ) );
  AN2P U2670 ( .A(n375), .B(n95), .Z(\ab[22][19] ) );
  AN2P U2671 ( .A(n371), .B(n95), .Z(\ab[22][18] ) );
  AN2P U2672 ( .A(n367), .B(n95), .Z(\ab[22][17] ) );
  AN2P U2673 ( .A(n363), .B(n95), .Z(\ab[22][16] ) );
  AN2P U2674 ( .A(n359), .B(n95), .Z(\ab[22][15] ) );
  AN2P U2675 ( .A(n355), .B(n96), .Z(\ab[22][14] ) );
  AN2P U2676 ( .A(n351), .B(n96), .Z(\ab[22][13] ) );
  AN2P U2677 ( .A(n347), .B(n96), .Z(\ab[22][12] ) );
  AN2P U2678 ( .A(n343), .B(n96), .Z(\ab[22][11] ) );
  AN2P U2679 ( .A(n339), .B(n96), .Z(\ab[22][10] ) );
  AN2P U2680 ( .A(n335), .B(n96), .Z(\ab[22][9] ) );
  AN2P U2681 ( .A(n331), .B(n96), .Z(\ab[22][8] ) );
  AN2P U2682 ( .A(n327), .B(n96), .Z(\ab[22][7] ) );
  AN2P U2683 ( .A(n323), .B(n97), .Z(\ab[22][6] ) );
  AN2P U2684 ( .A(n319), .B(n97), .Z(\ab[22][5] ) );
  AN2P U2685 ( .A(n315), .B(n97), .Z(\ab[22][4] ) );
  AN2P U2686 ( .A(n311), .B(n97), .Z(\ab[22][3] ) );
  AN2P U2687 ( .A(n307), .B(n97), .Z(\ab[22][2] ) );
  AN2P U2688 ( .A(n303), .B(n97), .Z(\ab[22][1] ) );
  AN2P U2689 ( .A(n299), .B(n97), .Z(\ab[22][0] ) );
  AN2P U2690 ( .A(n451), .B(n88), .Z(\ab[23][38] ) );
  AN2P U2691 ( .A(n447), .B(n88), .Z(\ab[23][37] ) );
  AN2P U2692 ( .A(n443), .B(n88), .Z(\ab[23][36] ) );
  AN2P U2693 ( .A(n439), .B(n88), .Z(\ab[23][35] ) );
  AN2P U2694 ( .A(n435), .B(n88), .Z(\ab[23][34] ) );
  AN2P U2695 ( .A(n431), .B(n88), .Z(\ab[23][33] ) );
  AN2P U2696 ( .A(n427), .B(n88), .Z(\ab[23][32] ) );
  AN2P U2697 ( .A(n423), .B(n88), .Z(\ab[23][31] ) );
  AN2P U2698 ( .A(n419), .B(n89), .Z(\ab[23][30] ) );
  AN2P U2699 ( .A(n415), .B(n89), .Z(\ab[23][29] ) );
  AN2P U2700 ( .A(n411), .B(n89), .Z(\ab[23][28] ) );
  AN2P U2701 ( .A(n407), .B(n89), .Z(\ab[23][27] ) );
  AN2P U2702 ( .A(n403), .B(n89), .Z(\ab[23][26] ) );
  AN2P U2703 ( .A(n399), .B(n89), .Z(\ab[23][25] ) );
  AN2P U2704 ( .A(n395), .B(n89), .Z(\ab[23][24] ) );
  AN2P U2705 ( .A(n391), .B(n89), .Z(\ab[23][23] ) );
  AN2P U2706 ( .A(n387), .B(n90), .Z(\ab[23][22] ) );
  AN2P U2707 ( .A(n383), .B(n90), .Z(\ab[23][21] ) );
  AN2P U2708 ( .A(n379), .B(n90), .Z(\ab[23][20] ) );
  AN2P U2709 ( .A(n375), .B(n90), .Z(\ab[23][19] ) );
  AN2P U2710 ( .A(n371), .B(n90), .Z(\ab[23][18] ) );
  AN2P U2711 ( .A(n367), .B(n90), .Z(\ab[23][17] ) );
  AN2P U2712 ( .A(n363), .B(n90), .Z(\ab[23][16] ) );
  AN2P U2713 ( .A(n359), .B(n90), .Z(\ab[23][15] ) );
  AN2P U2714 ( .A(n355), .B(n91), .Z(\ab[23][14] ) );
  AN2P U2715 ( .A(n351), .B(n91), .Z(\ab[23][13] ) );
  AN2P U2716 ( .A(n347), .B(n91), .Z(\ab[23][12] ) );
  AN2P U2717 ( .A(n343), .B(n91), .Z(\ab[23][11] ) );
  AN2P U2718 ( .A(n339), .B(n91), .Z(\ab[23][10] ) );
  AN2P U2719 ( .A(n335), .B(n91), .Z(\ab[23][9] ) );
  AN2P U2720 ( .A(n331), .B(n91), .Z(\ab[23][8] ) );
  AN2P U2721 ( .A(n327), .B(n91), .Z(\ab[23][7] ) );
  AN2P U2722 ( .A(n323), .B(n92), .Z(\ab[23][6] ) );
  AN2P U2723 ( .A(n319), .B(n92), .Z(\ab[23][5] ) );
  AN2P U2724 ( .A(n315), .B(n92), .Z(\ab[23][4] ) );
  AN2P U2725 ( .A(n311), .B(n92), .Z(\ab[23][3] ) );
  AN2P U2726 ( .A(n307), .B(n92), .Z(\ab[23][2] ) );
  AN2P U2727 ( .A(n303), .B(n92), .Z(\ab[23][1] ) );
  AN2P U2728 ( .A(n299), .B(n92), .Z(\ab[23][0] ) );
  AN2P U2729 ( .A(n451), .B(n77), .Z(\ab[24][38] ) );
  AN2P U2730 ( .A(n447), .B(n77), .Z(\ab[24][37] ) );
  AN2P U2731 ( .A(n443), .B(n77), .Z(\ab[24][36] ) );
  AN2P U2732 ( .A(n439), .B(n77), .Z(\ab[24][35] ) );
  AN2P U2733 ( .A(n435), .B(n77), .Z(\ab[24][34] ) );
  AN2P U2734 ( .A(n431), .B(n77), .Z(\ab[24][33] ) );
  AN2P U2735 ( .A(n427), .B(n77), .Z(\ab[24][32] ) );
  AN2P U2736 ( .A(n423), .B(n77), .Z(\ab[24][31] ) );
  AN2P U2737 ( .A(n419), .B(n78), .Z(\ab[24][30] ) );
  AN2P U2738 ( .A(n415), .B(n78), .Z(\ab[24][29] ) );
  AN2P U2739 ( .A(n411), .B(n78), .Z(\ab[24][28] ) );
  AN2P U2740 ( .A(n407), .B(n78), .Z(\ab[24][27] ) );
  AN2P U2741 ( .A(n403), .B(n78), .Z(\ab[24][26] ) );
  AN2P U2742 ( .A(n399), .B(n78), .Z(\ab[24][25] ) );
  AN2P U2743 ( .A(n395), .B(n78), .Z(\ab[24][24] ) );
  AN2P U2744 ( .A(n391), .B(n78), .Z(\ab[24][23] ) );
  AN2P U2745 ( .A(n387), .B(n79), .Z(\ab[24][22] ) );
  AN2P U2746 ( .A(n383), .B(n79), .Z(\ab[24][21] ) );
  AN2P U2747 ( .A(n379), .B(n79), .Z(\ab[24][20] ) );
  AN2P U2748 ( .A(n375), .B(n79), .Z(\ab[24][19] ) );
  AN2P U2749 ( .A(n371), .B(n79), .Z(\ab[24][18] ) );
  AN2P U2750 ( .A(n367), .B(n79), .Z(\ab[24][17] ) );
  AN2P U2751 ( .A(n363), .B(n79), .Z(\ab[24][16] ) );
  AN2P U2752 ( .A(n359), .B(n79), .Z(\ab[24][15] ) );
  AN2P U2753 ( .A(n355), .B(n80), .Z(\ab[24][14] ) );
  AN2P U2754 ( .A(n351), .B(n80), .Z(\ab[24][13] ) );
  AN2P U2755 ( .A(n347), .B(n80), .Z(\ab[24][12] ) );
  AN2P U2756 ( .A(n343), .B(n80), .Z(\ab[24][11] ) );
  AN2P U2757 ( .A(n339), .B(n80), .Z(\ab[24][10] ) );
  AN2P U2758 ( .A(n335), .B(n80), .Z(\ab[24][9] ) );
  AN2P U2759 ( .A(n331), .B(n80), .Z(\ab[24][8] ) );
  AN2P U2760 ( .A(n327), .B(n80), .Z(\ab[24][7] ) );
  AN2P U2761 ( .A(n323), .B(n81), .Z(\ab[24][6] ) );
  AN2P U2762 ( .A(n319), .B(n81), .Z(\ab[24][5] ) );
  AN2P U2763 ( .A(n315), .B(n81), .Z(\ab[24][4] ) );
  AN2P U2764 ( .A(n311), .B(n81), .Z(\ab[24][3] ) );
  AN2P U2765 ( .A(n307), .B(n81), .Z(\ab[24][2] ) );
  AN2P U2766 ( .A(n303), .B(n81), .Z(\ab[24][1] ) );
  AN2P U2767 ( .A(n299), .B(n81), .Z(\ab[24][0] ) );
  AN2P U2768 ( .A(n451), .B(n66), .Z(\ab[25][38] ) );
  AN2P U2769 ( .A(n447), .B(n66), .Z(\ab[25][37] ) );
  AN2P U2770 ( .A(n443), .B(n66), .Z(\ab[25][36] ) );
  AN2P U2771 ( .A(n439), .B(n66), .Z(\ab[25][35] ) );
  AN2P U2772 ( .A(n435), .B(n66), .Z(\ab[25][34] ) );
  AN2P U2773 ( .A(n431), .B(n66), .Z(\ab[25][33] ) );
  AN2P U2774 ( .A(n427), .B(n66), .Z(\ab[25][32] ) );
  AN2P U2775 ( .A(n423), .B(n66), .Z(\ab[25][31] ) );
  AN2P U2776 ( .A(n419), .B(n67), .Z(\ab[25][30] ) );
  AN2P U2777 ( .A(n415), .B(n67), .Z(\ab[25][29] ) );
  AN2P U2778 ( .A(n411), .B(n67), .Z(\ab[25][28] ) );
  AN2P U2779 ( .A(n407), .B(n67), .Z(\ab[25][27] ) );
  AN2P U2780 ( .A(n403), .B(n67), .Z(\ab[25][26] ) );
  AN2P U2781 ( .A(n399), .B(n67), .Z(\ab[25][25] ) );
  AN2P U2782 ( .A(n395), .B(n67), .Z(\ab[25][24] ) );
  AN2P U2783 ( .A(n391), .B(n67), .Z(\ab[25][23] ) );
  AN2P U2784 ( .A(n387), .B(n68), .Z(\ab[25][22] ) );
  AN2P U2785 ( .A(n383), .B(n68), .Z(\ab[25][21] ) );
  AN2P U2786 ( .A(n379), .B(n68), .Z(\ab[25][20] ) );
  AN2P U2787 ( .A(n375), .B(n68), .Z(\ab[25][19] ) );
  AN2P U2788 ( .A(n371), .B(n68), .Z(\ab[25][18] ) );
  AN2P U2789 ( .A(n367), .B(n68), .Z(\ab[25][17] ) );
  AN2P U2790 ( .A(n363), .B(n68), .Z(\ab[25][16] ) );
  AN2P U2791 ( .A(n359), .B(n68), .Z(\ab[25][15] ) );
  AN2P U2792 ( .A(n355), .B(n69), .Z(\ab[25][14] ) );
  AN2P U2793 ( .A(n351), .B(n69), .Z(\ab[25][13] ) );
  AN2P U2794 ( .A(n347), .B(n69), .Z(\ab[25][12] ) );
  AN2P U2795 ( .A(n343), .B(n69), .Z(\ab[25][11] ) );
  AN2P U2796 ( .A(n339), .B(n69), .Z(\ab[25][10] ) );
  AN2P U2797 ( .A(n335), .B(n69), .Z(\ab[25][9] ) );
  AN2P U2798 ( .A(n331), .B(n69), .Z(\ab[25][8] ) );
  AN2P U2799 ( .A(n327), .B(n69), .Z(\ab[25][7] ) );
  AN2P U2800 ( .A(n323), .B(n70), .Z(\ab[25][6] ) );
  AN2P U2801 ( .A(n319), .B(n70), .Z(\ab[25][5] ) );
  AN2P U2802 ( .A(n315), .B(n70), .Z(\ab[25][4] ) );
  AN2P U2803 ( .A(n311), .B(n70), .Z(\ab[25][3] ) );
  AN2P U2804 ( .A(n307), .B(n70), .Z(\ab[25][2] ) );
  AN2P U2805 ( .A(n303), .B(n70), .Z(\ab[25][1] ) );
  AN2P U2806 ( .A(n299), .B(n70), .Z(\ab[25][0] ) );
  AN2P U2807 ( .A(n451), .B(n55), .Z(\ab[26][38] ) );
  AN2P U2808 ( .A(n447), .B(n55), .Z(\ab[26][37] ) );
  AN2P U2809 ( .A(n443), .B(n55), .Z(\ab[26][36] ) );
  AN2P U2810 ( .A(n439), .B(n55), .Z(\ab[26][35] ) );
  AN2P U2811 ( .A(n435), .B(n55), .Z(\ab[26][34] ) );
  AN2P U2812 ( .A(n431), .B(n55), .Z(\ab[26][33] ) );
  AN2P U2813 ( .A(n427), .B(n55), .Z(\ab[26][32] ) );
  AN2P U2814 ( .A(n423), .B(n55), .Z(\ab[26][31] ) );
  AN2P U2815 ( .A(n419), .B(n56), .Z(\ab[26][30] ) );
  AN2P U2816 ( .A(n415), .B(n56), .Z(\ab[26][29] ) );
  AN2P U2817 ( .A(n411), .B(n56), .Z(\ab[26][28] ) );
  AN2P U2818 ( .A(n407), .B(n56), .Z(\ab[26][27] ) );
  AN2P U2819 ( .A(n403), .B(n56), .Z(\ab[26][26] ) );
  AN2P U2820 ( .A(n399), .B(n56), .Z(\ab[26][25] ) );
  AN2P U2821 ( .A(n395), .B(n56), .Z(\ab[26][24] ) );
  AN2P U2822 ( .A(n391), .B(n56), .Z(\ab[26][23] ) );
  AN2P U2823 ( .A(n387), .B(n57), .Z(\ab[26][22] ) );
  AN2P U2824 ( .A(n383), .B(n57), .Z(\ab[26][21] ) );
  AN2P U2825 ( .A(n379), .B(n57), .Z(\ab[26][20] ) );
  AN2P U2826 ( .A(n375), .B(n57), .Z(\ab[26][19] ) );
  AN2P U2827 ( .A(n371), .B(n57), .Z(\ab[26][18] ) );
  AN2P U2828 ( .A(n367), .B(n57), .Z(\ab[26][17] ) );
  AN2P U2829 ( .A(n363), .B(n57), .Z(\ab[26][16] ) );
  AN2P U2830 ( .A(n359), .B(n57), .Z(\ab[26][15] ) );
  AN2P U2831 ( .A(n355), .B(n58), .Z(\ab[26][14] ) );
  AN2P U2832 ( .A(n351), .B(n58), .Z(\ab[26][13] ) );
  AN2P U2833 ( .A(n347), .B(n58), .Z(\ab[26][12] ) );
  AN2P U2834 ( .A(n343), .B(n58), .Z(\ab[26][11] ) );
  AN2P U2835 ( .A(n339), .B(n58), .Z(\ab[26][10] ) );
  AN2P U2836 ( .A(n335), .B(n58), .Z(\ab[26][9] ) );
  AN2P U2837 ( .A(n331), .B(n58), .Z(\ab[26][8] ) );
  AN2P U2838 ( .A(n327), .B(n58), .Z(\ab[26][7] ) );
  AN2P U2839 ( .A(n323), .B(n59), .Z(\ab[26][6] ) );
  AN2P U2840 ( .A(n319), .B(n59), .Z(\ab[26][5] ) );
  AN2P U2841 ( .A(n315), .B(n59), .Z(\ab[26][4] ) );
  AN2P U2842 ( .A(n311), .B(n59), .Z(\ab[26][3] ) );
  AN2P U2843 ( .A(n307), .B(n59), .Z(\ab[26][2] ) );
  AN2P U2844 ( .A(n303), .B(n59), .Z(\ab[26][1] ) );
  AN2P U2845 ( .A(n299), .B(n59), .Z(\ab[26][0] ) );
  AN2P U2846 ( .A(n451), .B(n44), .Z(\ab[27][38] ) );
  AN2P U2847 ( .A(n447), .B(n44), .Z(\ab[27][37] ) );
  AN2P U2848 ( .A(n443), .B(n44), .Z(\ab[27][36] ) );
  AN2P U2849 ( .A(n439), .B(n44), .Z(\ab[27][35] ) );
  AN2P U2850 ( .A(n435), .B(n44), .Z(\ab[27][34] ) );
  AN2P U2851 ( .A(n431), .B(n44), .Z(\ab[27][33] ) );
  AN2P U2852 ( .A(n427), .B(n44), .Z(\ab[27][32] ) );
  AN2P U2853 ( .A(n423), .B(n44), .Z(\ab[27][31] ) );
  AN2P U2854 ( .A(n419), .B(n45), .Z(\ab[27][30] ) );
  AN2P U2855 ( .A(n415), .B(n45), .Z(\ab[27][29] ) );
  AN2P U2856 ( .A(n411), .B(n45), .Z(\ab[27][28] ) );
  AN2P U2857 ( .A(n407), .B(n45), .Z(\ab[27][27] ) );
  AN2P U2858 ( .A(n403), .B(n45), .Z(\ab[27][26] ) );
  AN2P U2859 ( .A(n399), .B(n45), .Z(\ab[27][25] ) );
  AN2P U2860 ( .A(n395), .B(n45), .Z(\ab[27][24] ) );
  AN2P U2861 ( .A(n391), .B(n45), .Z(\ab[27][23] ) );
  AN2P U2862 ( .A(n387), .B(n46), .Z(\ab[27][22] ) );
  AN2P U2863 ( .A(n383), .B(n46), .Z(\ab[27][21] ) );
  AN2P U2864 ( .A(n379), .B(n46), .Z(\ab[27][20] ) );
  AN2P U2865 ( .A(n375), .B(n46), .Z(\ab[27][19] ) );
  AN2P U2866 ( .A(n371), .B(n46), .Z(\ab[27][18] ) );
  AN2P U2867 ( .A(n367), .B(n46), .Z(\ab[27][17] ) );
  AN2P U2868 ( .A(n363), .B(n46), .Z(\ab[27][16] ) );
  AN2P U2869 ( .A(n359), .B(n46), .Z(\ab[27][15] ) );
  AN2P U2870 ( .A(n355), .B(n47), .Z(\ab[27][14] ) );
  AN2P U2871 ( .A(n351), .B(n47), .Z(\ab[27][13] ) );
  AN2P U2872 ( .A(n347), .B(n47), .Z(\ab[27][12] ) );
  AN2P U2873 ( .A(n343), .B(n47), .Z(\ab[27][11] ) );
  AN2P U2874 ( .A(n339), .B(n47), .Z(\ab[27][10] ) );
  AN2P U2875 ( .A(n335), .B(n47), .Z(\ab[27][9] ) );
  AN2P U2876 ( .A(n331), .B(n47), .Z(\ab[27][8] ) );
  AN2P U2877 ( .A(n327), .B(n47), .Z(\ab[27][7] ) );
  AN2P U2878 ( .A(n323), .B(n48), .Z(\ab[27][6] ) );
  AN2P U2879 ( .A(n319), .B(n48), .Z(\ab[27][5] ) );
  AN2P U2880 ( .A(n315), .B(n48), .Z(\ab[27][4] ) );
  AN2P U2881 ( .A(n311), .B(n48), .Z(\ab[27][3] ) );
  AN2P U2882 ( .A(n307), .B(n48), .Z(\ab[27][2] ) );
  AN2P U2883 ( .A(n303), .B(n48), .Z(\ab[27][1] ) );
  AN2P U2884 ( .A(n299), .B(n48), .Z(\ab[27][0] ) );
  AN2P U2885 ( .A(n451), .B(n33), .Z(\ab[28][38] ) );
  AN2P U2886 ( .A(n447), .B(n33), .Z(\ab[28][37] ) );
  AN2P U2887 ( .A(n443), .B(n33), .Z(\ab[28][36] ) );
  AN2P U2888 ( .A(n439), .B(n33), .Z(\ab[28][35] ) );
  AN2P U2889 ( .A(n435), .B(n33), .Z(\ab[28][34] ) );
  AN2P U2890 ( .A(n431), .B(n33), .Z(\ab[28][33] ) );
  AN2P U2891 ( .A(n427), .B(n33), .Z(\ab[28][32] ) );
  AN2P U2892 ( .A(n423), .B(n33), .Z(\ab[28][31] ) );
  AN2P U2893 ( .A(n419), .B(n34), .Z(\ab[28][30] ) );
  AN2P U2894 ( .A(n415), .B(n34), .Z(\ab[28][29] ) );
  AN2P U2895 ( .A(n411), .B(n34), .Z(\ab[28][28] ) );
  AN2P U2896 ( .A(n407), .B(n34), .Z(\ab[28][27] ) );
  AN2P U2897 ( .A(n403), .B(n34), .Z(\ab[28][26] ) );
  AN2P U2898 ( .A(n399), .B(n34), .Z(\ab[28][25] ) );
  AN2P U2899 ( .A(n395), .B(n34), .Z(\ab[28][24] ) );
  AN2P U2900 ( .A(n391), .B(n34), .Z(\ab[28][23] ) );
  AN2P U2901 ( .A(n387), .B(n35), .Z(\ab[28][22] ) );
  AN2P U2902 ( .A(n383), .B(n35), .Z(\ab[28][21] ) );
  AN2P U2903 ( .A(n379), .B(n35), .Z(\ab[28][20] ) );
  AN2P U2904 ( .A(n375), .B(n35), .Z(\ab[28][19] ) );
  AN2P U2905 ( .A(n371), .B(n35), .Z(\ab[28][18] ) );
  AN2P U2906 ( .A(n367), .B(n35), .Z(\ab[28][17] ) );
  AN2P U2907 ( .A(n363), .B(n35), .Z(\ab[28][16] ) );
  AN2P U2908 ( .A(n359), .B(n35), .Z(\ab[28][15] ) );
  AN2P U2909 ( .A(n355), .B(n36), .Z(\ab[28][14] ) );
  AN2P U2910 ( .A(n351), .B(n36), .Z(\ab[28][13] ) );
  AN2P U2911 ( .A(n347), .B(n36), .Z(\ab[28][12] ) );
  AN2P U2912 ( .A(n343), .B(n36), .Z(\ab[28][11] ) );
  AN2P U2913 ( .A(n339), .B(n36), .Z(\ab[28][10] ) );
  AN2P U2914 ( .A(n335), .B(n36), .Z(\ab[28][9] ) );
  AN2P U2915 ( .A(n331), .B(n36), .Z(\ab[28][8] ) );
  AN2P U2916 ( .A(n327), .B(n36), .Z(\ab[28][7] ) );
  AN2P U2917 ( .A(n323), .B(n37), .Z(\ab[28][6] ) );
  AN2P U2918 ( .A(n319), .B(n37), .Z(\ab[28][5] ) );
  AN2P U2919 ( .A(n315), .B(n37), .Z(\ab[28][4] ) );
  AN2P U2920 ( .A(n311), .B(n37), .Z(\ab[28][3] ) );
  AN2P U2921 ( .A(n307), .B(n37), .Z(\ab[28][2] ) );
  AN2P U2922 ( .A(n303), .B(n37), .Z(\ab[28][1] ) );
  AN2P U2923 ( .A(n299), .B(n37), .Z(\ab[28][0] ) );
  AN2P U2924 ( .A(n451), .B(n22), .Z(\ab[29][38] ) );
  AN2P U2925 ( .A(n447), .B(n22), .Z(\ab[29][37] ) );
  AN2P U2926 ( .A(n443), .B(n22), .Z(\ab[29][36] ) );
  AN2P U2927 ( .A(n439), .B(n22), .Z(\ab[29][35] ) );
  AN2P U2928 ( .A(n435), .B(n22), .Z(\ab[29][34] ) );
  AN2P U2929 ( .A(n431), .B(n22), .Z(\ab[29][33] ) );
  AN2P U2930 ( .A(n427), .B(n22), .Z(\ab[29][32] ) );
  AN2P U2931 ( .A(n423), .B(n22), .Z(\ab[29][31] ) );
  AN2P U2932 ( .A(n419), .B(n23), .Z(\ab[29][30] ) );
  AN2P U2933 ( .A(n415), .B(n23), .Z(\ab[29][29] ) );
  AN2P U2934 ( .A(n411), .B(n23), .Z(\ab[29][28] ) );
  AN2P U2935 ( .A(n407), .B(n23), .Z(\ab[29][27] ) );
  AN2P U2936 ( .A(n403), .B(n23), .Z(\ab[29][26] ) );
  AN2P U2937 ( .A(n399), .B(n23), .Z(\ab[29][25] ) );
  AN2P U2938 ( .A(n395), .B(n23), .Z(\ab[29][24] ) );
  AN2P U2939 ( .A(n391), .B(n23), .Z(\ab[29][23] ) );
  AN2P U2940 ( .A(n387), .B(n24), .Z(\ab[29][22] ) );
  AN2P U2941 ( .A(n383), .B(n24), .Z(\ab[29][21] ) );
  AN2P U2942 ( .A(n379), .B(n24), .Z(\ab[29][20] ) );
  AN2P U2943 ( .A(n375), .B(n24), .Z(\ab[29][19] ) );
  AN2P U2944 ( .A(n371), .B(n24), .Z(\ab[29][18] ) );
  AN2P U2945 ( .A(n367), .B(n24), .Z(\ab[29][17] ) );
  AN2P U2946 ( .A(n363), .B(n24), .Z(\ab[29][16] ) );
  AN2P U2947 ( .A(n359), .B(n24), .Z(\ab[29][15] ) );
  AN2P U2948 ( .A(n355), .B(n25), .Z(\ab[29][14] ) );
  AN2P U2949 ( .A(n351), .B(n25), .Z(\ab[29][13] ) );
  AN2P U2950 ( .A(n347), .B(n25), .Z(\ab[29][12] ) );
  AN2P U2951 ( .A(n343), .B(n25), .Z(\ab[29][11] ) );
  AN2P U2952 ( .A(n339), .B(n25), .Z(\ab[29][10] ) );
  AN2P U2953 ( .A(n335), .B(n25), .Z(\ab[29][9] ) );
  AN2P U2954 ( .A(n331), .B(n25), .Z(\ab[29][8] ) );
  AN2P U2955 ( .A(n327), .B(n25), .Z(\ab[29][7] ) );
  AN2P U2956 ( .A(n323), .B(n26), .Z(\ab[29][6] ) );
  AN2P U2957 ( .A(n319), .B(n26), .Z(\ab[29][5] ) );
  AN2P U2958 ( .A(n315), .B(n26), .Z(\ab[29][4] ) );
  AN2P U2959 ( .A(n311), .B(n26), .Z(\ab[29][3] ) );
  AN2P U2960 ( .A(n307), .B(n26), .Z(\ab[29][2] ) );
  AN2P U2961 ( .A(n303), .B(n26), .Z(\ab[29][1] ) );
  AN2P U2962 ( .A(n299), .B(n26), .Z(\ab[29][0] ) );
  NR2 U2964 ( .A(n492), .B(n16), .Z(\ab[29][95] ) );
  NR2 U2965 ( .A(n493), .B(n16), .Z(\ab[29][94] ) );
  NR2 U2966 ( .A(n494), .B(n16), .Z(\ab[29][93] ) );
  NR2 U2967 ( .A(n495), .B(n16), .Z(\ab[29][92] ) );
  NR2 U2968 ( .A(n496), .B(n16), .Z(\ab[29][91] ) );
  NR2 U2969 ( .A(n497), .B(n16), .Z(\ab[29][90] ) );
  NR2 U2970 ( .A(n498), .B(n16), .Z(\ab[29][89] ) );
  NR2 U2971 ( .A(n499), .B(n16), .Z(\ab[29][88] ) );
  NR2 U2972 ( .A(n500), .B(n16), .Z(\ab[29][87] ) );
  NR2 U2973 ( .A(n501), .B(n16), .Z(\ab[29][86] ) );
  NR2 U2974 ( .A(n502), .B(n16), .Z(\ab[29][85] ) );
  NR2 U2975 ( .A(n503), .B(n16), .Z(\ab[29][84] ) );
  NR2 U2976 ( .A(n504), .B(n17), .Z(\ab[29][83] ) );
  NR2 U2977 ( .A(n505), .B(n17), .Z(\ab[29][82] ) );
  NR2 U2978 ( .A(n506), .B(n17), .Z(\ab[29][81] ) );
  NR2 U2979 ( .A(n507), .B(n17), .Z(\ab[29][80] ) );
  NR2 U2980 ( .A(n508), .B(n17), .Z(\ab[29][79] ) );
  NR2 U2981 ( .A(n509), .B(n17), .Z(\ab[29][78] ) );
  NR2 U2982 ( .A(n510), .B(n17), .Z(\ab[29][77] ) );
  NR2 U2983 ( .A(n511), .B(n17), .Z(\ab[29][76] ) );
  NR2 U2984 ( .A(n512), .B(n17), .Z(\ab[29][75] ) );
  NR2 U2985 ( .A(n513), .B(n17), .Z(\ab[29][74] ) );
  NR2 U2986 ( .A(n514), .B(n17), .Z(\ab[29][73] ) );
  NR2 U2987 ( .A(n515), .B(n17), .Z(\ab[29][72] ) );
  NR2 U2988 ( .A(n516), .B(n18), .Z(\ab[29][71] ) );
  NR2 U2989 ( .A(n517), .B(n18), .Z(\ab[29][70] ) );
  NR2 U2990 ( .A(n518), .B(n18), .Z(\ab[29][69] ) );
  NR2 U2991 ( .A(n519), .B(n18), .Z(\ab[29][68] ) );
  NR2 U2992 ( .A(n520), .B(n18), .Z(\ab[29][67] ) );
  NR2 U2993 ( .A(n521), .B(n18), .Z(\ab[29][66] ) );
  NR2 U2994 ( .A(n522), .B(n18), .Z(\ab[29][65] ) );
  NR2 U2995 ( .A(n523), .B(n18), .Z(\ab[29][64] ) );
  NR2 U2996 ( .A(n524), .B(n18), .Z(\ab[29][63] ) );
  NR2 U2997 ( .A(n525), .B(n18), .Z(\ab[29][62] ) );
  NR2 U2998 ( .A(n526), .B(n18), .Z(\ab[29][61] ) );
  NR2 U2999 ( .A(n527), .B(n18), .Z(\ab[29][60] ) );
  NR2 U3000 ( .A(n528), .B(n19), .Z(\ab[29][59] ) );
  NR2 U3001 ( .A(n529), .B(n19), .Z(\ab[29][58] ) );
  NR2 U3002 ( .A(n530), .B(n19), .Z(\ab[29][57] ) );
  NR2 U3003 ( .A(n531), .B(n19), .Z(\ab[29][56] ) );
  NR2 U3004 ( .A(n532), .B(n19), .Z(\ab[29][55] ) );
  NR2 U3005 ( .A(n533), .B(n19), .Z(\ab[29][54] ) );
  NR2 U3006 ( .A(n534), .B(n19), .Z(\ab[29][53] ) );
  NR2 U3007 ( .A(n535), .B(n19), .Z(\ab[29][52] ) );
  NR2 U3008 ( .A(n536), .B(n19), .Z(\ab[29][51] ) );
  NR2 U3009 ( .A(n537), .B(n19), .Z(\ab[29][50] ) );
  NR2 U3010 ( .A(n538), .B(n19), .Z(\ab[29][49] ) );
  NR2 U3011 ( .A(n539), .B(n19), .Z(\ab[29][48] ) );
  NR2 U3012 ( .A(n540), .B(n20), .Z(\ab[29][47] ) );
  NR2 U3013 ( .A(n541), .B(n20), .Z(\ab[29][46] ) );
  NR2 U3014 ( .A(n542), .B(n20), .Z(\ab[29][45] ) );
  NR2 U3015 ( .A(n543), .B(n20), .Z(\ab[29][44] ) );
  NR2 U3016 ( .A(n544), .B(n20), .Z(\ab[29][43] ) );
  NR2 U3017 ( .A(n545), .B(n20), .Z(\ab[29][42] ) );
  NR2 U3018 ( .A(n546), .B(n20), .Z(\ab[29][41] ) );
  NR2 U3019 ( .A(n547), .B(n20), .Z(\ab[29][40] ) );
  NR2 U3020 ( .A(n548), .B(n20), .Z(\ab[29][39] ) );
  NR2 U3021 ( .A(n492), .B(n27), .Z(\ab[28][95] ) );
  NR2 U3022 ( .A(n493), .B(n27), .Z(\ab[28][94] ) );
  NR2 U3023 ( .A(n494), .B(n27), .Z(\ab[28][93] ) );
  NR2 U3024 ( .A(n495), .B(n27), .Z(\ab[28][92] ) );
  NR2 U3025 ( .A(n496), .B(n27), .Z(\ab[28][91] ) );
  NR2 U3026 ( .A(n497), .B(n27), .Z(\ab[28][90] ) );
  NR2 U3027 ( .A(n498), .B(n27), .Z(\ab[28][89] ) );
  NR2 U3028 ( .A(n499), .B(n27), .Z(\ab[28][88] ) );
  NR2 U3029 ( .A(n500), .B(n27), .Z(\ab[28][87] ) );
  NR2 U3030 ( .A(n501), .B(n27), .Z(\ab[28][86] ) );
  NR2 U3031 ( .A(n502), .B(n27), .Z(\ab[28][85] ) );
  NR2 U3032 ( .A(n503), .B(n27), .Z(\ab[28][84] ) );
  NR2 U3033 ( .A(n504), .B(n28), .Z(\ab[28][83] ) );
  NR2 U3034 ( .A(n505), .B(n28), .Z(\ab[28][82] ) );
  NR2 U3035 ( .A(n506), .B(n28), .Z(\ab[28][81] ) );
  NR2 U3036 ( .A(n507), .B(n28), .Z(\ab[28][80] ) );
  NR2 U3037 ( .A(n508), .B(n28), .Z(\ab[28][79] ) );
  NR2 U3038 ( .A(n509), .B(n28), .Z(\ab[28][78] ) );
  NR2 U3039 ( .A(n510), .B(n28), .Z(\ab[28][77] ) );
  NR2 U3040 ( .A(n511), .B(n28), .Z(\ab[28][76] ) );
  NR2 U3041 ( .A(n512), .B(n28), .Z(\ab[28][75] ) );
  NR2 U3042 ( .A(n513), .B(n28), .Z(\ab[28][74] ) );
  NR2 U3043 ( .A(n514), .B(n28), .Z(\ab[28][73] ) );
  NR2 U3044 ( .A(n515), .B(n28), .Z(\ab[28][72] ) );
  NR2 U3045 ( .A(n516), .B(n29), .Z(\ab[28][71] ) );
  NR2 U3046 ( .A(n517), .B(n29), .Z(\ab[28][70] ) );
  NR2 U3047 ( .A(n518), .B(n29), .Z(\ab[28][69] ) );
  NR2 U3048 ( .A(n519), .B(n29), .Z(\ab[28][68] ) );
  NR2 U3049 ( .A(n520), .B(n29), .Z(\ab[28][67] ) );
  NR2 U3050 ( .A(n521), .B(n29), .Z(\ab[28][66] ) );
  NR2 U3051 ( .A(n522), .B(n29), .Z(\ab[28][65] ) );
  NR2 U3052 ( .A(n523), .B(n29), .Z(\ab[28][64] ) );
  NR2 U3053 ( .A(n524), .B(n29), .Z(\ab[28][63] ) );
  NR2 U3054 ( .A(n525), .B(n29), .Z(\ab[28][62] ) );
  NR2 U3055 ( .A(n526), .B(n29), .Z(\ab[28][61] ) );
  NR2 U3056 ( .A(n527), .B(n29), .Z(\ab[28][60] ) );
  NR2 U3057 ( .A(n528), .B(n30), .Z(\ab[28][59] ) );
  NR2 U3058 ( .A(n529), .B(n30), .Z(\ab[28][58] ) );
  NR2 U3059 ( .A(n530), .B(n30), .Z(\ab[28][57] ) );
  NR2 U3060 ( .A(n531), .B(n30), .Z(\ab[28][56] ) );
  NR2 U3061 ( .A(n532), .B(n30), .Z(\ab[28][55] ) );
  NR2 U3062 ( .A(n533), .B(n30), .Z(\ab[28][54] ) );
  NR2 U3063 ( .A(n534), .B(n30), .Z(\ab[28][53] ) );
  NR2 U3064 ( .A(n535), .B(n30), .Z(\ab[28][52] ) );
  NR2 U3065 ( .A(n536), .B(n30), .Z(\ab[28][51] ) );
  NR2 U3066 ( .A(n537), .B(n30), .Z(\ab[28][50] ) );
  NR2 U3067 ( .A(n538), .B(n30), .Z(\ab[28][49] ) );
  NR2 U3068 ( .A(n539), .B(n30), .Z(\ab[28][48] ) );
  NR2 U3069 ( .A(n540), .B(n31), .Z(\ab[28][47] ) );
  NR2 U3070 ( .A(n541), .B(n31), .Z(\ab[28][46] ) );
  NR2 U3071 ( .A(n542), .B(n31), .Z(\ab[28][45] ) );
  NR2 U3072 ( .A(n543), .B(n31), .Z(\ab[28][44] ) );
  NR2 U3073 ( .A(n544), .B(n31), .Z(\ab[28][43] ) );
  NR2 U3074 ( .A(n545), .B(n31), .Z(\ab[28][42] ) );
  NR2 U3075 ( .A(n546), .B(n31), .Z(\ab[28][41] ) );
  NR2 U3076 ( .A(n547), .B(n31), .Z(\ab[28][40] ) );
  NR2 U3077 ( .A(n548), .B(n31), .Z(\ab[28][39] ) );
  NR2 U3078 ( .A(n492), .B(n38), .Z(\ab[27][95] ) );
  NR2 U3079 ( .A(n493), .B(n38), .Z(\ab[27][94] ) );
  NR2 U3080 ( .A(n494), .B(n38), .Z(\ab[27][93] ) );
  NR2 U3081 ( .A(n495), .B(n38), .Z(\ab[27][92] ) );
  NR2 U3082 ( .A(n496), .B(n38), .Z(\ab[27][91] ) );
  NR2 U3083 ( .A(n497), .B(n38), .Z(\ab[27][90] ) );
  NR2 U3084 ( .A(n498), .B(n38), .Z(\ab[27][89] ) );
  NR2 U3085 ( .A(n499), .B(n38), .Z(\ab[27][88] ) );
  NR2 U3086 ( .A(n500), .B(n38), .Z(\ab[27][87] ) );
  NR2 U3087 ( .A(n501), .B(n38), .Z(\ab[27][86] ) );
  NR2 U3088 ( .A(n502), .B(n38), .Z(\ab[27][85] ) );
  NR2 U3089 ( .A(n503), .B(n38), .Z(\ab[27][84] ) );
  NR2 U3090 ( .A(n504), .B(n39), .Z(\ab[27][83] ) );
  NR2 U3091 ( .A(n505), .B(n39), .Z(\ab[27][82] ) );
  NR2 U3092 ( .A(n506), .B(n39), .Z(\ab[27][81] ) );
  NR2 U3093 ( .A(n507), .B(n39), .Z(\ab[27][80] ) );
  NR2 U3094 ( .A(n508), .B(n39), .Z(\ab[27][79] ) );
  NR2 U3095 ( .A(n509), .B(n39), .Z(\ab[27][78] ) );
  NR2 U3096 ( .A(n510), .B(n39), .Z(\ab[27][77] ) );
  NR2 U3097 ( .A(n511), .B(n39), .Z(\ab[27][76] ) );
  NR2 U3098 ( .A(n512), .B(n39), .Z(\ab[27][75] ) );
  NR2 U3099 ( .A(n513), .B(n39), .Z(\ab[27][74] ) );
  NR2 U3100 ( .A(n514), .B(n39), .Z(\ab[27][73] ) );
  NR2 U3101 ( .A(n515), .B(n39), .Z(\ab[27][72] ) );
  NR2 U3102 ( .A(n516), .B(n40), .Z(\ab[27][71] ) );
  NR2 U3103 ( .A(n517), .B(n40), .Z(\ab[27][70] ) );
  NR2 U3104 ( .A(n518), .B(n40), .Z(\ab[27][69] ) );
  NR2 U3105 ( .A(n519), .B(n40), .Z(\ab[27][68] ) );
  NR2 U3106 ( .A(n520), .B(n40), .Z(\ab[27][67] ) );
  NR2 U3107 ( .A(n521), .B(n40), .Z(\ab[27][66] ) );
  NR2 U3108 ( .A(n522), .B(n40), .Z(\ab[27][65] ) );
  NR2 U3109 ( .A(n523), .B(n40), .Z(\ab[27][64] ) );
  NR2 U3110 ( .A(n524), .B(n40), .Z(\ab[27][63] ) );
  NR2 U3111 ( .A(n525), .B(n40), .Z(\ab[27][62] ) );
  NR2 U3112 ( .A(n526), .B(n40), .Z(\ab[27][61] ) );
  NR2 U3113 ( .A(n527), .B(n40), .Z(\ab[27][60] ) );
  NR2 U3114 ( .A(n528), .B(n41), .Z(\ab[27][59] ) );
  NR2 U3115 ( .A(n529), .B(n41), .Z(\ab[27][58] ) );
  NR2 U3116 ( .A(n530), .B(n41), .Z(\ab[27][57] ) );
  NR2 U3117 ( .A(n531), .B(n41), .Z(\ab[27][56] ) );
  NR2 U3118 ( .A(n532), .B(n41), .Z(\ab[27][55] ) );
  NR2 U3119 ( .A(n533), .B(n41), .Z(\ab[27][54] ) );
  NR2 U3120 ( .A(n534), .B(n41), .Z(\ab[27][53] ) );
  NR2 U3121 ( .A(n535), .B(n41), .Z(\ab[27][52] ) );
  NR2 U3122 ( .A(n536), .B(n41), .Z(\ab[27][51] ) );
  NR2 U3123 ( .A(n537), .B(n41), .Z(\ab[27][50] ) );
  NR2 U3124 ( .A(n538), .B(n41), .Z(\ab[27][49] ) );
  NR2 U3125 ( .A(n539), .B(n41), .Z(\ab[27][48] ) );
  NR2 U3126 ( .A(n540), .B(n42), .Z(\ab[27][47] ) );
  NR2 U3127 ( .A(n541), .B(n42), .Z(\ab[27][46] ) );
  NR2 U3128 ( .A(n542), .B(n42), .Z(\ab[27][45] ) );
  NR2 U3129 ( .A(n543), .B(n42), .Z(\ab[27][44] ) );
  NR2 U3130 ( .A(n544), .B(n42), .Z(\ab[27][43] ) );
  NR2 U3131 ( .A(n545), .B(n42), .Z(\ab[27][42] ) );
  NR2 U3132 ( .A(n546), .B(n42), .Z(\ab[27][41] ) );
  NR2 U3133 ( .A(n547), .B(n42), .Z(\ab[27][40] ) );
  NR2 U3134 ( .A(n548), .B(n42), .Z(\ab[27][39] ) );
  NR2 U3135 ( .A(n492), .B(n49), .Z(\ab[26][95] ) );
  NR2 U3136 ( .A(n493), .B(n49), .Z(\ab[26][94] ) );
  NR2 U3137 ( .A(n494), .B(n49), .Z(\ab[26][93] ) );
  NR2 U3138 ( .A(n495), .B(n49), .Z(\ab[26][92] ) );
  NR2 U3139 ( .A(n496), .B(n49), .Z(\ab[26][91] ) );
  NR2 U3140 ( .A(n497), .B(n49), .Z(\ab[26][90] ) );
  NR2 U3141 ( .A(n498), .B(n49), .Z(\ab[26][89] ) );
  NR2 U3142 ( .A(n499), .B(n49), .Z(\ab[26][88] ) );
  NR2 U3143 ( .A(n500), .B(n49), .Z(\ab[26][87] ) );
  NR2 U3144 ( .A(n501), .B(n49), .Z(\ab[26][86] ) );
  NR2 U3145 ( .A(n502), .B(n49), .Z(\ab[26][85] ) );
  NR2 U3146 ( .A(n503), .B(n49), .Z(\ab[26][84] ) );
  NR2 U3147 ( .A(n504), .B(n50), .Z(\ab[26][83] ) );
  NR2 U3148 ( .A(n505), .B(n50), .Z(\ab[26][82] ) );
  NR2 U3149 ( .A(n506), .B(n50), .Z(\ab[26][81] ) );
  NR2 U3150 ( .A(n507), .B(n50), .Z(\ab[26][80] ) );
  NR2 U3151 ( .A(n508), .B(n50), .Z(\ab[26][79] ) );
  NR2 U3152 ( .A(n509), .B(n50), .Z(\ab[26][78] ) );
  NR2 U3153 ( .A(n510), .B(n50), .Z(\ab[26][77] ) );
  NR2 U3154 ( .A(n511), .B(n50), .Z(\ab[26][76] ) );
  NR2 U3155 ( .A(n512), .B(n50), .Z(\ab[26][75] ) );
  NR2 U3156 ( .A(n513), .B(n50), .Z(\ab[26][74] ) );
  NR2 U3157 ( .A(n514), .B(n50), .Z(\ab[26][73] ) );
  NR2 U3158 ( .A(n515), .B(n50), .Z(\ab[26][72] ) );
  NR2 U3159 ( .A(n516), .B(n51), .Z(\ab[26][71] ) );
  NR2 U3160 ( .A(n517), .B(n51), .Z(\ab[26][70] ) );
  NR2 U3161 ( .A(n518), .B(n51), .Z(\ab[26][69] ) );
  NR2 U3162 ( .A(n519), .B(n51), .Z(\ab[26][68] ) );
  NR2 U3163 ( .A(n520), .B(n51), .Z(\ab[26][67] ) );
  NR2 U3164 ( .A(n521), .B(n51), .Z(\ab[26][66] ) );
  NR2 U3165 ( .A(n522), .B(n51), .Z(\ab[26][65] ) );
  NR2 U3166 ( .A(n523), .B(n51), .Z(\ab[26][64] ) );
  NR2 U3167 ( .A(n524), .B(n51), .Z(\ab[26][63] ) );
  NR2 U3168 ( .A(n525), .B(n51), .Z(\ab[26][62] ) );
  NR2 U3169 ( .A(n526), .B(n51), .Z(\ab[26][61] ) );
  NR2 U3170 ( .A(n527), .B(n51), .Z(\ab[26][60] ) );
  NR2 U3171 ( .A(n528), .B(n52), .Z(\ab[26][59] ) );
  NR2 U3172 ( .A(n529), .B(n52), .Z(\ab[26][58] ) );
  NR2 U3173 ( .A(n530), .B(n52), .Z(\ab[26][57] ) );
  NR2 U3174 ( .A(n531), .B(n52), .Z(\ab[26][56] ) );
  NR2 U3175 ( .A(n532), .B(n52), .Z(\ab[26][55] ) );
  NR2 U3176 ( .A(n533), .B(n52), .Z(\ab[26][54] ) );
  NR2 U3177 ( .A(n534), .B(n52), .Z(\ab[26][53] ) );
  NR2 U3178 ( .A(n535), .B(n52), .Z(\ab[26][52] ) );
  NR2 U3179 ( .A(n536), .B(n52), .Z(\ab[26][51] ) );
  NR2 U3180 ( .A(n537), .B(n52), .Z(\ab[26][50] ) );
  NR2 U3181 ( .A(n538), .B(n52), .Z(\ab[26][49] ) );
  NR2 U3182 ( .A(n539), .B(n52), .Z(\ab[26][48] ) );
  NR2 U3183 ( .A(n540), .B(n53), .Z(\ab[26][47] ) );
  NR2 U3184 ( .A(n541), .B(n53), .Z(\ab[26][46] ) );
  NR2 U3185 ( .A(n542), .B(n53), .Z(\ab[26][45] ) );
  NR2 U3186 ( .A(n543), .B(n53), .Z(\ab[26][44] ) );
  NR2 U3187 ( .A(n544), .B(n53), .Z(\ab[26][43] ) );
  NR2 U3188 ( .A(n545), .B(n53), .Z(\ab[26][42] ) );
  NR2 U3189 ( .A(n546), .B(n53), .Z(\ab[26][41] ) );
  NR2 U3190 ( .A(n547), .B(n53), .Z(\ab[26][40] ) );
  NR2 U3191 ( .A(n548), .B(n53), .Z(\ab[26][39] ) );
  NR2 U3192 ( .A(n492), .B(n60), .Z(\ab[25][95] ) );
  NR2 U3193 ( .A(n493), .B(n60), .Z(\ab[25][94] ) );
  NR2 U3194 ( .A(n494), .B(n60), .Z(\ab[25][93] ) );
  NR2 U3195 ( .A(n495), .B(n60), .Z(\ab[25][92] ) );
  NR2 U3196 ( .A(n496), .B(n60), .Z(\ab[25][91] ) );
  NR2 U3197 ( .A(n497), .B(n60), .Z(\ab[25][90] ) );
  NR2 U3198 ( .A(n498), .B(n60), .Z(\ab[25][89] ) );
  NR2 U3199 ( .A(n499), .B(n60), .Z(\ab[25][88] ) );
  NR2 U3200 ( .A(n500), .B(n60), .Z(\ab[25][87] ) );
  NR2 U3201 ( .A(n501), .B(n60), .Z(\ab[25][86] ) );
  NR2 U3202 ( .A(n502), .B(n60), .Z(\ab[25][85] ) );
  NR2 U3203 ( .A(n503), .B(n60), .Z(\ab[25][84] ) );
  NR2 U3204 ( .A(n504), .B(n61), .Z(\ab[25][83] ) );
  NR2 U3205 ( .A(n505), .B(n61), .Z(\ab[25][82] ) );
  NR2 U3206 ( .A(n506), .B(n61), .Z(\ab[25][81] ) );
  NR2 U3207 ( .A(n507), .B(n61), .Z(\ab[25][80] ) );
  NR2 U3208 ( .A(n508), .B(n61), .Z(\ab[25][79] ) );
  NR2 U3209 ( .A(n509), .B(n61), .Z(\ab[25][78] ) );
  NR2 U3210 ( .A(n510), .B(n61), .Z(\ab[25][77] ) );
  NR2 U3211 ( .A(n511), .B(n61), .Z(\ab[25][76] ) );
  NR2 U3212 ( .A(n512), .B(n61), .Z(\ab[25][75] ) );
  NR2 U3213 ( .A(n513), .B(n61), .Z(\ab[25][74] ) );
  NR2 U3214 ( .A(n514), .B(n61), .Z(\ab[25][73] ) );
  NR2 U3215 ( .A(n515), .B(n61), .Z(\ab[25][72] ) );
  NR2 U3216 ( .A(n516), .B(n62), .Z(\ab[25][71] ) );
  NR2 U3217 ( .A(n517), .B(n62), .Z(\ab[25][70] ) );
  NR2 U3218 ( .A(n518), .B(n62), .Z(\ab[25][69] ) );
  NR2 U3219 ( .A(n519), .B(n62), .Z(\ab[25][68] ) );
  NR2 U3220 ( .A(n520), .B(n62), .Z(\ab[25][67] ) );
  NR2 U3221 ( .A(n521), .B(n62), .Z(\ab[25][66] ) );
  NR2 U3222 ( .A(n522), .B(n62), .Z(\ab[25][65] ) );
  NR2 U3223 ( .A(n523), .B(n62), .Z(\ab[25][64] ) );
  NR2 U3224 ( .A(n524), .B(n62), .Z(\ab[25][63] ) );
  NR2 U3225 ( .A(n525), .B(n62), .Z(\ab[25][62] ) );
  NR2 U3226 ( .A(n526), .B(n62), .Z(\ab[25][61] ) );
  NR2 U3227 ( .A(n527), .B(n62), .Z(\ab[25][60] ) );
  NR2 U3228 ( .A(n528), .B(n63), .Z(\ab[25][59] ) );
  NR2 U3229 ( .A(n529), .B(n63), .Z(\ab[25][58] ) );
  NR2 U3230 ( .A(n530), .B(n63), .Z(\ab[25][57] ) );
  NR2 U3231 ( .A(n531), .B(n63), .Z(\ab[25][56] ) );
  NR2 U3232 ( .A(n532), .B(n63), .Z(\ab[25][55] ) );
  NR2 U3233 ( .A(n533), .B(n63), .Z(\ab[25][54] ) );
  NR2 U3234 ( .A(n534), .B(n63), .Z(\ab[25][53] ) );
  NR2 U3235 ( .A(n535), .B(n63), .Z(\ab[25][52] ) );
  NR2 U3236 ( .A(n536), .B(n63), .Z(\ab[25][51] ) );
  NR2 U3237 ( .A(n537), .B(n63), .Z(\ab[25][50] ) );
  NR2 U3238 ( .A(n538), .B(n63), .Z(\ab[25][49] ) );
  NR2 U3239 ( .A(n539), .B(n63), .Z(\ab[25][48] ) );
  NR2 U3240 ( .A(n540), .B(n64), .Z(\ab[25][47] ) );
  NR2 U3241 ( .A(n541), .B(n64), .Z(\ab[25][46] ) );
  NR2 U3242 ( .A(n542), .B(n64), .Z(\ab[25][45] ) );
  NR2 U3243 ( .A(n543), .B(n64), .Z(\ab[25][44] ) );
  NR2 U3244 ( .A(n544), .B(n64), .Z(\ab[25][43] ) );
  NR2 U3245 ( .A(n545), .B(n64), .Z(\ab[25][42] ) );
  NR2 U3246 ( .A(n546), .B(n64), .Z(\ab[25][41] ) );
  NR2 U3247 ( .A(n547), .B(n64), .Z(\ab[25][40] ) );
  NR2 U3248 ( .A(n548), .B(n64), .Z(\ab[25][39] ) );
  NR2 U3249 ( .A(n492), .B(n71), .Z(\ab[24][95] ) );
  NR2 U3250 ( .A(n493), .B(n71), .Z(\ab[24][94] ) );
  NR2 U3251 ( .A(n494), .B(n71), .Z(\ab[24][93] ) );
  NR2 U3252 ( .A(n495), .B(n71), .Z(\ab[24][92] ) );
  NR2 U3253 ( .A(n496), .B(n71), .Z(\ab[24][91] ) );
  NR2 U3254 ( .A(n497), .B(n71), .Z(\ab[24][90] ) );
  NR2 U3255 ( .A(n498), .B(n71), .Z(\ab[24][89] ) );
  NR2 U3256 ( .A(n499), .B(n71), .Z(\ab[24][88] ) );
  NR2 U3257 ( .A(n500), .B(n71), .Z(\ab[24][87] ) );
  NR2 U3258 ( .A(n501), .B(n71), .Z(\ab[24][86] ) );
  NR2 U3259 ( .A(n502), .B(n71), .Z(\ab[24][85] ) );
  NR2 U3260 ( .A(n503), .B(n71), .Z(\ab[24][84] ) );
  NR2 U3261 ( .A(n504), .B(n72), .Z(\ab[24][83] ) );
  NR2 U3262 ( .A(n505), .B(n72), .Z(\ab[24][82] ) );
  NR2 U3263 ( .A(n506), .B(n72), .Z(\ab[24][81] ) );
  NR2 U3264 ( .A(n507), .B(n72), .Z(\ab[24][80] ) );
  NR2 U3265 ( .A(n508), .B(n72), .Z(\ab[24][79] ) );
  NR2 U3266 ( .A(n509), .B(n72), .Z(\ab[24][78] ) );
  NR2 U3267 ( .A(n510), .B(n72), .Z(\ab[24][77] ) );
  NR2 U3268 ( .A(n511), .B(n72), .Z(\ab[24][76] ) );
  NR2 U3269 ( .A(n512), .B(n72), .Z(\ab[24][75] ) );
  NR2 U3270 ( .A(n513), .B(n72), .Z(\ab[24][74] ) );
  NR2 U3271 ( .A(n514), .B(n72), .Z(\ab[24][73] ) );
  NR2 U3272 ( .A(n515), .B(n72), .Z(\ab[24][72] ) );
  NR2 U3273 ( .A(n516), .B(n73), .Z(\ab[24][71] ) );
  NR2 U3274 ( .A(n517), .B(n73), .Z(\ab[24][70] ) );
  NR2 U3275 ( .A(n518), .B(n73), .Z(\ab[24][69] ) );
  NR2 U3276 ( .A(n519), .B(n73), .Z(\ab[24][68] ) );
  NR2 U3277 ( .A(n520), .B(n73), .Z(\ab[24][67] ) );
  NR2 U3278 ( .A(n521), .B(n73), .Z(\ab[24][66] ) );
  NR2 U3279 ( .A(n522), .B(n73), .Z(\ab[24][65] ) );
  NR2 U3280 ( .A(n523), .B(n73), .Z(\ab[24][64] ) );
  NR2 U3281 ( .A(n524), .B(n73), .Z(\ab[24][63] ) );
  NR2 U3282 ( .A(n525), .B(n73), .Z(\ab[24][62] ) );
  NR2 U3283 ( .A(n526), .B(n73), .Z(\ab[24][61] ) );
  NR2 U3284 ( .A(n527), .B(n73), .Z(\ab[24][60] ) );
  NR2 U3285 ( .A(n528), .B(n74), .Z(\ab[24][59] ) );
  NR2 U3286 ( .A(n529), .B(n74), .Z(\ab[24][58] ) );
  NR2 U3287 ( .A(n530), .B(n74), .Z(\ab[24][57] ) );
  NR2 U3288 ( .A(n531), .B(n74), .Z(\ab[24][56] ) );
  NR2 U3289 ( .A(n532), .B(n74), .Z(\ab[24][55] ) );
  NR2 U3290 ( .A(n533), .B(n74), .Z(\ab[24][54] ) );
  NR2 U3291 ( .A(n534), .B(n74), .Z(\ab[24][53] ) );
  NR2 U3292 ( .A(n535), .B(n74), .Z(\ab[24][52] ) );
  NR2 U3293 ( .A(n536), .B(n74), .Z(\ab[24][51] ) );
  NR2 U3294 ( .A(n537), .B(n74), .Z(\ab[24][50] ) );
  NR2 U3295 ( .A(n538), .B(n74), .Z(\ab[24][49] ) );
  NR2 U3296 ( .A(n539), .B(n74), .Z(\ab[24][48] ) );
  NR2 U3297 ( .A(n540), .B(n75), .Z(\ab[24][47] ) );
  NR2 U3298 ( .A(n541), .B(n75), .Z(\ab[24][46] ) );
  NR2 U3299 ( .A(n542), .B(n75), .Z(\ab[24][45] ) );
  NR2 U3300 ( .A(n543), .B(n75), .Z(\ab[24][44] ) );
  NR2 U3301 ( .A(n544), .B(n75), .Z(\ab[24][43] ) );
  NR2 U3302 ( .A(n545), .B(n75), .Z(\ab[24][42] ) );
  NR2 U3303 ( .A(n546), .B(n75), .Z(\ab[24][41] ) );
  NR2 U3304 ( .A(n547), .B(n75), .Z(\ab[24][40] ) );
  NR2 U3305 ( .A(n548), .B(n75), .Z(\ab[24][39] ) );
  NR2 U3306 ( .A(n492), .B(n82), .Z(\ab[23][95] ) );
  NR2 U3307 ( .A(n493), .B(n82), .Z(\ab[23][94] ) );
  NR2 U3308 ( .A(n494), .B(n82), .Z(\ab[23][93] ) );
  NR2 U3309 ( .A(n495), .B(n82), .Z(\ab[23][92] ) );
  NR2 U3310 ( .A(n496), .B(n82), .Z(\ab[23][91] ) );
  NR2 U3311 ( .A(n497), .B(n82), .Z(\ab[23][90] ) );
  NR2 U3312 ( .A(n498), .B(n82), .Z(\ab[23][89] ) );
  NR2 U3313 ( .A(n499), .B(n82), .Z(\ab[23][88] ) );
  NR2 U3314 ( .A(n500), .B(n82), .Z(\ab[23][87] ) );
  NR2 U3315 ( .A(n501), .B(n82), .Z(\ab[23][86] ) );
  NR2 U3316 ( .A(n502), .B(n82), .Z(\ab[23][85] ) );
  NR2 U3317 ( .A(n503), .B(n82), .Z(\ab[23][84] ) );
  NR2 U3318 ( .A(n504), .B(n83), .Z(\ab[23][83] ) );
  NR2 U3319 ( .A(n505), .B(n83), .Z(\ab[23][82] ) );
  NR2 U3320 ( .A(n506), .B(n83), .Z(\ab[23][81] ) );
  NR2 U3321 ( .A(n507), .B(n83), .Z(\ab[23][80] ) );
  NR2 U3322 ( .A(n508), .B(n83), .Z(\ab[23][79] ) );
  NR2 U3323 ( .A(n509), .B(n83), .Z(\ab[23][78] ) );
  NR2 U3324 ( .A(n510), .B(n83), .Z(\ab[23][77] ) );
  NR2 U3325 ( .A(n511), .B(n83), .Z(\ab[23][76] ) );
  NR2 U3326 ( .A(n512), .B(n83), .Z(\ab[23][75] ) );
  NR2 U3327 ( .A(n513), .B(n83), .Z(\ab[23][74] ) );
  NR2 U3328 ( .A(n514), .B(n83), .Z(\ab[23][73] ) );
  NR2 U3329 ( .A(n515), .B(n83), .Z(\ab[23][72] ) );
  NR2 U3330 ( .A(n516), .B(n84), .Z(\ab[23][71] ) );
  NR2 U3331 ( .A(n517), .B(n84), .Z(\ab[23][70] ) );
  NR2 U3332 ( .A(n518), .B(n84), .Z(\ab[23][69] ) );
  NR2 U3333 ( .A(n519), .B(n84), .Z(\ab[23][68] ) );
  NR2 U3334 ( .A(n520), .B(n84), .Z(\ab[23][67] ) );
  NR2 U3335 ( .A(n521), .B(n84), .Z(\ab[23][66] ) );
  NR2 U3336 ( .A(n522), .B(n84), .Z(\ab[23][65] ) );
  NR2 U3337 ( .A(n523), .B(n84), .Z(\ab[23][64] ) );
  NR2 U3338 ( .A(n524), .B(n84), .Z(\ab[23][63] ) );
  NR2 U3339 ( .A(n525), .B(n84), .Z(\ab[23][62] ) );
  NR2 U3340 ( .A(n526), .B(n84), .Z(\ab[23][61] ) );
  NR2 U3341 ( .A(n527), .B(n84), .Z(\ab[23][60] ) );
  NR2 U3342 ( .A(n528), .B(n85), .Z(\ab[23][59] ) );
  NR2 U3343 ( .A(n529), .B(n85), .Z(\ab[23][58] ) );
  NR2 U3344 ( .A(n530), .B(n85), .Z(\ab[23][57] ) );
  NR2 U3345 ( .A(n531), .B(n85), .Z(\ab[23][56] ) );
  NR2 U3346 ( .A(n532), .B(n85), .Z(\ab[23][55] ) );
  NR2 U3347 ( .A(n533), .B(n85), .Z(\ab[23][54] ) );
  NR2 U3348 ( .A(n534), .B(n85), .Z(\ab[23][53] ) );
  NR2 U3349 ( .A(n535), .B(n85), .Z(\ab[23][52] ) );
  NR2 U3350 ( .A(n536), .B(n85), .Z(\ab[23][51] ) );
  NR2 U3351 ( .A(n537), .B(n85), .Z(\ab[23][50] ) );
  NR2 U3352 ( .A(n538), .B(n85), .Z(\ab[23][49] ) );
  NR2 U3353 ( .A(n539), .B(n85), .Z(\ab[23][48] ) );
  NR2 U3354 ( .A(n540), .B(n86), .Z(\ab[23][47] ) );
  NR2 U3355 ( .A(n541), .B(n86), .Z(\ab[23][46] ) );
  NR2 U3356 ( .A(n542), .B(n86), .Z(\ab[23][45] ) );
  NR2 U3357 ( .A(n543), .B(n86), .Z(\ab[23][44] ) );
  NR2 U3358 ( .A(n544), .B(n86), .Z(\ab[23][43] ) );
  NR2 U3359 ( .A(n545), .B(n86), .Z(\ab[23][42] ) );
  NR2 U3360 ( .A(n546), .B(n86), .Z(\ab[23][41] ) );
  NR2 U3361 ( .A(n547), .B(n86), .Z(\ab[23][40] ) );
  NR2 U3362 ( .A(n548), .B(n86), .Z(\ab[23][39] ) );
  NR2 U3363 ( .A(n492), .B(n4), .Z(\ab[22][95] ) );
  NR2 U3364 ( .A(n493), .B(n4), .Z(\ab[22][94] ) );
  NR2 U3365 ( .A(n494), .B(n4), .Z(\ab[22][93] ) );
  NR2 U3366 ( .A(n495), .B(n4), .Z(\ab[22][92] ) );
  NR2 U3367 ( .A(n496), .B(n4), .Z(\ab[22][91] ) );
  NR2 U3368 ( .A(n497), .B(n4), .Z(\ab[22][90] ) );
  NR2 U3369 ( .A(n498), .B(n4), .Z(\ab[22][89] ) );
  NR2 U3370 ( .A(n499), .B(n4), .Z(\ab[22][88] ) );
  NR2 U3371 ( .A(n500), .B(n4), .Z(\ab[22][87] ) );
  NR2 U3372 ( .A(n501), .B(n4), .Z(\ab[22][86] ) );
  NR2 U3373 ( .A(n502), .B(n4), .Z(\ab[22][85] ) );
  NR2 U3374 ( .A(n503), .B(n4), .Z(\ab[22][84] ) );
  NR2 U3375 ( .A(n504), .B(n557), .Z(\ab[22][83] ) );
  NR2 U3376 ( .A(n505), .B(n4), .Z(\ab[22][82] ) );
  NR2 U3377 ( .A(n506), .B(n557), .Z(\ab[22][81] ) );
  NR2 U3378 ( .A(n507), .B(n4), .Z(\ab[22][80] ) );
  NR2 U3379 ( .A(n508), .B(n4), .Z(\ab[22][79] ) );
  NR2 U3380 ( .A(n509), .B(n4), .Z(\ab[22][78] ) );
  NR2 U3381 ( .A(n510), .B(n4), .Z(\ab[22][77] ) );
  NR2 U3382 ( .A(n511), .B(n4), .Z(\ab[22][76] ) );
  NR2 U3383 ( .A(n512), .B(n4), .Z(\ab[22][75] ) );
  NR2 U3384 ( .A(n513), .B(n4), .Z(\ab[22][74] ) );
  NR2 U3385 ( .A(n514), .B(n4), .Z(\ab[22][73] ) );
  NR2 U3386 ( .A(n515), .B(n4), .Z(\ab[22][72] ) );
  NR2 U3387 ( .A(n516), .B(n557), .Z(\ab[22][71] ) );
  NR2 U3388 ( .A(n517), .B(n557), .Z(\ab[22][70] ) );
  NR2 U3389 ( .A(n518), .B(n557), .Z(\ab[22][69] ) );
  NR2 U3390 ( .A(n519), .B(n4), .Z(\ab[22][68] ) );
  NR2 U3391 ( .A(n520), .B(n557), .Z(\ab[22][67] ) );
  NR2 U3392 ( .A(n521), .B(n557), .Z(\ab[22][66] ) );
  NR2 U3393 ( .A(n522), .B(n557), .Z(\ab[22][65] ) );
  NR2 U3394 ( .A(n523), .B(n4), .Z(\ab[22][64] ) );
  NR2 U3395 ( .A(n524), .B(n557), .Z(\ab[22][63] ) );
  NR2 U3396 ( .A(n525), .B(n557), .Z(\ab[22][62] ) );
  NR2 U3397 ( .A(n526), .B(n557), .Z(\ab[22][61] ) );
  NR2 U3398 ( .A(n527), .B(n4), .Z(\ab[22][60] ) );
  NR2 U3399 ( .A(n528), .B(n557), .Z(\ab[22][59] ) );
  NR2 U3400 ( .A(n529), .B(n557), .Z(\ab[22][58] ) );
  NR2 U3401 ( .A(n530), .B(n557), .Z(\ab[22][57] ) );
  NR2 U3402 ( .A(n531), .B(n557), .Z(\ab[22][56] ) );
  NR2 U3403 ( .A(n532), .B(n557), .Z(\ab[22][55] ) );
  NR2 U3404 ( .A(n533), .B(n557), .Z(\ab[22][54] ) );
  NR2 U3405 ( .A(n534), .B(n557), .Z(\ab[22][53] ) );
  NR2 U3406 ( .A(n535), .B(n557), .Z(\ab[22][52] ) );
  NR2 U3407 ( .A(n536), .B(n557), .Z(\ab[22][51] ) );
  NR2 U3408 ( .A(n537), .B(n557), .Z(\ab[22][50] ) );
  NR2 U3409 ( .A(n538), .B(n557), .Z(\ab[22][49] ) );
  NR2 U3410 ( .A(n539), .B(n557), .Z(\ab[22][48] ) );
  NR2 U3411 ( .A(n540), .B(n557), .Z(\ab[22][47] ) );
  NR2 U3412 ( .A(n541), .B(n557), .Z(\ab[22][46] ) );
  NR2 U3413 ( .A(n542), .B(n557), .Z(\ab[22][45] ) );
  NR2 U3414 ( .A(n543), .B(n557), .Z(\ab[22][44] ) );
  NR2 U3415 ( .A(n544), .B(n557), .Z(\ab[22][43] ) );
  NR2 U3416 ( .A(n545), .B(n557), .Z(\ab[22][42] ) );
  NR2 U3417 ( .A(n546), .B(n557), .Z(\ab[22][41] ) );
  NR2 U3418 ( .A(n547), .B(n557), .Z(\ab[22][40] ) );
  NR2 U3419 ( .A(n548), .B(n557), .Z(\ab[22][39] ) );
  NR2 U3420 ( .A(n492), .B(n98), .Z(\ab[21][95] ) );
  NR2 U3421 ( .A(n493), .B(n98), .Z(\ab[21][94] ) );
  NR2 U3422 ( .A(n494), .B(n98), .Z(\ab[21][93] ) );
  NR2 U3423 ( .A(n495), .B(n98), .Z(\ab[21][92] ) );
  NR2 U3424 ( .A(n496), .B(n98), .Z(\ab[21][91] ) );
  NR2 U3425 ( .A(n497), .B(n98), .Z(\ab[21][90] ) );
  NR2 U3426 ( .A(n498), .B(n98), .Z(\ab[21][89] ) );
  NR2 U3427 ( .A(n499), .B(n98), .Z(\ab[21][88] ) );
  NR2 U3428 ( .A(n500), .B(n98), .Z(\ab[21][87] ) );
  NR2 U3429 ( .A(n501), .B(n98), .Z(\ab[21][86] ) );
  NR2 U3430 ( .A(n502), .B(n98), .Z(\ab[21][85] ) );
  NR2 U3431 ( .A(n503), .B(n98), .Z(\ab[21][84] ) );
  NR2 U3432 ( .A(n504), .B(n99), .Z(\ab[21][83] ) );
  NR2 U3433 ( .A(n505), .B(n99), .Z(\ab[21][82] ) );
  NR2 U3434 ( .A(n506), .B(n99), .Z(\ab[21][81] ) );
  NR2 U3435 ( .A(n507), .B(n99), .Z(\ab[21][80] ) );
  NR2 U3436 ( .A(n508), .B(n99), .Z(\ab[21][79] ) );
  NR2 U3437 ( .A(n509), .B(n99), .Z(\ab[21][78] ) );
  NR2 U3438 ( .A(n510), .B(n99), .Z(\ab[21][77] ) );
  NR2 U3439 ( .A(n511), .B(n99), .Z(\ab[21][76] ) );
  NR2 U3440 ( .A(n512), .B(n99), .Z(\ab[21][75] ) );
  NR2 U3441 ( .A(n513), .B(n99), .Z(\ab[21][74] ) );
  NR2 U3442 ( .A(n514), .B(n99), .Z(\ab[21][73] ) );
  NR2 U3443 ( .A(n515), .B(n99), .Z(\ab[21][72] ) );
  NR2 U3444 ( .A(n516), .B(n100), .Z(\ab[21][71] ) );
  NR2 U3445 ( .A(n517), .B(n100), .Z(\ab[21][70] ) );
  NR2 U3446 ( .A(n518), .B(n100), .Z(\ab[21][69] ) );
  NR2 U3447 ( .A(n519), .B(n100), .Z(\ab[21][68] ) );
  NR2 U3448 ( .A(n520), .B(n100), .Z(\ab[21][67] ) );
  NR2 U3449 ( .A(n521), .B(n100), .Z(\ab[21][66] ) );
  NR2 U3450 ( .A(n522), .B(n100), .Z(\ab[21][65] ) );
  NR2 U3451 ( .A(n523), .B(n100), .Z(\ab[21][64] ) );
  NR2 U3452 ( .A(n524), .B(n100), .Z(\ab[21][63] ) );
  NR2 U3453 ( .A(n525), .B(n100), .Z(\ab[21][62] ) );
  NR2 U3454 ( .A(n526), .B(n100), .Z(\ab[21][61] ) );
  NR2 U3455 ( .A(n527), .B(n100), .Z(\ab[21][60] ) );
  NR2 U3456 ( .A(n528), .B(n101), .Z(\ab[21][59] ) );
  NR2 U3457 ( .A(n529), .B(n101), .Z(\ab[21][58] ) );
  NR2 U3458 ( .A(n530), .B(n101), .Z(\ab[21][57] ) );
  NR2 U3459 ( .A(n531), .B(n101), .Z(\ab[21][56] ) );
  NR2 U3460 ( .A(n532), .B(n101), .Z(\ab[21][55] ) );
  NR2 U3461 ( .A(n533), .B(n101), .Z(\ab[21][54] ) );
  NR2 U3462 ( .A(n534), .B(n101), .Z(\ab[21][53] ) );
  NR2 U3463 ( .A(n535), .B(n101), .Z(\ab[21][52] ) );
  NR2 U3464 ( .A(n536), .B(n101), .Z(\ab[21][51] ) );
  NR2 U3465 ( .A(n537), .B(n101), .Z(\ab[21][50] ) );
  NR2 U3466 ( .A(n538), .B(n101), .Z(\ab[21][49] ) );
  NR2 U3467 ( .A(n539), .B(n101), .Z(\ab[21][48] ) );
  NR2 U3468 ( .A(n540), .B(n102), .Z(\ab[21][47] ) );
  NR2 U3469 ( .A(n541), .B(n102), .Z(\ab[21][46] ) );
  NR2 U3470 ( .A(n542), .B(n102), .Z(\ab[21][45] ) );
  NR2 U3471 ( .A(n543), .B(n102), .Z(\ab[21][44] ) );
  NR2 U3472 ( .A(n544), .B(n102), .Z(\ab[21][43] ) );
  NR2 U3473 ( .A(n545), .B(n102), .Z(\ab[21][42] ) );
  NR2 U3474 ( .A(n546), .B(n102), .Z(\ab[21][41] ) );
  NR2 U3475 ( .A(n547), .B(n102), .Z(\ab[21][40] ) );
  NR2 U3476 ( .A(n548), .B(n102), .Z(\ab[21][39] ) );
  NR2 U3477 ( .A(n492), .B(n109), .Z(\ab[20][95] ) );
  NR2 U3478 ( .A(n493), .B(n109), .Z(\ab[20][94] ) );
  NR2 U3479 ( .A(n494), .B(n109), .Z(\ab[20][93] ) );
  NR2 U3480 ( .A(n495), .B(n109), .Z(\ab[20][92] ) );
  NR2 U3481 ( .A(n496), .B(n109), .Z(\ab[20][91] ) );
  NR2 U3482 ( .A(n497), .B(n109), .Z(\ab[20][90] ) );
  NR2 U3483 ( .A(n498), .B(n109), .Z(\ab[20][89] ) );
  NR2 U3484 ( .A(n499), .B(n109), .Z(\ab[20][88] ) );
  NR2 U3485 ( .A(n500), .B(n109), .Z(\ab[20][87] ) );
  NR2 U3486 ( .A(n501), .B(n109), .Z(\ab[20][86] ) );
  NR2 U3487 ( .A(n502), .B(n109), .Z(\ab[20][85] ) );
  NR2 U3488 ( .A(n503), .B(n109), .Z(\ab[20][84] ) );
  NR2 U3489 ( .A(n504), .B(n110), .Z(\ab[20][83] ) );
  NR2 U3490 ( .A(n505), .B(n110), .Z(\ab[20][82] ) );
  NR2 U3491 ( .A(n506), .B(n110), .Z(\ab[20][81] ) );
  NR2 U3492 ( .A(n507), .B(n110), .Z(\ab[20][80] ) );
  NR2 U3493 ( .A(n508), .B(n110), .Z(\ab[20][79] ) );
  NR2 U3494 ( .A(n509), .B(n110), .Z(\ab[20][78] ) );
  NR2 U3495 ( .A(n510), .B(n110), .Z(\ab[20][77] ) );
  NR2 U3496 ( .A(n511), .B(n110), .Z(\ab[20][76] ) );
  NR2 U3497 ( .A(n512), .B(n110), .Z(\ab[20][75] ) );
  NR2 U3498 ( .A(n513), .B(n110), .Z(\ab[20][74] ) );
  NR2 U3499 ( .A(n514), .B(n110), .Z(\ab[20][73] ) );
  NR2 U3500 ( .A(n515), .B(n110), .Z(\ab[20][72] ) );
  NR2 U3501 ( .A(n516), .B(n111), .Z(\ab[20][71] ) );
  NR2 U3502 ( .A(n517), .B(n111), .Z(\ab[20][70] ) );
  NR2 U3503 ( .A(n518), .B(n111), .Z(\ab[20][69] ) );
  NR2 U3504 ( .A(n519), .B(n111), .Z(\ab[20][68] ) );
  NR2 U3505 ( .A(n520), .B(n111), .Z(\ab[20][67] ) );
  NR2 U3506 ( .A(n521), .B(n111), .Z(\ab[20][66] ) );
  NR2 U3507 ( .A(n522), .B(n111), .Z(\ab[20][65] ) );
  NR2 U3508 ( .A(n523), .B(n111), .Z(\ab[20][64] ) );
  NR2 U3509 ( .A(n524), .B(n111), .Z(\ab[20][63] ) );
  NR2 U3510 ( .A(n525), .B(n111), .Z(\ab[20][62] ) );
  NR2 U3511 ( .A(n526), .B(n111), .Z(\ab[20][61] ) );
  NR2 U3512 ( .A(n527), .B(n111), .Z(\ab[20][60] ) );
  NR2 U3513 ( .A(n528), .B(n112), .Z(\ab[20][59] ) );
  NR2 U3514 ( .A(n529), .B(n112), .Z(\ab[20][58] ) );
  NR2 U3515 ( .A(n530), .B(n112), .Z(\ab[20][57] ) );
  NR2 U3516 ( .A(n531), .B(n112), .Z(\ab[20][56] ) );
  NR2 U3517 ( .A(n532), .B(n112), .Z(\ab[20][55] ) );
  NR2 U3518 ( .A(n533), .B(n112), .Z(\ab[20][54] ) );
  NR2 U3519 ( .A(n534), .B(n112), .Z(\ab[20][53] ) );
  NR2 U3520 ( .A(n535), .B(n112), .Z(\ab[20][52] ) );
  NR2 U3521 ( .A(n536), .B(n112), .Z(\ab[20][51] ) );
  NR2 U3522 ( .A(n537), .B(n112), .Z(\ab[20][50] ) );
  NR2 U3523 ( .A(n538), .B(n112), .Z(\ab[20][49] ) );
  NR2 U3524 ( .A(n539), .B(n112), .Z(\ab[20][48] ) );
  NR2 U3525 ( .A(n540), .B(n113), .Z(\ab[20][47] ) );
  NR2 U3526 ( .A(n541), .B(n113), .Z(\ab[20][46] ) );
  NR2 U3527 ( .A(n542), .B(n113), .Z(\ab[20][45] ) );
  NR2 U3528 ( .A(n543), .B(n113), .Z(\ab[20][44] ) );
  NR2 U3529 ( .A(n544), .B(n113), .Z(\ab[20][43] ) );
  NR2 U3530 ( .A(n545), .B(n113), .Z(\ab[20][42] ) );
  NR2 U3531 ( .A(n546), .B(n113), .Z(\ab[20][41] ) );
  NR2 U3532 ( .A(n547), .B(n113), .Z(\ab[20][40] ) );
  NR2 U3533 ( .A(n548), .B(n113), .Z(\ab[20][39] ) );
  NR2 U3534 ( .A(n492), .B(n120), .Z(\ab[19][95] ) );
  NR2 U3535 ( .A(n493), .B(n120), .Z(\ab[19][94] ) );
  NR2 U3536 ( .A(n494), .B(n120), .Z(\ab[19][93] ) );
  NR2 U3537 ( .A(n495), .B(n120), .Z(\ab[19][92] ) );
  NR2 U3538 ( .A(n496), .B(n120), .Z(\ab[19][91] ) );
  NR2 U3539 ( .A(n497), .B(n120), .Z(\ab[19][90] ) );
  NR2 U3540 ( .A(n498), .B(n120), .Z(\ab[19][89] ) );
  NR2 U3541 ( .A(n499), .B(n120), .Z(\ab[19][88] ) );
  NR2 U3542 ( .A(n500), .B(n120), .Z(\ab[19][87] ) );
  NR2 U3543 ( .A(n501), .B(n120), .Z(\ab[19][86] ) );
  NR2 U3544 ( .A(n502), .B(n120), .Z(\ab[19][85] ) );
  NR2 U3545 ( .A(n503), .B(n120), .Z(\ab[19][84] ) );
  NR2 U3546 ( .A(n504), .B(n121), .Z(\ab[19][83] ) );
  NR2 U3547 ( .A(n505), .B(n121), .Z(\ab[19][82] ) );
  NR2 U3548 ( .A(n506), .B(n121), .Z(\ab[19][81] ) );
  NR2 U3549 ( .A(n507), .B(n121), .Z(\ab[19][80] ) );
  NR2 U3550 ( .A(n508), .B(n121), .Z(\ab[19][79] ) );
  NR2 U3551 ( .A(n509), .B(n121), .Z(\ab[19][78] ) );
  NR2 U3552 ( .A(n510), .B(n121), .Z(\ab[19][77] ) );
  NR2 U3553 ( .A(n511), .B(n121), .Z(\ab[19][76] ) );
  NR2 U3554 ( .A(n512), .B(n121), .Z(\ab[19][75] ) );
  NR2 U3555 ( .A(n513), .B(n121), .Z(\ab[19][74] ) );
  NR2 U3556 ( .A(n514), .B(n121), .Z(\ab[19][73] ) );
  NR2 U3557 ( .A(n515), .B(n121), .Z(\ab[19][72] ) );
  NR2 U3558 ( .A(n516), .B(n122), .Z(\ab[19][71] ) );
  NR2 U3559 ( .A(n517), .B(n122), .Z(\ab[19][70] ) );
  NR2 U3560 ( .A(n518), .B(n122), .Z(\ab[19][69] ) );
  NR2 U3561 ( .A(n519), .B(n122), .Z(\ab[19][68] ) );
  NR2 U3562 ( .A(n520), .B(n122), .Z(\ab[19][67] ) );
  NR2 U3563 ( .A(n521), .B(n122), .Z(\ab[19][66] ) );
  NR2 U3564 ( .A(n522), .B(n122), .Z(\ab[19][65] ) );
  NR2 U3565 ( .A(n523), .B(n122), .Z(\ab[19][64] ) );
  NR2 U3566 ( .A(n524), .B(n122), .Z(\ab[19][63] ) );
  NR2 U3567 ( .A(n525), .B(n122), .Z(\ab[19][62] ) );
  NR2 U3568 ( .A(n526), .B(n122), .Z(\ab[19][61] ) );
  NR2 U3569 ( .A(n527), .B(n122), .Z(\ab[19][60] ) );
  NR2 U3570 ( .A(n528), .B(n123), .Z(\ab[19][59] ) );
  NR2 U3571 ( .A(n529), .B(n123), .Z(\ab[19][58] ) );
  NR2 U3572 ( .A(n530), .B(n123), .Z(\ab[19][57] ) );
  NR2 U3573 ( .A(n531), .B(n123), .Z(\ab[19][56] ) );
  NR2 U3574 ( .A(n532), .B(n123), .Z(\ab[19][55] ) );
  NR2 U3575 ( .A(n533), .B(n123), .Z(\ab[19][54] ) );
  NR2 U3576 ( .A(n534), .B(n123), .Z(\ab[19][53] ) );
  NR2 U3577 ( .A(n535), .B(n123), .Z(\ab[19][52] ) );
  NR2 U3578 ( .A(n536), .B(n123), .Z(\ab[19][51] ) );
  NR2 U3579 ( .A(n537), .B(n123), .Z(\ab[19][50] ) );
  NR2 U3580 ( .A(n538), .B(n123), .Z(\ab[19][49] ) );
  NR2 U3581 ( .A(n539), .B(n123), .Z(\ab[19][48] ) );
  NR2 U3582 ( .A(n540), .B(n124), .Z(\ab[19][47] ) );
  NR2 U3583 ( .A(n541), .B(n124), .Z(\ab[19][46] ) );
  NR2 U3584 ( .A(n542), .B(n124), .Z(\ab[19][45] ) );
  NR2 U3585 ( .A(n543), .B(n124), .Z(\ab[19][44] ) );
  NR2 U3586 ( .A(n544), .B(n124), .Z(\ab[19][43] ) );
  NR2 U3587 ( .A(n545), .B(n124), .Z(\ab[19][42] ) );
  NR2 U3588 ( .A(n546), .B(n124), .Z(\ab[19][41] ) );
  NR2 U3589 ( .A(n547), .B(n124), .Z(\ab[19][40] ) );
  NR2 U3590 ( .A(n548), .B(n124), .Z(\ab[19][39] ) );
  NR2 U3591 ( .A(n492), .B(n131), .Z(\ab[18][95] ) );
  NR2 U3592 ( .A(n493), .B(n131), .Z(\ab[18][94] ) );
  NR2 U3593 ( .A(n494), .B(n131), .Z(\ab[18][93] ) );
  NR2 U3594 ( .A(n495), .B(n131), .Z(\ab[18][92] ) );
  NR2 U3595 ( .A(n496), .B(n131), .Z(\ab[18][91] ) );
  NR2 U3596 ( .A(n497), .B(n131), .Z(\ab[18][90] ) );
  NR2 U3597 ( .A(n498), .B(n131), .Z(\ab[18][89] ) );
  NR2 U3598 ( .A(n499), .B(n131), .Z(\ab[18][88] ) );
  NR2 U3599 ( .A(n500), .B(n131), .Z(\ab[18][87] ) );
  NR2 U3600 ( .A(n501), .B(n131), .Z(\ab[18][86] ) );
  NR2 U3601 ( .A(n502), .B(n131), .Z(\ab[18][85] ) );
  NR2 U3602 ( .A(n503), .B(n131), .Z(\ab[18][84] ) );
  NR2 U3603 ( .A(n504), .B(n132), .Z(\ab[18][83] ) );
  NR2 U3604 ( .A(n505), .B(n132), .Z(\ab[18][82] ) );
  NR2 U3605 ( .A(n506), .B(n132), .Z(\ab[18][81] ) );
  NR2 U3606 ( .A(n507), .B(n132), .Z(\ab[18][80] ) );
  NR2 U3607 ( .A(n508), .B(n132), .Z(\ab[18][79] ) );
  NR2 U3608 ( .A(n509), .B(n132), .Z(\ab[18][78] ) );
  NR2 U3609 ( .A(n510), .B(n132), .Z(\ab[18][77] ) );
  NR2 U3610 ( .A(n511), .B(n132), .Z(\ab[18][76] ) );
  NR2 U3611 ( .A(n512), .B(n132), .Z(\ab[18][75] ) );
  NR2 U3612 ( .A(n513), .B(n132), .Z(\ab[18][74] ) );
  NR2 U3613 ( .A(n514), .B(n132), .Z(\ab[18][73] ) );
  NR2 U3614 ( .A(n515), .B(n132), .Z(\ab[18][72] ) );
  NR2 U3615 ( .A(n516), .B(n133), .Z(\ab[18][71] ) );
  NR2 U3616 ( .A(n517), .B(n133), .Z(\ab[18][70] ) );
  NR2 U3617 ( .A(n518), .B(n133), .Z(\ab[18][69] ) );
  NR2 U3618 ( .A(n519), .B(n133), .Z(\ab[18][68] ) );
  NR2 U3619 ( .A(n520), .B(n133), .Z(\ab[18][67] ) );
  NR2 U3620 ( .A(n521), .B(n133), .Z(\ab[18][66] ) );
  NR2 U3621 ( .A(n522), .B(n133), .Z(\ab[18][65] ) );
  NR2 U3622 ( .A(n523), .B(n133), .Z(\ab[18][64] ) );
  NR2 U3623 ( .A(n524), .B(n133), .Z(\ab[18][63] ) );
  NR2 U3624 ( .A(n525), .B(n133), .Z(\ab[18][62] ) );
  NR2 U3625 ( .A(n526), .B(n133), .Z(\ab[18][61] ) );
  NR2 U3626 ( .A(n527), .B(n133), .Z(\ab[18][60] ) );
  NR2 U3627 ( .A(n528), .B(n134), .Z(\ab[18][59] ) );
  NR2 U3628 ( .A(n529), .B(n134), .Z(\ab[18][58] ) );
  NR2 U3629 ( .A(n530), .B(n134), .Z(\ab[18][57] ) );
  NR2 U3630 ( .A(n531), .B(n134), .Z(\ab[18][56] ) );
  NR2 U3631 ( .A(n532), .B(n134), .Z(\ab[18][55] ) );
  NR2 U3632 ( .A(n533), .B(n134), .Z(\ab[18][54] ) );
  NR2 U3633 ( .A(n534), .B(n134), .Z(\ab[18][53] ) );
  NR2 U3634 ( .A(n535), .B(n134), .Z(\ab[18][52] ) );
  NR2 U3635 ( .A(n536), .B(n134), .Z(\ab[18][51] ) );
  NR2 U3636 ( .A(n537), .B(n134), .Z(\ab[18][50] ) );
  NR2 U3637 ( .A(n538), .B(n134), .Z(\ab[18][49] ) );
  NR2 U3638 ( .A(n539), .B(n134), .Z(\ab[18][48] ) );
  NR2 U3639 ( .A(n540), .B(n135), .Z(\ab[18][47] ) );
  NR2 U3640 ( .A(n541), .B(n135), .Z(\ab[18][46] ) );
  NR2 U3641 ( .A(n542), .B(n135), .Z(\ab[18][45] ) );
  NR2 U3642 ( .A(n543), .B(n135), .Z(\ab[18][44] ) );
  NR2 U3643 ( .A(n544), .B(n135), .Z(\ab[18][43] ) );
  NR2 U3644 ( .A(n545), .B(n135), .Z(\ab[18][42] ) );
  NR2 U3645 ( .A(n546), .B(n135), .Z(\ab[18][41] ) );
  NR2 U3646 ( .A(n547), .B(n135), .Z(\ab[18][40] ) );
  NR2 U3647 ( .A(n548), .B(n135), .Z(\ab[18][39] ) );
  NR2 U3648 ( .A(n492), .B(n142), .Z(\ab[17][95] ) );
  NR2 U3649 ( .A(n493), .B(n142), .Z(\ab[17][94] ) );
  NR2 U3650 ( .A(n494), .B(n142), .Z(\ab[17][93] ) );
  NR2 U3651 ( .A(n495), .B(n142), .Z(\ab[17][92] ) );
  NR2 U3652 ( .A(n496), .B(n142), .Z(\ab[17][91] ) );
  NR2 U3653 ( .A(n497), .B(n142), .Z(\ab[17][90] ) );
  NR2 U3654 ( .A(n498), .B(n142), .Z(\ab[17][89] ) );
  NR2 U3655 ( .A(n499), .B(n142), .Z(\ab[17][88] ) );
  NR2 U3656 ( .A(n500), .B(n142), .Z(\ab[17][87] ) );
  NR2 U3657 ( .A(n501), .B(n142), .Z(\ab[17][86] ) );
  NR2 U3658 ( .A(n502), .B(n142), .Z(\ab[17][85] ) );
  NR2 U3659 ( .A(n503), .B(n142), .Z(\ab[17][84] ) );
  NR2 U3660 ( .A(n504), .B(n143), .Z(\ab[17][83] ) );
  NR2 U3661 ( .A(n505), .B(n143), .Z(\ab[17][82] ) );
  NR2 U3662 ( .A(n506), .B(n143), .Z(\ab[17][81] ) );
  NR2 U3663 ( .A(n507), .B(n143), .Z(\ab[17][80] ) );
  NR2 U3664 ( .A(n508), .B(n143), .Z(\ab[17][79] ) );
  NR2 U3665 ( .A(n509), .B(n143), .Z(\ab[17][78] ) );
  NR2 U3666 ( .A(n510), .B(n143), .Z(\ab[17][77] ) );
  NR2 U3667 ( .A(n511), .B(n143), .Z(\ab[17][76] ) );
  NR2 U3668 ( .A(n512), .B(n143), .Z(\ab[17][75] ) );
  NR2 U3669 ( .A(n513), .B(n143), .Z(\ab[17][74] ) );
  NR2 U3670 ( .A(n514), .B(n143), .Z(\ab[17][73] ) );
  NR2 U3671 ( .A(n515), .B(n143), .Z(\ab[17][72] ) );
  NR2 U3672 ( .A(n516), .B(n144), .Z(\ab[17][71] ) );
  NR2 U3673 ( .A(n517), .B(n144), .Z(\ab[17][70] ) );
  NR2 U3674 ( .A(n518), .B(n144), .Z(\ab[17][69] ) );
  NR2 U3675 ( .A(n519), .B(n144), .Z(\ab[17][68] ) );
  NR2 U3676 ( .A(n520), .B(n144), .Z(\ab[17][67] ) );
  NR2 U3677 ( .A(n521), .B(n144), .Z(\ab[17][66] ) );
  NR2 U3678 ( .A(n522), .B(n144), .Z(\ab[17][65] ) );
  NR2 U3679 ( .A(n523), .B(n144), .Z(\ab[17][64] ) );
  NR2 U3680 ( .A(n524), .B(n144), .Z(\ab[17][63] ) );
  NR2 U3681 ( .A(n525), .B(n144), .Z(\ab[17][62] ) );
  NR2 U3682 ( .A(n526), .B(n144), .Z(\ab[17][61] ) );
  NR2 U3683 ( .A(n527), .B(n144), .Z(\ab[17][60] ) );
  NR2 U3684 ( .A(n528), .B(n145), .Z(\ab[17][59] ) );
  NR2 U3685 ( .A(n529), .B(n145), .Z(\ab[17][58] ) );
  NR2 U3686 ( .A(n530), .B(n145), .Z(\ab[17][57] ) );
  NR2 U3687 ( .A(n531), .B(n145), .Z(\ab[17][56] ) );
  NR2 U3688 ( .A(n532), .B(n145), .Z(\ab[17][55] ) );
  NR2 U3689 ( .A(n533), .B(n145), .Z(\ab[17][54] ) );
  NR2 U3690 ( .A(n534), .B(n145), .Z(\ab[17][53] ) );
  NR2 U3691 ( .A(n535), .B(n145), .Z(\ab[17][52] ) );
  NR2 U3692 ( .A(n536), .B(n145), .Z(\ab[17][51] ) );
  NR2 U3693 ( .A(n537), .B(n145), .Z(\ab[17][50] ) );
  NR2 U3694 ( .A(n538), .B(n145), .Z(\ab[17][49] ) );
  NR2 U3695 ( .A(n539), .B(n145), .Z(\ab[17][48] ) );
  NR2 U3696 ( .A(n540), .B(n146), .Z(\ab[17][47] ) );
  NR2 U3697 ( .A(n541), .B(n146), .Z(\ab[17][46] ) );
  NR2 U3698 ( .A(n542), .B(n146), .Z(\ab[17][45] ) );
  NR2 U3699 ( .A(n543), .B(n146), .Z(\ab[17][44] ) );
  NR2 U3700 ( .A(n544), .B(n146), .Z(\ab[17][43] ) );
  NR2 U3701 ( .A(n545), .B(n146), .Z(\ab[17][42] ) );
  NR2 U3702 ( .A(n546), .B(n146), .Z(\ab[17][41] ) );
  NR2 U3703 ( .A(n547), .B(n146), .Z(\ab[17][40] ) );
  NR2 U3704 ( .A(n548), .B(n146), .Z(\ab[17][39] ) );
  NR2 U3705 ( .A(n492), .B(n153), .Z(\ab[16][95] ) );
  NR2 U3706 ( .A(n493), .B(n153), .Z(\ab[16][94] ) );
  NR2 U3707 ( .A(n494), .B(n153), .Z(\ab[16][93] ) );
  NR2 U3708 ( .A(n495), .B(n153), .Z(\ab[16][92] ) );
  NR2 U3709 ( .A(n496), .B(n153), .Z(\ab[16][91] ) );
  NR2 U3710 ( .A(n497), .B(n153), .Z(\ab[16][90] ) );
  NR2 U3711 ( .A(n498), .B(n153), .Z(\ab[16][89] ) );
  NR2 U3712 ( .A(n499), .B(n153), .Z(\ab[16][88] ) );
  NR2 U3713 ( .A(n500), .B(n153), .Z(\ab[16][87] ) );
  NR2 U3714 ( .A(n501), .B(n153), .Z(\ab[16][86] ) );
  NR2 U3715 ( .A(n502), .B(n153), .Z(\ab[16][85] ) );
  NR2 U3716 ( .A(n503), .B(n153), .Z(\ab[16][84] ) );
  NR2 U3717 ( .A(n504), .B(n154), .Z(\ab[16][83] ) );
  NR2 U3718 ( .A(n505), .B(n154), .Z(\ab[16][82] ) );
  NR2 U3719 ( .A(n506), .B(n154), .Z(\ab[16][81] ) );
  NR2 U3720 ( .A(n507), .B(n154), .Z(\ab[16][80] ) );
  NR2 U3721 ( .A(n508), .B(n154), .Z(\ab[16][79] ) );
  NR2 U3722 ( .A(n509), .B(n154), .Z(\ab[16][78] ) );
  NR2 U3723 ( .A(n510), .B(n154), .Z(\ab[16][77] ) );
  NR2 U3724 ( .A(n511), .B(n154), .Z(\ab[16][76] ) );
  NR2 U3725 ( .A(n512), .B(n154), .Z(\ab[16][75] ) );
  NR2 U3726 ( .A(n513), .B(n154), .Z(\ab[16][74] ) );
  NR2 U3727 ( .A(n514), .B(n154), .Z(\ab[16][73] ) );
  NR2 U3728 ( .A(n515), .B(n154), .Z(\ab[16][72] ) );
  NR2 U3729 ( .A(n516), .B(n155), .Z(\ab[16][71] ) );
  NR2 U3730 ( .A(n517), .B(n155), .Z(\ab[16][70] ) );
  NR2 U3731 ( .A(n518), .B(n155), .Z(\ab[16][69] ) );
  NR2 U3732 ( .A(n519), .B(n155), .Z(\ab[16][68] ) );
  NR2 U3733 ( .A(n520), .B(n155), .Z(\ab[16][67] ) );
  NR2 U3734 ( .A(n521), .B(n155), .Z(\ab[16][66] ) );
  NR2 U3735 ( .A(n522), .B(n155), .Z(\ab[16][65] ) );
  NR2 U3736 ( .A(n523), .B(n155), .Z(\ab[16][64] ) );
  NR2 U3737 ( .A(n524), .B(n155), .Z(\ab[16][63] ) );
  NR2 U3738 ( .A(n525), .B(n155), .Z(\ab[16][62] ) );
  NR2 U3739 ( .A(n526), .B(n155), .Z(\ab[16][61] ) );
  NR2 U3740 ( .A(n527), .B(n155), .Z(\ab[16][60] ) );
  NR2 U3741 ( .A(n528), .B(n156), .Z(\ab[16][59] ) );
  NR2 U3742 ( .A(n529), .B(n156), .Z(\ab[16][58] ) );
  NR2 U3743 ( .A(n530), .B(n156), .Z(\ab[16][57] ) );
  NR2 U3744 ( .A(n531), .B(n156), .Z(\ab[16][56] ) );
  NR2 U3745 ( .A(n532), .B(n156), .Z(\ab[16][55] ) );
  NR2 U3746 ( .A(n533), .B(n156), .Z(\ab[16][54] ) );
  NR2 U3747 ( .A(n534), .B(n156), .Z(\ab[16][53] ) );
  NR2 U3748 ( .A(n535), .B(n156), .Z(\ab[16][52] ) );
  NR2 U3749 ( .A(n536), .B(n156), .Z(\ab[16][51] ) );
  NR2 U3750 ( .A(n537), .B(n156), .Z(\ab[16][50] ) );
  NR2 U3751 ( .A(n538), .B(n156), .Z(\ab[16][49] ) );
  NR2 U3752 ( .A(n539), .B(n156), .Z(\ab[16][48] ) );
  NR2 U3753 ( .A(n540), .B(n157), .Z(\ab[16][47] ) );
  NR2 U3754 ( .A(n541), .B(n157), .Z(\ab[16][46] ) );
  NR2 U3755 ( .A(n542), .B(n157), .Z(\ab[16][45] ) );
  NR2 U3756 ( .A(n543), .B(n157), .Z(\ab[16][44] ) );
  NR2 U3757 ( .A(n544), .B(n157), .Z(\ab[16][43] ) );
  NR2 U3758 ( .A(n545), .B(n157), .Z(\ab[16][42] ) );
  NR2 U3759 ( .A(n546), .B(n157), .Z(\ab[16][41] ) );
  NR2 U3760 ( .A(n547), .B(n157), .Z(\ab[16][40] ) );
  NR2 U3761 ( .A(n548), .B(n157), .Z(\ab[16][39] ) );
  NR2 U3762 ( .A(n492), .B(n5), .Z(\ab[15][95] ) );
  NR2 U3763 ( .A(n493), .B(n5), .Z(\ab[15][94] ) );
  NR2 U3764 ( .A(n494), .B(n5), .Z(\ab[15][93] ) );
  NR2 U3765 ( .A(n495), .B(n5), .Z(\ab[15][92] ) );
  NR2 U3766 ( .A(n496), .B(n5), .Z(\ab[15][91] ) );
  NR2 U3767 ( .A(n497), .B(n5), .Z(\ab[15][90] ) );
  NR2 U3768 ( .A(n498), .B(n5), .Z(\ab[15][89] ) );
  NR2 U3769 ( .A(n499), .B(n5), .Z(\ab[15][88] ) );
  NR2 U3770 ( .A(n500), .B(n5), .Z(\ab[15][87] ) );
  NR2 U3771 ( .A(n501), .B(n5), .Z(\ab[15][86] ) );
  NR2 U3772 ( .A(n502), .B(n5), .Z(\ab[15][85] ) );
  NR2 U3773 ( .A(n503), .B(n5), .Z(\ab[15][84] ) );
  NR2 U3774 ( .A(n504), .B(n6), .Z(\ab[15][83] ) );
  NR2 U3775 ( .A(n505), .B(n6), .Z(\ab[15][82] ) );
  NR2 U3776 ( .A(n506), .B(n6), .Z(\ab[15][81] ) );
  NR2 U3777 ( .A(n507), .B(n6), .Z(\ab[15][80] ) );
  NR2 U3778 ( .A(n508), .B(n6), .Z(\ab[15][79] ) );
  NR2 U3779 ( .A(n509), .B(n6), .Z(\ab[15][78] ) );
  NR2 U3780 ( .A(n510), .B(n6), .Z(\ab[15][77] ) );
  NR2 U3781 ( .A(n511), .B(n6), .Z(\ab[15][76] ) );
  NR2 U3782 ( .A(n512), .B(n6), .Z(\ab[15][75] ) );
  NR2 U3783 ( .A(n513), .B(n6), .Z(\ab[15][74] ) );
  NR2 U3784 ( .A(n514), .B(n6), .Z(\ab[15][73] ) );
  NR2 U3785 ( .A(n515), .B(n6), .Z(\ab[15][72] ) );
  NR2 U3786 ( .A(n516), .B(n7), .Z(\ab[15][71] ) );
  NR2 U3787 ( .A(n517), .B(n7), .Z(\ab[15][70] ) );
  NR2 U3788 ( .A(n518), .B(n7), .Z(\ab[15][69] ) );
  NR2 U3789 ( .A(n519), .B(n7), .Z(\ab[15][68] ) );
  NR2 U3790 ( .A(n520), .B(n7), .Z(\ab[15][67] ) );
  NR2 U3791 ( .A(n521), .B(n7), .Z(\ab[15][66] ) );
  NR2 U3792 ( .A(n522), .B(n7), .Z(\ab[15][65] ) );
  NR2 U3793 ( .A(n523), .B(n7), .Z(\ab[15][64] ) );
  NR2 U3794 ( .A(n524), .B(n7), .Z(\ab[15][63] ) );
  NR2 U3795 ( .A(n525), .B(n7), .Z(\ab[15][62] ) );
  NR2 U3796 ( .A(n526), .B(n7), .Z(\ab[15][61] ) );
  NR2 U3797 ( .A(n527), .B(n7), .Z(\ab[15][60] ) );
  NR2 U3798 ( .A(n528), .B(n8), .Z(\ab[15][59] ) );
  NR2 U3799 ( .A(n529), .B(n8), .Z(\ab[15][58] ) );
  NR2 U3800 ( .A(n530), .B(n8), .Z(\ab[15][57] ) );
  NR2 U3801 ( .A(n531), .B(n8), .Z(\ab[15][56] ) );
  NR2 U3802 ( .A(n532), .B(n8), .Z(\ab[15][55] ) );
  NR2 U3803 ( .A(n533), .B(n8), .Z(\ab[15][54] ) );
  NR2 U3804 ( .A(n534), .B(n8), .Z(\ab[15][53] ) );
  NR2 U3805 ( .A(n535), .B(n8), .Z(\ab[15][52] ) );
  NR2 U3806 ( .A(n536), .B(n8), .Z(\ab[15][51] ) );
  NR2 U3807 ( .A(n537), .B(n8), .Z(\ab[15][50] ) );
  NR2 U3808 ( .A(n538), .B(n8), .Z(\ab[15][49] ) );
  NR2 U3809 ( .A(n539), .B(n8), .Z(\ab[15][48] ) );
  NR2 U3810 ( .A(n540), .B(n9), .Z(\ab[15][47] ) );
  NR2 U3811 ( .A(n541), .B(n9), .Z(\ab[15][46] ) );
  NR2 U3812 ( .A(n542), .B(n9), .Z(\ab[15][45] ) );
  NR2 U3813 ( .A(n543), .B(n9), .Z(\ab[15][44] ) );
  NR2 U3814 ( .A(n544), .B(n9), .Z(\ab[15][43] ) );
  NR2 U3815 ( .A(n545), .B(n9), .Z(\ab[15][42] ) );
  NR2 U3816 ( .A(n546), .B(n9), .Z(\ab[15][41] ) );
  NR2 U3817 ( .A(n547), .B(n9), .Z(\ab[15][40] ) );
  NR2 U3818 ( .A(n548), .B(n9), .Z(\ab[15][39] ) );
endmodule


module LOG_POLY_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:0] carry;

  EO3P U2_6 ( .A(A[6]), .B(n3), .C(carry[6]), .Z(DIFF[6]) );
  FA1A U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1A U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1A U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1A U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA1A U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  IVP U1 ( .A(A[0]), .Z(n1) );
  EN U2 ( .A(A[0]), .B(n9), .Z(DIFF[0]) );
  IVP U3 ( .A(B[1]), .Z(n8) );
  ND2 U4 ( .A(n1), .B(n2), .Z(carry[1]) );
  IVP U5 ( .A(n9), .Z(n2) );
  IVP U6 ( .A(B[2]), .Z(n7) );
  IVP U7 ( .A(B[3]), .Z(n6) );
  IVP U8 ( .A(B[4]), .Z(n5) );
  IVP U9 ( .A(B[5]), .Z(n4) );
  IVP U10 ( .A(B[6]), .Z(n3) );
  IVP U11 ( .A(B[0]), .Z(n9) );
endmodule


module LOG_POLY_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [24:0] carry;

  FA1A U2_22 ( .A(A[22]), .B(n3), .CI(carry[22]), .CO(carry[23]), .S(DIFF[22])
         );
  FA1A U2_21 ( .A(A[21]), .B(n4), .CI(carry[21]), .CO(carry[22]), .S(DIFF[21])
         );
  FA1A U2_20 ( .A(A[20]), .B(n5), .CI(carry[20]), .CO(carry[21]), .S(DIFF[20])
         );
  FA1A U2_19 ( .A(A[19]), .B(n6), .CI(carry[19]), .CO(carry[20]), .S(DIFF[19])
         );
  FA1A U2_18 ( .A(A[18]), .B(n7), .CI(carry[18]), .CO(carry[19]), .S(DIFF[18])
         );
  FA1A U2_17 ( .A(A[17]), .B(n8), .CI(carry[17]), .CO(carry[18]), .S(DIFF[17])
         );
  FA1A U2_16 ( .A(A[16]), .B(n9), .CI(carry[16]), .CO(carry[17]), .S(DIFF[16])
         );
  FA1A U2_15 ( .A(A[15]), .B(n10), .CI(carry[15]), .CO(carry[16]), .S(DIFF[15]) );
  FA1A U2_14 ( .A(A[14]), .B(n11), .CI(carry[14]), .CO(carry[15]), .S(DIFF[14]) );
  FA1A U2_13 ( .A(A[13]), .B(n12), .CI(carry[13]), .CO(carry[14]), .S(DIFF[13]) );
  FA1A U2_12 ( .A(A[12]), .B(n13), .CI(carry[12]), .CO(carry[13]), .S(DIFF[12]) );
  FA1A U2_11 ( .A(A[11]), .B(n14), .CI(carry[11]), .CO(carry[12]), .S(DIFF[11]) );
  FA1A U2_10 ( .A(A[10]), .B(n15), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  FA1A U2_9 ( .A(A[9]), .B(n16), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]) );
  FA1A U2_8 ( .A(A[8]), .B(n17), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA1A U2_7 ( .A(A[7]), .B(n18), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA1A U2_6 ( .A(A[6]), .B(n19), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1A U2_5 ( .A(A[5]), .B(n20), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1A U2_4 ( .A(A[4]), .B(n21), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1A U2_3 ( .A(A[3]), .B(n22), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1A U2_2 ( .A(A[2]), .B(n23), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA1A U2_1 ( .A(A[1]), .B(n24), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  EN U1 ( .A(A[23]), .B(carry[23]), .Z(DIFF[23]) );
  IVP U2 ( .A(n25), .Z(n2) );
  IVP U3 ( .A(B[0]), .Z(n25) );
  ND2 U4 ( .A(n1), .B(n2), .Z(carry[1]) );
  IVP U5 ( .A(B[1]), .Z(n24) );
  IVP U6 ( .A(A[0]), .Z(n1) );
  IVP U7 ( .A(B[2]), .Z(n23) );
  IVP U8 ( .A(B[3]), .Z(n22) );
  IVP U9 ( .A(B[4]), .Z(n21) );
  IVP U10 ( .A(B[5]), .Z(n20) );
  IVP U11 ( .A(B[6]), .Z(n19) );
  IVP U12 ( .A(B[7]), .Z(n18) );
  IVP U13 ( .A(B[8]), .Z(n17) );
  IVP U14 ( .A(B[9]), .Z(n16) );
  IVP U15 ( .A(B[10]), .Z(n15) );
  IVP U16 ( .A(B[11]), .Z(n14) );
  IVP U17 ( .A(B[12]), .Z(n13) );
  IVP U18 ( .A(B[13]), .Z(n12) );
  IVP U19 ( .A(B[14]), .Z(n11) );
  IVP U20 ( .A(B[15]), .Z(n10) );
  IVP U21 ( .A(B[16]), .Z(n9) );
  IVP U22 ( .A(B[17]), .Z(n8) );
  IVP U23 ( .A(B[18]), .Z(n7) );
  IVP U24 ( .A(B[19]), .Z(n6) );
  IVP U25 ( .A(B[20]), .Z(n5) );
  IVP U26 ( .A(B[21]), .Z(n4) );
  IVP U27 ( .A(B[22]), .Z(n3) );
  EN U28 ( .A(A[0]), .B(n25), .Z(DIFF[0]) );
endmodule


module LOG_POLY_DW01_add_5 ( A, B, CI, SUM, CO );
  input [93:0] A;
  input [93:0] B;
  output [93:0] SUM;
  input CI;
  output CO;
  wire   \A[46] , \A[45] , \A[44] , \A[43] , \A[42] , \A[41] , \A[40] ,
         \A[39] , \A[38] , \A[37] , \A[36] , \A[35] , \A[34] , \A[33] ,
         \A[32] , \A[31] , \A[30] , \A[29] , \A[28] , \A[27] , \A[26] ,
         \A[25] , \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] ,
         \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] ,
         \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] ,
         \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474;
  assign SUM[46] = \A[46] ;
  assign \A[46]  = A[46];
  assign SUM[45] = \A[45] ;
  assign \A[45]  = A[45];
  assign SUM[44] = \A[44] ;
  assign \A[44]  = A[44];
  assign SUM[43] = \A[43] ;
  assign \A[43]  = A[43];
  assign SUM[42] = \A[42] ;
  assign \A[42]  = A[42];
  assign SUM[41] = \A[41] ;
  assign \A[41]  = A[41];
  assign SUM[40] = \A[40] ;
  assign \A[40]  = A[40];
  assign SUM[39] = \A[39] ;
  assign \A[39]  = A[39];
  assign SUM[38] = \A[38] ;
  assign \A[38]  = A[38];
  assign SUM[37] = \A[37] ;
  assign \A[37]  = A[37];
  assign SUM[36] = \A[36] ;
  assign \A[36]  = A[36];
  assign SUM[35] = \A[35] ;
  assign \A[35]  = A[35];
  assign SUM[34] = \A[34] ;
  assign \A[34]  = A[34];
  assign SUM[33] = \A[33] ;
  assign \A[33]  = A[33];
  assign SUM[32] = \A[32] ;
  assign \A[32]  = A[32];
  assign SUM[31] = \A[31] ;
  assign \A[31]  = A[31];
  assign SUM[30] = \A[30] ;
  assign \A[30]  = A[30];
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  IVAP U2 ( .A(n405), .Z(n404) );
  ND2P U3 ( .A(n415), .B(n416), .Z(n403) );
  IV U4 ( .A(n136), .Z(n135) );
  ND2 U5 ( .A(n388), .B(n41), .Z(n379) );
  AN3P U6 ( .A(n355), .B(n381), .C(n356), .Z(n3) );
  ND2P U7 ( .A(n434), .B(n425), .Z(n432) );
  ND2P U8 ( .A(n269), .B(n5), .Z(n293) );
  ND2 U9 ( .A(n223), .B(n224), .Z(n1) );
  IVAP U10 ( .A(B[78]), .Z(n250) );
  ND2 U11 ( .A(n302), .B(n303), .Z(n2) );
  AO2P U12 ( .A(B[58]), .B(A[58]), .C(B[59]), .D(A[59]), .Z(n397) );
  IVP U13 ( .A(n323), .Z(n310) );
  ND4P U14 ( .A(n327), .B(n49), .C(n328), .D(n329), .Z(n323) );
  ND2P U15 ( .A(n382), .B(n34), .Z(n380) );
  ND2P U16 ( .A(n210), .B(n211), .Z(n197) );
  ND2P U17 ( .A(n62), .B(n105), .Z(n94) );
  IV U18 ( .A(n209), .Z(n207) );
  AO7P U19 ( .A(n86), .B(n87), .C(n88), .Z(n85) );
  ND2P U20 ( .A(n447), .B(n448), .Z(n363) );
  AO3 U21 ( .A(n96), .B(n97), .C(n98), .D(n99), .Z(n104) );
  ND2 U22 ( .A(n357), .B(n358), .Z(n331) );
  NR2P U23 ( .A(n364), .B(n365), .Z(n361) );
  IVA U24 ( .A(n205), .Z(n221) );
  IVAP U25 ( .A(A[82]), .Z(n181) );
  ND3P U26 ( .A(n361), .B(n362), .C(n363), .Z(n39) );
  IVA U27 ( .A(A[80]), .Z(n193) );
  EOP U28 ( .A(n252), .B(n253), .Z(SUM[77]) );
  IV U29 ( .A(n247), .Z(n254) );
  AO7P U30 ( .A(n212), .B(n213), .C(n5), .Z(n211) );
  IVP U31 ( .A(n37), .Z(n38) );
  IVDAP U32 ( .A(A[74]), .Y(n37), .Z(n40) );
  ND2 U33 ( .A(n267), .B(n268), .Z(n261) );
  ND4P U34 ( .A(n220), .B(n221), .C(n222), .D(n352), .Z(n141) );
  ND2P U35 ( .A(n446), .B(n428), .Z(n443) );
  AN2 U36 ( .A(n237), .B(n223), .Z(n20) );
  OR2P U37 ( .A(A[74]), .B(B[74]), .Z(n270) );
  OR2P U38 ( .A(n141), .B(n142), .Z(n194) );
  IVP U39 ( .A(n206), .Z(n201) );
  OR2 U40 ( .A(A[50]), .B(B[50]), .Z(n36) );
  NR2P U41 ( .A(n228), .B(n229), .Z(n220) );
  OR2P U42 ( .A(A[49]), .B(B[49]), .Z(n446) );
  NR2P U43 ( .A(A[49]), .B(B[49]), .Z(n453) );
  IV U44 ( .A(n287), .Z(n284) );
  EOP U45 ( .A(n343), .B(n342), .Z(SUM[66]) );
  OR2 U46 ( .A(n196), .B(n195), .Z(n139) );
  ND2 U47 ( .A(B[77]), .B(A[77]), .Z(n217) );
  ND2 U48 ( .A(n36), .B(n445), .Z(n444) );
  IVAP U49 ( .A(A[81]), .Z(n189) );
  ND3P U50 ( .A(n355), .B(n16), .C(n356), .Z(n328) );
  NR2P U51 ( .A(B[60]), .B(A[60]), .Z(n16) );
  IV U52 ( .A(n104), .Z(n86) );
  NR2P U53 ( .A(n449), .B(n450), .Z(n448) );
  NR3P U54 ( .A(n451), .B(n452), .C(n453), .Z(n450) );
  IV U55 ( .A(n133), .Z(n147) );
  IVAP U56 ( .A(n137), .Z(n96) );
  NR2P U57 ( .A(n473), .B(n31), .Z(n51) );
  ND2P U58 ( .A(n397), .B(n27), .Z(n388) );
  IV U59 ( .A(n473), .Z(n471) );
  ND2P U60 ( .A(B[87]), .B(A[87]), .Z(n129) );
  ND2P U61 ( .A(n192), .B(n193), .Z(n186) );
  AN2 U62 ( .A(n126), .B(n127), .Z(n4) );
  IV U63 ( .A(n120), .Z(n124) );
  ND2P U64 ( .A(n120), .B(n117), .Z(n118) );
  AO7P U65 ( .A(n128), .B(n129), .C(n130), .Z(n120) );
  IV U66 ( .A(n108), .Z(n110) );
  ND2P U67 ( .A(n108), .B(n105), .Z(n106) );
  AO7P U68 ( .A(n113), .B(n59), .C(n114), .Z(n108) );
  IVP U69 ( .A(A[56]), .Z(n416) );
  IVP U70 ( .A(B[56]), .Z(n415) );
  IVP U71 ( .A(B[81]), .Z(n188) );
  ND4 U72 ( .A(n389), .B(n399), .C(n402), .D(n403), .Z(n25) );
  ND2 U73 ( .A(n420), .B(n28), .Z(n372) );
  ND3 U74 ( .A(n157), .B(n158), .C(n159), .Z(n152) );
  ND2 U75 ( .A(n148), .B(n149), .Z(n133) );
  ND3 U76 ( .A(n150), .B(n151), .C(n152), .Z(n148) );
  IVP U77 ( .A(B[80]), .Z(n192) );
  EO U78 ( .A(n457), .B(n458), .Z(SUM[51]) );
  EN U79 ( .A(n410), .B(n52), .Z(SUM[58]) );
  EN U80 ( .A(n317), .B(n66), .Z(SUM[69]) );
  EO U81 ( .A(n295), .B(n296), .Z(SUM[72]) );
  EO U82 ( .A(n288), .B(n289), .Z(SUM[73]) );
  EO U83 ( .A(n282), .B(n283), .Z(SUM[74]) );
  EO U84 ( .A(n314), .B(n60), .Z(SUM[70]) );
  EN U85 ( .A(n406), .B(n407), .Z(SUM[59]) );
  EN U86 ( .A(n95), .B(n76), .Z(SUM[87]) );
  EN U87 ( .A(n179), .B(n78), .Z(SUM[82]) );
  EN U88 ( .A(n171), .B(n79), .Z(SUM[83]) );
  EO U89 ( .A(n57), .B(n80), .Z(SUM[62]) );
  EN U90 ( .A(n187), .B(n81), .Z(SUM[81]) );
  EN U91 ( .A(n162), .B(n163), .Z(SUM[84]) );
  EN U92 ( .A(n155), .B(n82), .Z(SUM[85]) );
  EN U93 ( .A(n143), .B(n83), .Z(SUM[86]) );
  EN U94 ( .A(n313), .B(n84), .Z(SUM[71]) );
  OR2P U95 ( .A(B[71]), .B(A[71]), .Z(n5) );
  AN2P U96 ( .A(n424), .B(n425), .Z(n6) );
  IVDA U97 ( .A(n321), .Y(n7), .Z(n8) );
  IVDA U98 ( .A(n302), .Y(n9), .Z(n10) );
  IVDA U99 ( .A(n305), .Y(n11), .Z(n12) );
  IVDA U100 ( .A(n446), .Y(n13), .Z(n14) );
  IVDA U101 ( .A(n16), .Y(n15), .Z(n42) );
  ND2 U102 ( .A(n374), .B(n375), .Z(n371) );
  OR2 U103 ( .A(A[58]), .B(B[58]), .Z(n399) );
  OR2 U104 ( .A(A[58]), .B(B[58]), .Z(n17) );
  NR2P U105 ( .A(A[50]), .B(B[50]), .Z(n452) );
  ND2 U106 ( .A(n463), .B(n445), .Z(n18) );
  IV U107 ( .A(A[57]), .Z(n412) );
  B5I U108 ( .A(n227), .Z(n216) );
  ND2 U109 ( .A(n311), .B(n235), .Z(n309) );
  IVDA U110 ( .A(n385), .Z(n21) );
  IV U111 ( .A(B[57]), .Z(n411) );
  ND2 U112 ( .A(n446), .B(n428), .Z(n22) );
  IVDA U113 ( .A(n387), .Z(n23) );
  ND2 U114 ( .A(n411), .B(n412), .Z(n402) );
  IVDA U115 ( .A(n399), .Z(n24) );
  IV U116 ( .A(n142), .Z(n297) );
  NR2 U117 ( .A(A[58]), .B(B[58]), .Z(n26) );
  NR2 U118 ( .A(n215), .B(n206), .Z(n210) );
  OR2 U119 ( .A(A[55]), .B(B[55]), .Z(n28) );
  B5I U120 ( .A(n422), .Z(n420) );
  AN2P U121 ( .A(n411), .B(n412), .Z(n27) );
  ND2 U122 ( .A(n420), .B(n421), .Z(n29) );
  B3I U123 ( .A(A[69]), .Z1(n319) );
  IVDA U124 ( .A(n271), .Z(n30) );
  ND2P U125 ( .A(B[74]), .B(n38), .Z(n268) );
  OR2 U126 ( .A(n22), .B(n18), .Z(n31) );
  OR2 U127 ( .A(n22), .B(n18), .Z(n32) );
  ND4P U128 ( .A(n384), .B(n385), .C(n386), .D(n387), .Z(n382) );
  OR2P U129 ( .A(B[65]), .B(A[65]), .Z(n337) );
  IV U130 ( .A(n270), .Z(n281) );
  ND2 U131 ( .A(n447), .B(n448), .Z(n33) );
  ND2 U132 ( .A(n26), .B(n398), .Z(n34) );
  ND2 U133 ( .A(n26), .B(n398), .Z(n383) );
  OR2P U134 ( .A(B[66]), .B(A[66]), .Z(n338) );
  IV U135 ( .A(n362), .Z(n35) );
  OR2P U136 ( .A(A[48]), .B(B[48]), .Z(n445) );
  ND4P U137 ( .A(B[64]), .B(A[64]), .C(n337), .D(n338), .Z(n335) );
  NR2P U138 ( .A(n330), .B(n47), .Z(n329) );
  ND2P U139 ( .A(n238), .B(n20), .Z(n233) );
  ND2P U140 ( .A(n339), .B(n232), .Z(n334) );
  B5I U141 ( .A(n368), .Z(n362) );
  ND2P U142 ( .A(n318), .B(n319), .Z(n303) );
  B5I U143 ( .A(B[69]), .Z(n318) );
  IVDA U144 ( .A(n427), .Y(n437), .Z(n19) );
  ND3P U145 ( .A(n231), .B(n230), .C(n232), .Z(n330) );
  ND3 U146 ( .A(n361), .B(n362), .C(n363), .Z(n238) );
  ND4P U147 ( .A(n383), .B(n388), .C(n41), .D(n382), .Z(n237) );
  OR2 U148 ( .A(A[59]), .B(B[59]), .Z(n41) );
  OR2 U149 ( .A(A[59]), .B(B[59]), .Z(n389) );
  ND2 U150 ( .A(B[57]), .B(A[57]), .Z(n387) );
  NR2P U151 ( .A(n473), .B(n25), .Z(n367) );
  NR2 U152 ( .A(n233), .B(n234), .Z(n43) );
  ND2 U153 ( .A(n415), .B(n416), .Z(n44) );
  ND2 U154 ( .A(n58), .B(n249), .Z(n248) );
  ND2 U155 ( .A(B[63]), .B(A[63]), .Z(n223) );
  ND2P U156 ( .A(n318), .B(n319), .Z(n45) );
  ND2 U157 ( .A(n318), .B(n319), .Z(n46) );
  ND2P U158 ( .A(n223), .B(n224), .Z(n352) );
  IVP U159 ( .A(n161), .Z(n160) );
  AO3P U160 ( .A(n96), .B(n97), .C(n98), .D(n99), .Z(n95) );
  OR2P U161 ( .A(B[70]), .B(A[70]), .Z(n302) );
  IVDAP U162 ( .A(n331), .Y(n48), .Z(n47) );
  IV U163 ( .A(A[78]), .Z(n251) );
  ND2 U164 ( .A(B[69]), .B(A[69]), .Z(n305) );
  OR2P U165 ( .A(B[62]), .B(A[62]), .Z(n357) );
  AO6P U166 ( .A(n46), .B(n315), .C(n11), .Z(n314) );
  IVA U167 ( .A(B[76]), .Z(n273) );
  OR2P U168 ( .A(B[63]), .B(A[63]), .Z(n358) );
  ND4 U169 ( .A(n311), .B(n235), .C(n236), .D(n39), .Z(n321) );
  AO7P U170 ( .A(n391), .B(n57), .C(n356), .Z(n390) );
  AO6P U171 ( .A(n201), .B(n195), .C(n202), .Z(n200) );
  ND3P U172 ( .A(n235), .B(n3), .C(n236), .Z(n234) );
  NR2P U173 ( .A(n365), .B(n69), .Z(n366) );
  ND4P U174 ( .A(n225), .B(n226), .C(n227), .D(n203), .Z(n195) );
  AO6P U175 ( .A(n279), .B(n280), .C(n281), .Z(n278) );
  NR2P U176 ( .A(n277), .B(n278), .Z(n276) );
  IVP U177 ( .A(n170), .Z(n169) );
  IV U178 ( .A(n306), .Z(n320) );
  OR2P U179 ( .A(A[54]), .B(B[54]), .Z(n426) );
  AO7P U180 ( .A(n55), .B(n2), .C(n299), .Z(n269) );
  IVA U181 ( .A(n213), .Z(n299) );
  AO3 U182 ( .A(n351), .B(n321), .C(n1), .D(n230), .Z(n347) );
  AO7 U183 ( .A(n27), .B(n56), .C(n387), .Z(n409) );
  AO7P U184 ( .A(n51), .B(n33), .C(n404), .Z(n401) );
  ND2 U185 ( .A(B[71]), .B(A[71]), .Z(n300) );
  ND2P U186 ( .A(n122), .B(n123), .Z(n117) );
  IVP U187 ( .A(A[89]), .Z(n123) );
  IV U188 ( .A(B[86]), .Z(n144) );
  IV U189 ( .A(n346), .Z(n345) );
  AN2P U190 ( .A(n392), .B(n355), .Z(n57) );
  AO7 U191 ( .A(n417), .B(n405), .C(n400), .Z(n414) );
  EO U192 ( .A(n56), .B(n61), .Z(SUM[57]) );
  ND2 U193 ( .A(n462), .B(n463), .Z(n461) );
  AN2P U194 ( .A(n118), .B(n119), .Z(n59) );
  ND3 U195 ( .A(n166), .B(n167), .C(n168), .Z(n159) );
  ND2 U196 ( .A(n175), .B(n176), .Z(n168) );
  ND2 U197 ( .A(n106), .B(n107), .Z(n89) );
  OR2 U198 ( .A(B[88]), .B(A[88]), .Z(n127) );
  IVA U199 ( .A(B[89]), .Z(n122) );
  ND2 U200 ( .A(n333), .B(n232), .Z(n343) );
  AO3P U201 ( .A(n284), .B(n249), .C(n30), .D(n285), .Z(n279) );
  IVDA U202 ( .A(n217), .Y(n243) );
  IV U203 ( .A(n286), .Z(n290) );
  AN2 U204 ( .A(n63), .B(n112), .Z(n62) );
  AN2 U205 ( .A(n4), .B(n117), .Z(n63) );
  AN2 U206 ( .A(n53), .B(n225), .Z(n58) );
  AO7P U207 ( .A(n13), .B(n465), .C(n466), .Z(n462) );
  IVP U208 ( .A(n467), .Z(n465) );
  AO7P U209 ( .A(n332), .B(n209), .C(n49), .Z(n306) );
  ND2P U210 ( .A(n359), .B(n356), .Z(n327) );
  OR2P U211 ( .A(B[68]), .B(A[68]), .Z(n312) );
  OR2P U212 ( .A(B[67]), .B(A[67]), .Z(n49) );
  OR2P U213 ( .A(B[85]), .B(A[85]), .Z(n151) );
  OR2P U214 ( .A(B[61]), .B(A[61]), .Z(n360) );
  IV U215 ( .A(A[86]), .Z(n145) );
  OR2P U216 ( .A(B[79]), .B(A[79]), .Z(n203) );
  OR2P U217 ( .A(B[75]), .B(A[75]), .Z(n263) );
  IVA U218 ( .A(n474), .Z(SUM[47]) );
  EOP U219 ( .A(n275), .B(n276), .Z(SUM[75]) );
  ENP U220 ( .A(n340), .B(n77), .Z(SUM[67]) );
  ENP U221 ( .A(n131), .B(n70), .Z(SUM[88]) );
  ENP U222 ( .A(n121), .B(n71), .Z(SUM[89]) );
  ENP U223 ( .A(n115), .B(n72), .Z(SUM[90]) );
  ENP U224 ( .A(n109), .B(n73), .Z(SUM[91]) );
  ENP U225 ( .A(n100), .B(n74), .Z(SUM[92]) );
  ENP U226 ( .A(n390), .B(n75), .Z(SUM[63]) );
  EOP U227 ( .A(n85), .B(B[93]), .Z(SUM[93]) );
  ENP U228 ( .A(n244), .B(n245), .Z(SUM[78]) );
  ENP U229 ( .A(n239), .B(n240), .Z(SUM[79]) );
  AO3P U230 ( .A(n96), .B(n97), .C(n98), .D(n99), .Z(n50) );
  AO6P U231 ( .A(n231), .B(n344), .C(n345), .Z(n342) );
  OR2P U232 ( .A(n443), .B(n444), .Z(n69) );
  AO7 U233 ( .A(n27), .B(n56), .C(n23), .Z(n52) );
  AO7 U234 ( .A(n146), .B(n136), .C(n147), .Z(n143) );
  NR2 U235 ( .A(n142), .B(n205), .Z(n53) );
  ND2 U236 ( .A(n286), .B(n287), .Z(n285) );
  IV U237 ( .A(n237), .Z(n396) );
  AO3 U238 ( .A(n320), .B(n321), .C(n322), .D(n312), .Z(n316) );
  ND2 U239 ( .A(n168), .B(n167), .Z(n174) );
  ND2 U240 ( .A(n246), .B(n226), .Z(n241) );
  ND2 U241 ( .A(n247), .B(n248), .Z(n246) );
  ND2 U242 ( .A(n291), .B(n272), .Z(n287) );
  ND2 U243 ( .A(n292), .B(n293), .Z(n291) );
  NR2 U244 ( .A(n473), .B(n32), .Z(n54) );
  AN2P U245 ( .A(n304), .B(n305), .Z(n55) );
  AN2P U246 ( .A(n386), .B(n413), .Z(n56) );
  AO7 U247 ( .A(n341), .B(n342), .C(n333), .Z(n340) );
  AO3 U248 ( .A(n216), .B(n241), .C(n219), .D(n242), .Z(n239) );
  AO7 U249 ( .A(n190), .B(n146), .C(n185), .Z(n187) );
  AO3 U250 ( .A(n146), .B(n161), .C(n159), .D(n158), .Z(n162) );
  AO7 U251 ( .A(n146), .B(n154), .C(n156), .Z(n155) );
  ND2 U252 ( .A(n152), .B(n150), .Z(n156) );
  ND2 U253 ( .A(n241), .B(n217), .Z(n245) );
  ND2 U254 ( .A(n408), .B(n21), .Z(n406) );
  ND2 U255 ( .A(n409), .B(n24), .Z(n408) );
  ND2 U256 ( .A(n300), .B(n301), .Z(n213) );
  ND2 U257 ( .A(n260), .B(n196), .Z(n255) );
  ND3 U258 ( .A(n5), .B(n221), .C(n269), .Z(n260) );
  ND2 U259 ( .A(n226), .B(n217), .Z(n252) );
  ND2 U260 ( .A(n10), .B(n301), .Z(n60) );
  NR2 U261 ( .A(n277), .B(n281), .Z(n283) );
  ND2 U262 ( .A(n292), .B(n272), .Z(n295) );
  EO U263 ( .A(n258), .B(n259), .Z(SUM[76]) );
  ND2 U264 ( .A(n402), .B(n23), .Z(n61) );
  ND2 U265 ( .A(n182), .B(n183), .Z(n175) );
  ND2 U266 ( .A(n184), .B(n185), .Z(n182) );
  EN U267 ( .A(n191), .B(n64), .Z(SUM[80]) );
  ND2 U268 ( .A(n185), .B(n186), .Z(n64) );
  EN U269 ( .A(n393), .B(n65), .Z(SUM[61]) );
  ND2 U270 ( .A(n360), .B(n355), .Z(n65) );
  EN U271 ( .A(n349), .B(n350), .Z(SUM[65]) );
  ND2 U272 ( .A(n346), .B(n231), .Z(n350) );
  ND2 U273 ( .A(n348), .B(n347), .Z(n349) );
  ND2 U274 ( .A(n45), .B(n12), .Z(n66) );
  EN U275 ( .A(n353), .B(n354), .Z(SUM[64]) );
  EO U276 ( .A(n324), .B(n325), .Z(SUM[68]) );
  ND2 U277 ( .A(n310), .B(n8), .Z(n326) );
  EO U278 ( .A(n394), .B(n67), .Z(SUM[60]) );
  ND2 U279 ( .A(n15), .B(n381), .Z(n67) );
  ND2 U280 ( .A(n469), .B(n470), .Z(n467) );
  EN U281 ( .A(n414), .B(n68), .Z(SUM[56]) );
  ND2 U282 ( .A(n44), .B(n386), .Z(n68) );
  EN U283 ( .A(n464), .B(n462), .Z(SUM[50]) );
  ND2 U284 ( .A(n455), .B(n463), .Z(n464) );
  EN U285 ( .A(n440), .B(n439), .Z(SUM[52]) );
  EN U286 ( .A(n468), .B(n467), .Z(SUM[49]) );
  ND2 U287 ( .A(n466), .B(n14), .Z(n468) );
  EO U288 ( .A(n472), .B(n473), .Z(SUM[48]) );
  ND2 U289 ( .A(n376), .B(n377), .Z(n374) );
  AO3 U290 ( .A(n6), .B(n419), .C(n373), .D(n29), .Z(n418) );
  ND2 U291 ( .A(B[70]), .B(A[70]), .Z(n301) );
  ND2 U292 ( .A(B[52]), .B(A[52]), .Z(n376) );
  EN U293 ( .A(n429), .B(n430), .Z(SUM[55]) );
  ND2 U294 ( .A(n28), .B(n373), .Z(n430) );
  ND2 U295 ( .A(n422), .B(n431), .Z(n429) );
  AO7 U296 ( .A(n261), .B(n262), .C(n263), .Z(n196) );
  AO7 U297 ( .A(n264), .B(n265), .C(n266), .Z(n262) );
  ND2 U298 ( .A(B[72]), .B(A[72]), .Z(n265) );
  IV U299 ( .A(B[77]), .Z(n256) );
  IV U300 ( .A(B[83]), .Z(n172) );
  ND2 U301 ( .A(B[52]), .B(A[52]), .Z(n424) );
  ND2 U302 ( .A(B[78]), .B(A[78]), .Z(n219) );
  ND2 U303 ( .A(B[60]), .B(A[60]), .Z(n381) );
  ND2 U304 ( .A(B[80]), .B(A[80]), .Z(n185) );
  ND2 U305 ( .A(B[58]), .B(A[58]), .Z(n385) );
  ND2 U306 ( .A(B[59]), .B(A[59]), .Z(n384) );
  ND2 U307 ( .A(B[59]), .B(A[59]), .Z(n398) );
  ND2 U308 ( .A(B[75]), .B(A[75]), .Z(n267) );
  ND2 U309 ( .A(B[79]), .B(A[79]), .Z(n218) );
  ND2 U310 ( .A(B[76]), .B(A[76]), .Z(n204) );
  ND2 U311 ( .A(B[67]), .B(A[67]), .Z(n336) );
  ND2 U312 ( .A(B[81]), .B(A[81]), .Z(n184) );
  IV U313 ( .A(B[82]), .Z(n180) );
  EN U314 ( .A(n433), .B(n432), .Z(SUM[54]) );
  IV U315 ( .A(B[84]), .Z(n164) );
  OR2 U316 ( .A(B[90]), .B(A[90]), .Z(n112) );
  ND2 U317 ( .A(B[84]), .B(A[84]), .Z(n157) );
  ND2 U318 ( .A(B[82]), .B(A[82]), .Z(n176) );
  OR2 U319 ( .A(B[87]), .B(A[87]), .Z(n126) );
  ND2 U320 ( .A(B[89]), .B(A[89]), .Z(n119) );
  ND2 U321 ( .A(B[90]), .B(A[90]), .Z(n114) );
  EN U322 ( .A(n436), .B(n435), .Z(SUM[53]) );
  ND2 U323 ( .A(B[83]), .B(A[83]), .Z(n158) );
  ND2 U324 ( .A(B[72]), .B(A[72]), .Z(n292) );
  ND2 U325 ( .A(B[86]), .B(A[86]), .Z(n99) );
  ND2 U326 ( .A(B[49]), .B(A[49]), .Z(n466) );
  ND2 U327 ( .A(B[73]), .B(A[73]), .Z(n280) );
  ND2 U328 ( .A(B[85]), .B(A[85]), .Z(n149) );
  AO6 U329 ( .A(n89), .B(n90), .C(n91), .Z(n88) );
  OR2 U330 ( .A(B[91]), .B(A[91]), .Z(n105) );
  ND2 U331 ( .A(B[91]), .B(A[91]), .Z(n107) );
  OR2 U332 ( .A(B[92]), .B(A[92]), .Z(n90) );
  ND2 U333 ( .A(B[92]), .B(A[92]), .Z(n92) );
  ND2 U334 ( .A(n41), .B(n398), .Z(n407) );
  ND2 U335 ( .A(n127), .B(n130), .Z(n70) );
  ND2 U336 ( .A(n117), .B(n119), .Z(n71) );
  ND2 U337 ( .A(n112), .B(n114), .Z(n72) );
  ND2 U338 ( .A(n105), .B(n107), .Z(n73) );
  ND2 U339 ( .A(n92), .B(n90), .Z(n74) );
  ND2 U340 ( .A(n358), .B(n223), .Z(n75) );
  ND2 U341 ( .A(n126), .B(n129), .Z(n76) );
  ND2 U342 ( .A(n336), .B(n49), .Z(n77) );
  ND2 U343 ( .A(n176), .B(n167), .Z(n78) );
  ND2 U344 ( .A(n158), .B(n166), .Z(n79) );
  ND2 U345 ( .A(n218), .B(n203), .Z(n240) );
  ND2 U346 ( .A(n357), .B(n356), .Z(n80) );
  ND2 U347 ( .A(n184), .B(n183), .Z(n81) );
  ND2 U348 ( .A(n157), .B(n150), .Z(n163) );
  ND2 U349 ( .A(n151), .B(n149), .Z(n82) );
  ND2 U350 ( .A(n134), .B(n99), .Z(n83) );
  ND2 U351 ( .A(n267), .B(n263), .Z(n275) );
  ND2 U352 ( .A(n300), .B(n5), .Z(n84) );
  IVP U353 ( .A(n428), .Z(n364) );
  ND2 U354 ( .A(n33), .B(n428), .Z(n441) );
  AN2 U355 ( .A(n454), .B(n428), .Z(n458) );
  AO7 U356 ( .A(n146), .B(n178), .C(n175), .Z(n179) );
  ND2 U357 ( .A(B[64]), .B(A[64]), .Z(n348) );
  ND2 U358 ( .A(n424), .B(n19), .Z(n440) );
  AO7 U359 ( .A(n146), .B(n170), .C(n174), .Z(n171) );
  ND2 U360 ( .A(B[65]), .B(A[65]), .Z(n346) );
  AN2 U361 ( .A(A[65]), .B(B[65]), .Z(n339) );
  AO3 U362 ( .A(n370), .B(n371), .C(n372), .D(n373), .Z(n369) );
  ND2 U363 ( .A(n230), .B(n231), .Z(n229) );
  AO7 U364 ( .A(A[47]), .B(B[47]), .C(n473), .Z(n474) );
  AO7 U365 ( .A(n7), .B(n224), .C(n223), .Z(n353) );
  OR2P U366 ( .A(A[50]), .B(B[50]), .Z(n463) );
  ND2 U367 ( .A(B[50]), .B(A[50]), .Z(n455) );
  AO3 U368 ( .A(A[50]), .B(B[50]), .C(A[49]), .D(B[49]), .Z(n456) );
  NR2 U369 ( .A(n330), .B(n223), .Z(n332) );
  ND2 U370 ( .A(B[88]), .B(A[88]), .Z(n130) );
  IV U371 ( .A(A[77]), .Z(n257) );
  ND3 U372 ( .A(n204), .B(n205), .C(n201), .Z(n199) );
  ND2 U373 ( .A(B[53]), .B(A[53]), .Z(n425) );
  ND2 U374 ( .A(B[53]), .B(A[53]), .Z(n377) );
  ND2P U375 ( .A(n366), .B(n367), .Z(n236) );
  ND2 U376 ( .A(B[51]), .B(A[51]), .Z(n454) );
  AO7 U377 ( .A(n9), .B(n314), .C(n301), .Z(n313) );
  ND2 U378 ( .A(B[66]), .B(A[66]), .Z(n333) );
  ND2 U379 ( .A(n101), .B(n102), .Z(n100) );
  IVAP U380 ( .A(n178), .Z(n177) );
  ND2 U381 ( .A(B[55]), .B(A[55]), .Z(n373) );
  AO4 U382 ( .A(A[55]), .B(B[55]), .C(A[54]), .D(B[54]), .Z(n370) );
  OR2P U383 ( .A(A[52]), .B(B[52]), .Z(n427) );
  AO3 U384 ( .A(n40), .B(B[74]), .C(A[73]), .D(B[73]), .Z(n266) );
  AO4 U385 ( .A(A[74]), .B(B[74]), .C(A[73]), .D(B[73]), .Z(n264) );
  NR2 U386 ( .A(n54), .B(n33), .Z(n417) );
  ND2 U387 ( .A(n30), .B(n280), .Z(n288) );
  OR2P U388 ( .A(A[53]), .B(B[53]), .Z(n375) );
  IV U389 ( .A(A[76]), .Z(n274) );
  ND2 U390 ( .A(B[61]), .B(A[61]), .Z(n355) );
  ND2 U391 ( .A(n347), .B(n348), .Z(n344) );
  ND2 U392 ( .A(n225), .B(n204), .Z(n258) );
  AO7 U393 ( .A(n215), .B(n255), .C(n225), .Z(n247) );
  ND2 U394 ( .A(n306), .B(n326), .Z(n324) );
  ND2 U395 ( .A(n304), .B(n316), .Z(n317) );
  ND2 U396 ( .A(n348), .B(n230), .Z(n354) );
  ND2 U397 ( .A(n316), .B(n304), .Z(n315) );
  IV U398 ( .A(A[51]), .Z(n460) );
  IVA U399 ( .A(B[51]), .Z(n459) );
  IV U400 ( .A(A[83]), .Z(n173) );
  ND2 U401 ( .A(n445), .B(n469), .Z(n472) );
  ND2 U402 ( .A(n445), .B(n471), .Z(n470) );
  ND2 U403 ( .A(B[48]), .B(A[48]), .Z(n469) );
  ND2 U404 ( .A(B[48]), .B(A[48]), .Z(n451) );
  ND2 U405 ( .A(n110), .B(n111), .Z(n109) );
  IVDA U406 ( .A(n90), .Y(n93) );
  ND2 U407 ( .A(n59), .B(n116), .Z(n115) );
  ND2 U408 ( .A(n124), .B(n125), .Z(n121) );
  ND2 U409 ( .A(n129), .B(n132), .Z(n131) );
  IV U410 ( .A(n89), .Z(n101) );
  ND2P U411 ( .A(n160), .B(n150), .Z(n154) );
  IV U412 ( .A(n151), .Z(n153) );
  IV U413 ( .A(A[84]), .Z(n165) );
  IV U414 ( .A(n94), .Z(n103) );
  IV U415 ( .A(n360), .Z(n359) );
  OR2P U416 ( .A(A[65]), .B(B[65]), .Z(n231) );
  OR2P U417 ( .A(A[64]), .B(B[64]), .Z(n230) );
  IVA U418 ( .A(n195), .Z(n222) );
  OR2P U419 ( .A(A[73]), .B(B[73]), .Z(n271) );
  OR2P U420 ( .A(A[72]), .B(B[72]), .Z(n272) );
  ND2 U421 ( .A(n426), .B(n422), .Z(n433) );
  ND2 U422 ( .A(n432), .B(n426), .Z(n431) );
  OR2P U423 ( .A(A[55]), .B(B[55]), .Z(n421) );
  ND2 U424 ( .A(n227), .B(n219), .Z(n244) );
  ND2 U425 ( .A(n243), .B(n227), .Z(n242) );
  ND2 U426 ( .A(n21), .B(n24), .Z(n410) );
  ND2 U427 ( .A(n279), .B(n280), .Z(n282) );
  AO6 U428 ( .A(n58), .B(n249), .C(n254), .Z(n253) );
  AO6 U429 ( .A(n53), .B(n249), .C(n255), .Z(n259) );
  AO6 U430 ( .A(n290), .B(n249), .C(n284), .Z(n289) );
  AO6 U431 ( .A(n297), .B(n249), .C(n298), .Z(n296) );
  OR2P U432 ( .A(n153), .B(n154), .Z(n136) );
  ND2 U433 ( .A(n425), .B(n375), .Z(n436) );
  ND2 U434 ( .A(n435), .B(n375), .Z(n434) );
  ND2 U435 ( .A(n236), .B(n39), .Z(n308) );
  ND2 U436 ( .A(n375), .B(n423), .Z(n419) );
  OR2P U437 ( .A(n364), .B(n365), .Z(n405) );
  ND2 U438 ( .A(n103), .B(n50), .Z(n102) );
  ND2 U439 ( .A(n62), .B(n50), .Z(n111) );
  ND2 U440 ( .A(n63), .B(n95), .Z(n116) );
  ND2 U441 ( .A(n4), .B(n50), .Z(n125) );
  ND2 U442 ( .A(n95), .B(n126), .Z(n132) );
  AO3 U443 ( .A(n43), .B(n194), .C(n140), .D(n139), .Z(n191) );
  ND2 U444 ( .A(n232), .B(n49), .Z(n228) );
  OR2P U445 ( .A(A[66]), .B(B[66]), .Z(n232) );
  IVA U446 ( .A(n92), .Z(n91) );
  OR2 U447 ( .A(n93), .B(n94), .Z(n87) );
  IVA U448 ( .A(n112), .Z(n113) );
  IVA U449 ( .A(n127), .Z(n128) );
  ND2P U450 ( .A(n133), .B(n134), .Z(n98) );
  ND2P U451 ( .A(n135), .B(n134), .Z(n97) );
  AO3P U452 ( .A(n138), .B(n194), .C(n139), .D(n140), .Z(n137) );
  ND2P U453 ( .A(n144), .B(n145), .Z(n134) );
  ND2P U454 ( .A(n164), .B(n165), .Z(n150) );
  ND2P U455 ( .A(n169), .B(n166), .Z(n161) );
  ND2P U456 ( .A(n172), .B(n173), .Z(n166) );
  ND2P U457 ( .A(n177), .B(n167), .Z(n170) );
  ND2P U458 ( .A(n180), .B(n181), .Z(n167) );
  ND2P U459 ( .A(n186), .B(n183), .Z(n178) );
  ND2P U460 ( .A(n188), .B(n189), .Z(n183) );
  IVA U461 ( .A(n191), .Z(n146) );
  IVA U462 ( .A(n186), .Z(n190) );
  AO3P U463 ( .A(n197), .B(n198), .C(n199), .D(n200), .Z(n140) );
  IVA U464 ( .A(n203), .Z(n202) );
  NR3P U465 ( .A(n207), .B(n208), .C(n142), .Z(n198) );
  IVA U466 ( .A(n49), .Z(n208) );
  NR2P U467 ( .A(n55), .B(n214), .Z(n212) );
  AO3P U468 ( .A(n216), .B(n217), .C(n218), .D(n219), .Z(n206) );
  NR2P U469 ( .A(n233), .B(n234), .Z(n138) );
  ND2P U470 ( .A(n250), .B(n251), .Z(n227) );
  IVA U471 ( .A(n204), .Z(n215) );
  ND2P U472 ( .A(n256), .B(n257), .Z(n226) );
  ND4P U473 ( .A(n263), .B(n270), .C(n271), .D(n272), .Z(n205) );
  ND2P U474 ( .A(n273), .B(n274), .Z(n225) );
  IVA U475 ( .A(n268), .Z(n277) );
  OR2 U476 ( .A(n294), .B(n142), .Z(n286) );
  IVA U477 ( .A(n272), .Z(n294) );
  IVA U478 ( .A(n293), .Z(n298) );
  ND2P U479 ( .A(n302), .B(n303), .Z(n214) );
  ND2P U480 ( .A(n306), .B(n307), .Z(n249) );
  AO7P U481 ( .A(n308), .B(n309), .C(n310), .Z(n307) );
  ND4P U482 ( .A(n5), .B(n302), .C(n45), .D(n312), .Z(n142) );
  ND2 U483 ( .A(n323), .B(n306), .Z(n322) );
  AN2P U484 ( .A(n312), .B(n304), .Z(n325) );
  ND2P U485 ( .A(B[68]), .B(A[68]), .Z(n304) );
  ND4P U486 ( .A(n333), .B(n334), .C(n335), .D(n336), .Z(n209) );
  IVA U487 ( .A(n232), .Z(n341) );
  IVA U488 ( .A(n223), .Z(n351) );
  ND3P U489 ( .A(n327), .B(n48), .C(n328), .Z(n224) );
  ND2P U490 ( .A(n362), .B(n369), .Z(n235) );
  IVA U491 ( .A(n378), .Z(n311) );
  AO7P U492 ( .A(n379), .B(n380), .C(n3), .Z(n378) );
  IVA U493 ( .A(n357), .Z(n391) );
  ND2P U494 ( .A(B[62]), .B(A[62]), .Z(n356) );
  ND2 U495 ( .A(n393), .B(n360), .Z(n392) );
  AO7P U496 ( .A(n42), .B(n394), .C(n381), .Z(n393) );
  NR2P U497 ( .A(n395), .B(n396), .Z(n394) );
  AO6P U498 ( .A(n400), .B(n401), .C(n35), .Z(n395) );
  ND4P U499 ( .A(n389), .B(n17), .C(n402), .D(n403), .Z(n368) );
  ND2 U500 ( .A(n414), .B(n44), .Z(n413) );
  ND2P U501 ( .A(B[56]), .B(A[56]), .Z(n386) );
  IVA U502 ( .A(n418), .Z(n400) );
  IVA U503 ( .A(n370), .Z(n423) );
  ND4P U504 ( .A(n421), .B(n426), .C(n375), .D(n427), .Z(n365) );
  ND2P U505 ( .A(B[54]), .B(A[54]), .Z(n422) );
  AO7P U506 ( .A(n437), .B(n438), .C(n424), .Z(n435) );
  IVA U507 ( .A(n439), .Z(n438) );
  ND2P U508 ( .A(n441), .B(n442), .Z(n439) );
  OR2 U509 ( .A(n473), .B(n31), .Z(n442) );
  IVA U510 ( .A(n454), .Z(n449) );
  AN2P U511 ( .A(n455), .B(n456), .Z(n447) );
  ND2P U512 ( .A(n459), .B(n460), .Z(n428) );
  ND2 U513 ( .A(n455), .B(n461), .Z(n457) );
  ND2P U514 ( .A(B[47]), .B(A[47]), .Z(n473) );
endmodule


module LOG_POLY_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [47:0] A;
  input [47:0] B;
  output [95:0] PRODUCT;
  input TC;
  wire   \ab[47][47] , \ab[47][45] , \ab[47][44] , \ab[47][43] , \ab[47][42] ,
         \ab[47][41] , \ab[47][40] , \ab[47][39] , \ab[47][38] , \ab[47][37] ,
         \ab[47][36] , \ab[47][35] , \ab[47][34] , \ab[47][33] , \ab[47][32] ,
         \ab[47][31] , \ab[47][30] , \ab[47][29] , \ab[47][28] , \ab[47][27] ,
         \ab[47][26] , \ab[47][25] , \ab[47][24] , \ab[47][23] , \ab[47][22] ,
         \ab[47][21] , \ab[47][20] , \ab[47][19] , \ab[47][18] , \ab[47][17] ,
         \ab[47][16] , \ab[47][15] , \ab[47][14] , \ab[47][13] , \ab[47][12] ,
         \ab[47][11] , \ab[47][10] , \ab[46][46] , \ab[46][45] , \ab[46][44] ,
         \ab[46][43] , \ab[46][42] , \ab[46][41] , \ab[46][40] , \ab[46][39] ,
         \ab[46][38] , \ab[46][37] , \ab[46][36] , \ab[46][35] , \ab[46][34] ,
         \ab[46][33] , \ab[46][32] , \ab[46][31] , \ab[46][30] , \ab[46][29] ,
         \ab[46][28] , \ab[46][27] , \ab[46][26] , \ab[46][25] , \ab[46][24] ,
         \ab[46][23] , \ab[46][22] , \ab[46][21] , \ab[46][20] , \ab[46][19] ,
         \ab[46][18] , \ab[46][17] , \ab[46][16] , \ab[46][15] , \ab[46][14] ,
         \ab[46][13] , \ab[46][12] , \ab[46][11] , \ab[46][10] , \ab[45][45] ,
         \ab[45][44] , \ab[45][43] , \ab[45][42] , \ab[45][41] , \ab[45][40] ,
         \ab[45][39] , \ab[45][38] , \ab[45][37] , \ab[45][36] , \ab[45][35] ,
         \ab[45][34] , \ab[45][33] , \ab[45][32] , \ab[45][31] , \ab[45][30] ,
         \ab[45][29] , \ab[45][28] , \ab[45][27] , \ab[45][26] , \ab[45][25] ,
         \ab[45][24] , \ab[45][23] , \ab[45][22] , \ab[45][21] , \ab[45][20] ,
         \ab[45][19] , \ab[45][18] , \ab[45][17] , \ab[45][16] , \ab[45][15] ,
         \ab[45][14] , \ab[45][13] , \ab[45][12] , \ab[45][11] , \ab[45][10] ,
         \ab[44][44] , \ab[44][43] , \ab[44][42] , \ab[44][41] , \ab[44][40] ,
         \ab[44][39] , \ab[44][38] , \ab[44][37] , \ab[44][36] , \ab[44][35] ,
         \ab[44][34] , \ab[44][33] , \ab[44][32] , \ab[44][31] , \ab[44][30] ,
         \ab[44][29] , \ab[44][28] , \ab[44][27] , \ab[44][26] , \ab[44][25] ,
         \ab[44][24] , \ab[44][23] , \ab[44][22] , \ab[44][21] , \ab[44][20] ,
         \ab[44][19] , \ab[44][18] , \ab[44][17] , \ab[44][16] , \ab[44][15] ,
         \ab[44][14] , \ab[44][13] , \ab[44][12] , \ab[44][11] , \ab[44][10] ,
         \ab[43][43] , \ab[43][42] , \ab[43][41] , \ab[43][40] , \ab[43][39] ,
         \ab[43][38] , \ab[43][37] , \ab[43][36] , \ab[43][35] , \ab[43][34] ,
         \ab[43][33] , \ab[43][32] , \ab[43][31] , \ab[43][30] , \ab[43][29] ,
         \ab[43][28] , \ab[43][27] , \ab[43][26] , \ab[43][25] , \ab[43][24] ,
         \ab[43][23] , \ab[43][22] , \ab[43][21] , \ab[43][20] , \ab[43][19] ,
         \ab[43][18] , \ab[43][17] , \ab[43][16] , \ab[43][15] , \ab[43][14] ,
         \ab[43][13] , \ab[43][12] , \ab[43][11] , \ab[43][10] , \ab[42][42] ,
         \ab[42][41] , \ab[42][40] , \ab[42][39] , \ab[42][38] , \ab[42][37] ,
         \ab[42][36] , \ab[42][35] , \ab[42][34] , \ab[42][33] , \ab[42][32] ,
         \ab[42][31] , \ab[42][30] , \ab[42][29] , \ab[42][28] , \ab[42][27] ,
         \ab[42][26] , \ab[42][25] , \ab[42][24] , \ab[42][23] , \ab[42][22] ,
         \ab[42][21] , \ab[42][20] , \ab[42][19] , \ab[42][18] , \ab[42][17] ,
         \ab[42][16] , \ab[42][15] , \ab[42][14] , \ab[42][13] , \ab[42][12] ,
         \ab[42][11] , \ab[42][10] , \ab[41][41] , \ab[41][40] , \ab[41][39] ,
         \ab[41][38] , \ab[41][37] , \ab[41][36] , \ab[41][35] , \ab[41][34] ,
         \ab[41][33] , \ab[41][32] , \ab[41][31] , \ab[41][30] , \ab[41][29] ,
         \ab[41][28] , \ab[41][27] , \ab[41][26] , \ab[41][25] , \ab[41][24] ,
         \ab[41][23] , \ab[41][22] , \ab[41][21] , \ab[41][20] , \ab[41][19] ,
         \ab[41][18] , \ab[41][17] , \ab[41][16] , \ab[41][15] , \ab[41][14] ,
         \ab[41][13] , \ab[41][12] , \ab[41][11] , \ab[41][10] , \ab[40][40] ,
         \ab[40][39] , \ab[40][38] , \ab[40][37] , \ab[40][36] , \ab[40][35] ,
         \ab[40][34] , \ab[40][33] , \ab[40][32] , \ab[40][31] , \ab[40][30] ,
         \ab[40][29] , \ab[40][28] , \ab[40][27] , \ab[40][26] , \ab[40][25] ,
         \ab[40][24] , \ab[40][23] , \ab[40][22] , \ab[40][21] , \ab[40][20] ,
         \ab[40][19] , \ab[40][18] , \ab[40][17] , \ab[40][16] , \ab[40][15] ,
         \ab[40][14] , \ab[40][13] , \ab[40][12] , \ab[40][11] , \ab[39][39] ,
         \ab[39][38] , \ab[39][37] , \ab[39][36] , \ab[39][35] , \ab[39][34] ,
         \ab[39][33] , \ab[39][32] , \ab[39][31] , \ab[39][30] , \ab[39][29] ,
         \ab[39][28] , \ab[39][27] , \ab[39][26] , \ab[39][25] , \ab[39][24] ,
         \ab[39][23] , \ab[39][22] , \ab[39][21] , \ab[39][20] , \ab[39][19] ,
         \ab[39][18] , \ab[39][17] , \ab[39][16] , \ab[39][15] , \ab[39][14] ,
         \ab[39][13] , \ab[39][12] , \ab[39][11] , \ab[38][38] , \ab[38][37] ,
         \ab[38][36] , \ab[38][35] , \ab[38][34] , \ab[38][33] , \ab[38][32] ,
         \ab[38][31] , \ab[38][30] , \ab[38][29] , \ab[38][28] , \ab[38][27] ,
         \ab[38][26] , \ab[38][25] , \ab[38][24] , \ab[38][23] , \ab[38][22] ,
         \ab[38][21] , \ab[38][20] , \ab[38][19] , \ab[38][18] , \ab[38][17] ,
         \ab[38][16] , \ab[38][15] , \ab[38][14] , \ab[38][13] , \ab[38][12] ,
         \ab[38][11] , \ab[37][37] , \ab[37][36] , \ab[37][35] , \ab[37][34] ,
         \ab[37][33] , \ab[37][32] , \ab[37][31] , \ab[37][30] , \ab[37][29] ,
         \ab[37][28] , \ab[37][27] , \ab[37][26] , \ab[37][25] , \ab[37][24] ,
         \ab[37][23] , \ab[37][22] , \ab[37][21] , \ab[37][20] , \ab[37][19] ,
         \ab[37][18] , \ab[37][17] , \ab[37][16] , \ab[37][15] , \ab[37][14] ,
         \ab[37][13] , \ab[37][12] , \ab[36][36] , \ab[36][35] , \ab[36][34] ,
         \ab[36][33] , \ab[36][32] , \ab[36][31] , \ab[36][30] , \ab[36][29] ,
         \ab[36][28] , \ab[36][27] , \ab[36][26] , \ab[36][25] , \ab[36][24] ,
         \ab[36][23] , \ab[36][22] , \ab[36][21] , \ab[36][20] , \ab[36][19] ,
         \ab[36][18] , \ab[36][17] , \ab[36][16] , \ab[36][15] , \ab[36][14] ,
         \ab[36][13] , \ab[36][12] , \ab[35][35] , \ab[35][34] , \ab[35][33] ,
         \ab[35][32] , \ab[35][31] , \ab[35][30] , \ab[35][29] , \ab[35][28] ,
         \ab[35][27] , \ab[35][26] , \ab[35][25] , \ab[35][24] , \ab[35][23] ,
         \ab[35][22] , \ab[35][21] , \ab[35][20] , \ab[35][19] , \ab[35][18] ,
         \ab[35][17] , \ab[35][16] , \ab[35][15] , \ab[35][14] , \ab[35][13] ,
         \ab[34][34] , \ab[34][33] , \ab[34][32] , \ab[34][31] , \ab[34][30] ,
         \ab[34][29] , \ab[34][28] , \ab[34][27] , \ab[34][26] , \ab[34][25] ,
         \ab[34][24] , \ab[34][23] , \ab[34][22] , \ab[34][21] , \ab[34][20] ,
         \ab[34][19] , \ab[34][18] , \ab[34][17] , \ab[34][16] , \ab[34][15] ,
         \ab[34][14] , \ab[34][13] , \ab[33][33] , \ab[33][32] , \ab[33][31] ,
         \ab[33][30] , \ab[33][29] , \ab[33][28] , \ab[33][27] , \ab[33][26] ,
         \ab[33][25] , \ab[33][24] , \ab[33][23] , \ab[33][22] , \ab[33][21] ,
         \ab[33][20] , \ab[33][19] , \ab[33][18] , \ab[33][17] , \ab[33][16] ,
         \ab[33][15] , \ab[33][14] , \ab[33][13] , \ab[32][32] , \ab[32][31] ,
         \ab[32][30] , \ab[32][29] , \ab[32][28] , \ab[32][27] , \ab[32][26] ,
         \ab[32][25] , \ab[32][24] , \ab[32][23] , \ab[32][22] , \ab[32][21] ,
         \ab[32][20] , \ab[32][19] , \ab[32][18] , \ab[32][17] , \ab[32][16] ,
         \ab[32][15] , \ab[32][14] , \ab[31][31] , \ab[31][30] , \ab[31][29] ,
         \ab[31][28] , \ab[31][27] , \ab[31][26] , \ab[31][25] , \ab[31][24] ,
         \ab[31][23] , \ab[31][22] , \ab[31][21] , \ab[31][20] , \ab[31][19] ,
         \ab[31][18] , \ab[31][17] , \ab[31][16] , \ab[31][15] , \ab[31][14] ,
         \ab[30][30] , \ab[30][29] , \ab[30][28] , \ab[30][27] , \ab[30][26] ,
         \ab[30][25] , \ab[30][24] , \ab[30][23] , \ab[30][22] , \ab[30][21] ,
         \ab[30][20] , \ab[30][19] , \ab[30][18] , \ab[30][17] , \ab[30][16] ,
         \ab[30][15] , \ab[29][29] , \ab[29][28] , \ab[29][27] , \ab[29][26] ,
         \ab[29][25] , \ab[29][24] , \ab[29][23] , \ab[29][22] , \ab[29][21] ,
         \ab[29][20] , \ab[29][19] , \ab[29][18] , \ab[29][17] , \ab[29][16] ,
         \ab[28][28] , \ab[28][27] , \ab[28][26] , \ab[28][25] , \ab[28][24] ,
         \ab[28][23] , \ab[28][22] , \ab[28][21] , \ab[28][20] , \ab[28][19] ,
         \ab[28][18] , \ab[28][17] , \ab[28][16] , \ab[27][27] , \ab[27][26] ,
         \ab[27][25] , \ab[27][24] , \ab[27][23] , \ab[27][22] , \ab[27][21] ,
         \ab[27][20] , \ab[27][19] , \ab[27][18] , \ab[27][17] , \ab[27][16] ,
         \ab[26][26] , \ab[26][25] , \ab[26][24] , \ab[26][23] , \ab[26][22] ,
         \ab[26][21] , \ab[26][20] , \ab[26][19] , \ab[26][18] , \ab[26][17] ,
         \ab[26][16] , \ab[25][25] , \ab[25][24] , \ab[25][23] , \ab[25][22] ,
         \ab[25][21] , \ab[25][20] , \ab[25][19] , \ab[25][18] , \ab[25][17] ,
         \ab[25][16] , \ab[24][24] , \ab[24][23] , \ab[24][22] , \ab[24][21] ,
         \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] , \ab[24][16] ,
         \ab[23][23] , \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] ,
         \ab[23][18] , \ab[23][17] , \ab[23][16] , \ab[22][22] , \ab[22][21] ,
         \ab[22][20] , \ab[22][19] , \ab[22][18] , \ab[22][17] , \ab[22][16] ,
         \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] ,
         \ab[21][16] , \ab[20][20] , \ab[20][19] , \ab[20][18] , \ab[20][17] ,
         \ab[20][16] , \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] ,
         \ab[18][18] , \ab[18][17] , \ab[18][16] , \ab[17][17] , \ab[17][16] ,
         \ab[16][16] , \ab[15][15] , \ab[14][14] , \ab[13][13] , \ab[12][12] ,
         \ab[11][11] , \ab[10][10] , \ab[9][47] , \ab[9][46] , \ab[9][45] ,
         \ab[9][44] , \ab[9][9] , \ab[8][47] , \ab[8][8] , \ab[7][47] ,
         \ab[7][7] , \ab[6][6] , \ab[5][5] , \ab[4][4] , \ab[3][3] ,
         \ab[2][2] , \ab[1][1] , \ab[1][0] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][46] , \CARRYB[4][45] ,
         \CARRYB[4][44] , \CARRYB[4][43] , \CARRYB[4][42] , \CARRYB[4][41] ,
         \CARRYB[4][40] , \CARRYB[4][39] , \CARRYB[4][38] , \CARRYB[4][37] ,
         \CARRYB[4][36] , \CARRYB[4][35] , \CARRYB[4][34] , \CARRYB[4][33] ,
         \CARRYB[4][32] , \CARRYB[4][31] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][46] , \CARRYB[3][45] , \CARRYB[3][44] ,
         \CARRYB[3][43] , \CARRYB[3][42] , \CARRYB[3][41] , \CARRYB[3][40] ,
         \CARRYB[3][39] , \CARRYB[3][38] , \CARRYB[3][37] , \CARRYB[3][36] ,
         \CARRYB[3][35] , \CARRYB[3][34] , \CARRYB[3][33] , \CARRYB[3][32] ,
         \CARRYB[3][31] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][46] , \CARRYB[2][45] , \CARRYB[2][44] , \CARRYB[2][43] ,
         \CARRYB[2][42] , \CARRYB[2][41] , \CARRYB[2][40] , \CARRYB[2][39] ,
         \CARRYB[2][38] , \CARRYB[2][37] , \CARRYB[2][36] , \CARRYB[2][35] ,
         \CARRYB[2][34] , \CARRYB[2][33] , \CARRYB[2][32] , \CARRYB[2][31] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][46] ,
         \CARRYB[1][45] , \CARRYB[1][43] , \CARRYB[1][42] , \CARRYB[1][41] ,
         \CARRYB[1][40] , \CARRYB[1][39] , \CARRYB[1][38] , \CARRYB[1][37] ,
         \CARRYB[1][36] , \CARRYB[1][35] , \CARRYB[1][34] , \CARRYB[1][33] ,
         \CARRYB[1][32] , \CARRYB[1][31] , \CARRYB[1][30] , \CARRYB[1][29] ,
         \CARRYB[1][28] , \CARRYB[1][27] , \CARRYB[1][26] , \CARRYB[1][25] ,
         \CARRYB[1][24] , \CARRYB[1][23] , \CARRYB[1][22] , \CARRYB[1][21] ,
         \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] , \CARRYB[1][17] ,
         \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][46] , \SUMB[4][45] ,
         \SUMB[4][44] , \SUMB[4][43] , \SUMB[4][42] , \SUMB[4][41] ,
         \SUMB[4][40] , \SUMB[4][39] , \SUMB[4][38] , \SUMB[4][37] ,
         \SUMB[4][36] , \SUMB[4][35] , \SUMB[4][34] , \SUMB[4][33] ,
         \SUMB[4][32] , \SUMB[4][31] , \SUMB[4][30] , \SUMB[4][29] ,
         \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] , \SUMB[4][25] ,
         \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] , \SUMB[4][21] ,
         \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] , \SUMB[4][17] ,
         \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] ,
         \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] ,
         \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][46] ,
         \SUMB[3][45] , \SUMB[3][44] , \SUMB[3][43] , \SUMB[3][42] ,
         \SUMB[3][41] , \SUMB[3][40] , \SUMB[3][39] , \SUMB[3][38] ,
         \SUMB[3][37] , \SUMB[3][36] , \SUMB[3][35] , \SUMB[3][34] ,
         \SUMB[3][33] , \SUMB[3][32] , \SUMB[3][31] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][46] ,
         \SUMB[2][45] , \SUMB[2][44] , \SUMB[2][43] , \SUMB[2][42] ,
         \SUMB[2][41] , \SUMB[2][40] , \SUMB[2][39] , \SUMB[2][38] ,
         \SUMB[2][37] , \SUMB[2][36] , \SUMB[2][35] , \SUMB[2][34] ,
         \SUMB[2][33] , \SUMB[2][32] , \SUMB[2][31] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][46] ,
         \SUMB[1][45] , \SUMB[1][44] , \SUMB[1][43] , \SUMB[1][42] ,
         \SUMB[1][41] , \SUMB[1][40] , \SUMB[1][39] , \SUMB[1][38] ,
         \SUMB[1][37] , \SUMB[1][36] , \SUMB[1][35] , \SUMB[1][34] ,
         \SUMB[1][33] , \SUMB[1][32] , \SUMB[1][31] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[15][46] , \CARRYB[15][45] , \CARRYB[15][44] ,
         \CARRYB[15][43] , \CARRYB[15][42] , \CARRYB[15][41] ,
         \CARRYB[15][40] , \CARRYB[15][39] , \CARRYB[15][38] ,
         \CARRYB[15][37] , \CARRYB[15][36] , \CARRYB[15][35] ,
         \CARRYB[15][34] , \CARRYB[15][33] , \CARRYB[15][32] ,
         \CARRYB[15][31] , \CARRYB[15][30] , \CARRYB[15][29] ,
         \CARRYB[15][28] , \CARRYB[15][27] , \CARRYB[15][26] ,
         \CARRYB[15][25] , \CARRYB[15][24] , \CARRYB[15][23] ,
         \CARRYB[15][22] , \CARRYB[15][21] , \CARRYB[15][20] ,
         \CARRYB[15][19] , \CARRYB[15][18] , \CARRYB[15][17] ,
         \CARRYB[15][16] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][46] ,
         \CARRYB[14][45] , \CARRYB[14][44] , \CARRYB[14][43] ,
         \CARRYB[14][42] , \CARRYB[14][41] , \CARRYB[14][40] ,
         \CARRYB[14][39] , \CARRYB[14][38] , \CARRYB[14][37] ,
         \CARRYB[14][36] , \CARRYB[14][35] , \CARRYB[14][34] ,
         \CARRYB[14][33] , \CARRYB[14][32] , \CARRYB[14][31] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][46] , \CARRYB[13][45] , \CARRYB[13][44] ,
         \CARRYB[13][43] , \CARRYB[13][42] , \CARRYB[13][41] ,
         \CARRYB[13][40] , \CARRYB[13][39] , \CARRYB[13][38] ,
         \CARRYB[13][37] , \CARRYB[13][36] , \CARRYB[13][35] ,
         \CARRYB[13][34] , \CARRYB[13][33] , \CARRYB[13][32] ,
         \CARRYB[13][31] , \CARRYB[13][30] , \CARRYB[13][29] ,
         \CARRYB[13][28] , \CARRYB[13][27] , \CARRYB[13][26] ,
         \CARRYB[13][25] , \CARRYB[13][24] , \CARRYB[13][23] ,
         \CARRYB[13][22] , \CARRYB[13][21] , \CARRYB[13][20] ,
         \CARRYB[13][19] , \CARRYB[13][18] , \CARRYB[13][17] ,
         \CARRYB[13][16] , \CARRYB[13][15] , \CARRYB[13][14] ,
         \CARRYB[13][13] , \CARRYB[13][12] , \CARRYB[13][11] ,
         \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] , \CARRYB[13][7] ,
         \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] , \CARRYB[13][3] ,
         \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] , \CARRYB[12][46] ,
         \CARRYB[12][45] , \CARRYB[12][44] , \CARRYB[12][43] ,
         \CARRYB[12][42] , \CARRYB[12][41] , \CARRYB[12][40] ,
         \CARRYB[12][39] , \CARRYB[12][38] , \CARRYB[12][37] ,
         \CARRYB[12][36] , \CARRYB[12][35] , \CARRYB[12][34] ,
         \CARRYB[12][33] , \CARRYB[12][32] , \CARRYB[12][31] ,
         \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][46] , \CARRYB[11][45] , \CARRYB[11][44] ,
         \CARRYB[11][43] , \CARRYB[11][42] , \CARRYB[11][41] ,
         \CARRYB[11][40] , \CARRYB[11][39] , \CARRYB[11][38] ,
         \CARRYB[11][37] , \CARRYB[11][36] , \CARRYB[11][35] ,
         \CARRYB[11][34] , \CARRYB[11][33] , \CARRYB[11][32] ,
         \CARRYB[11][31] , \CARRYB[11][30] , \CARRYB[11][29] ,
         \CARRYB[11][28] , \CARRYB[11][27] , \CARRYB[11][26] ,
         \CARRYB[11][25] , \CARRYB[11][24] , \CARRYB[11][23] ,
         \CARRYB[11][22] , \CARRYB[11][21] , \CARRYB[11][20] ,
         \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \CARRYB[11][15] , \CARRYB[11][14] ,
         \CARRYB[11][13] , \CARRYB[11][12] , \CARRYB[11][11] ,
         \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] , \CARRYB[11][7] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][46] ,
         \CARRYB[10][45] , \CARRYB[10][44] , \CARRYB[10][43] ,
         \CARRYB[10][42] , \CARRYB[10][41] , \CARRYB[10][40] ,
         \CARRYB[10][39] , \CARRYB[10][38] , \CARRYB[10][37] ,
         \CARRYB[10][36] , \CARRYB[10][35] , \CARRYB[10][34] ,
         \CARRYB[10][33] , \CARRYB[10][32] , \CARRYB[10][31] ,
         \CARRYB[10][30] , \CARRYB[10][29] , \CARRYB[10][28] ,
         \CARRYB[10][27] , \CARRYB[10][26] , \CARRYB[10][25] ,
         \CARRYB[10][24] , \CARRYB[10][23] , \CARRYB[10][22] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][46] , \CARRYB[9][45] , \CARRYB[9][44] ,
         \CARRYB[9][43] , \CARRYB[9][42] , \CARRYB[9][41] , \CARRYB[9][40] ,
         \CARRYB[9][39] , \CARRYB[9][38] , \CARRYB[9][37] , \CARRYB[9][36] ,
         \CARRYB[9][35] , \CARRYB[9][34] , \CARRYB[9][33] , \CARRYB[9][32] ,
         \CARRYB[9][31] , \CARRYB[9][30] , \CARRYB[9][29] , \CARRYB[9][28] ,
         \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][25] , \CARRYB[9][24] ,
         \CARRYB[9][23] , \CARRYB[9][22] , \CARRYB[9][21] , \CARRYB[9][20] ,
         \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] , \CARRYB[9][16] ,
         \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] ,
         \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] ,
         \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] ,
         \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] ,
         \CARRYB[8][46] , \CARRYB[8][45] , \CARRYB[8][44] , \CARRYB[8][43] ,
         \CARRYB[8][42] , \CARRYB[8][41] , \CARRYB[8][40] , \CARRYB[8][39] ,
         \CARRYB[8][38] , \CARRYB[8][37] , \CARRYB[8][36] , \CARRYB[8][35] ,
         \CARRYB[8][34] , \CARRYB[8][33] , \CARRYB[8][32] , \CARRYB[8][31] ,
         \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] , \CARRYB[8][27] ,
         \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] , \CARRYB[8][23] ,
         \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] , \CARRYB[8][19] ,
         \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] ,
         \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] ,
         \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] ,
         \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][46] ,
         \CARRYB[7][45] , \CARRYB[7][44] , \CARRYB[7][43] , \CARRYB[7][42] ,
         \CARRYB[7][41] , \CARRYB[7][40] , \CARRYB[7][39] , \CARRYB[7][38] ,
         \CARRYB[7][37] , \CARRYB[7][36] , \CARRYB[7][35] , \CARRYB[7][34] ,
         \CARRYB[7][33] , \CARRYB[7][32] , \CARRYB[7][31] , \CARRYB[7][30] ,
         \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] ,
         \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] ,
         \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] ,
         \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][46] , \CARRYB[6][45] ,
         \CARRYB[6][44] , \CARRYB[6][43] , \CARRYB[6][42] , \CARRYB[6][41] ,
         \CARRYB[6][40] , \CARRYB[6][39] , \CARRYB[6][38] , \CARRYB[6][37] ,
         \CARRYB[6][36] , \CARRYB[6][35] , \CARRYB[6][34] , \CARRYB[6][33] ,
         \CARRYB[6][32] , \CARRYB[6][31] , \CARRYB[6][30] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][46] , \CARRYB[5][45] , \CARRYB[5][44] ,
         \CARRYB[5][43] , \CARRYB[5][42] , \CARRYB[5][41] , \CARRYB[5][40] ,
         \CARRYB[5][39] , \CARRYB[5][38] , \CARRYB[5][37] , \CARRYB[5][36] ,
         \CARRYB[5][35] , \CARRYB[5][34] , \CARRYB[5][33] , \CARRYB[5][32] ,
         \CARRYB[5][31] , \CARRYB[5][30] , \CARRYB[5][29] , \CARRYB[5][28] ,
         \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] , \CARRYB[5][24] ,
         \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] , \CARRYB[5][20] ,
         \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] , \CARRYB[5][16] ,
         \SUMB[15][46] , \SUMB[15][45] , \SUMB[15][44] , \SUMB[15][43] ,
         \SUMB[15][42] , \SUMB[15][41] , \SUMB[15][40] , \SUMB[15][39] ,
         \SUMB[15][38] , \SUMB[15][37] , \SUMB[15][36] , \SUMB[15][35] ,
         \SUMB[15][34] , \SUMB[15][33] , \SUMB[15][32] , \SUMB[15][31] ,
         \SUMB[15][30] , \SUMB[15][29] , \SUMB[15][28] , \SUMB[15][27] ,
         \SUMB[15][26] , \SUMB[15][25] , \SUMB[15][24] , \SUMB[15][23] ,
         \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] , \SUMB[15][19] ,
         \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] , \SUMB[15][15] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][46] , \SUMB[14][45] ,
         \SUMB[14][44] , \SUMB[14][43] , \SUMB[14][42] , \SUMB[14][41] ,
         \SUMB[14][40] , \SUMB[14][39] , \SUMB[14][38] , \SUMB[14][37] ,
         \SUMB[14][36] , \SUMB[14][35] , \SUMB[14][34] , \SUMB[14][33] ,
         \SUMB[14][32] , \SUMB[14][31] , \SUMB[14][30] , \SUMB[14][29] ,
         \SUMB[14][28] , \SUMB[14][27] , \SUMB[14][26] , \SUMB[14][25] ,
         \SUMB[14][24] , \SUMB[14][23] , \SUMB[14][22] , \SUMB[14][21] ,
         \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] , \SUMB[14][17] ,
         \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][46] , \SUMB[13][45] , \SUMB[13][44] , \SUMB[13][43] ,
         \SUMB[13][42] , \SUMB[13][41] , \SUMB[13][40] , \SUMB[13][39] ,
         \SUMB[13][38] , \SUMB[13][37] , \SUMB[13][36] , \SUMB[13][35] ,
         \SUMB[13][34] , \SUMB[13][33] , \SUMB[13][32] , \SUMB[13][31] ,
         \SUMB[13][30] , \SUMB[13][29] , \SUMB[13][28] , \SUMB[13][27] ,
         \SUMB[13][26] , \SUMB[13][25] , \SUMB[13][24] , \SUMB[13][23] ,
         \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] , \SUMB[13][19] ,
         \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] , \SUMB[13][15] ,
         \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] ,
         \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][46] , \SUMB[12][45] ,
         \SUMB[12][44] , \SUMB[12][43] , \SUMB[12][42] , \SUMB[12][41] ,
         \SUMB[12][40] , \SUMB[12][39] , \SUMB[12][38] , \SUMB[12][37] ,
         \SUMB[12][36] , \SUMB[12][35] , \SUMB[12][34] , \SUMB[12][33] ,
         \SUMB[12][32] , \SUMB[12][31] , \SUMB[12][30] , \SUMB[12][29] ,
         \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] , \SUMB[12][25] ,
         \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] , \SUMB[12][21] ,
         \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] , \SUMB[12][17] ,
         \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] ,
         \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] ,
         \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][46] , \SUMB[11][45] , \SUMB[11][44] , \SUMB[11][43] ,
         \SUMB[11][42] , \SUMB[11][41] , \SUMB[11][40] , \SUMB[11][39] ,
         \SUMB[11][38] , \SUMB[11][37] , \SUMB[11][36] , \SUMB[11][35] ,
         \SUMB[11][34] , \SUMB[11][33] , \SUMB[11][32] , \SUMB[11][31] ,
         \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] , \SUMB[11][27] ,
         \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] , \SUMB[11][23] ,
         \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] , \SUMB[11][19] ,
         \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][46] , \SUMB[10][45] ,
         \SUMB[10][44] , \SUMB[10][43] , \SUMB[10][42] , \SUMB[10][41] ,
         \SUMB[10][40] , \SUMB[10][39] , \SUMB[10][38] , \SUMB[10][37] ,
         \SUMB[10][36] , \SUMB[10][35] , \SUMB[10][34] , \SUMB[10][33] ,
         \SUMB[10][32] , \SUMB[10][31] , \SUMB[10][30] , \SUMB[10][29] ,
         \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] , \SUMB[10][25] ,
         \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] , \SUMB[10][21] ,
         \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] ,
         \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][46] , \SUMB[9][45] , \SUMB[9][44] , \SUMB[9][43] ,
         \SUMB[9][42] , \SUMB[9][41] , \SUMB[9][40] , \SUMB[9][39] ,
         \SUMB[9][38] , \SUMB[9][37] , \SUMB[9][36] , \SUMB[9][35] ,
         \SUMB[9][34] , \SUMB[9][33] , \SUMB[9][32] , \SUMB[9][31] ,
         \SUMB[9][30] , \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] ,
         \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] ,
         \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] ,
         \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] ,
         \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] ,
         \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][46] , \SUMB[8][45] , \SUMB[8][44] , \SUMB[8][43] ,
         \SUMB[8][42] , \SUMB[8][41] , \SUMB[8][40] , \SUMB[8][39] ,
         \SUMB[8][38] , \SUMB[8][37] , \SUMB[8][36] , \SUMB[8][35] ,
         \SUMB[8][34] , \SUMB[8][33] , \SUMB[8][32] , \SUMB[8][31] ,
         \SUMB[8][30] , \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] ,
         \SUMB[8][26] , \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] ,
         \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][46] , \SUMB[7][45] , \SUMB[7][44] , \SUMB[7][43] ,
         \SUMB[7][42] , \SUMB[7][41] , \SUMB[7][40] , \SUMB[7][39] ,
         \SUMB[7][38] , \SUMB[7][37] , \SUMB[7][36] , \SUMB[7][35] ,
         \SUMB[7][34] , \SUMB[7][33] , \SUMB[7][32] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][46] , \SUMB[6][45] , \SUMB[6][44] , \SUMB[6][43] ,
         \SUMB[6][42] , \SUMB[6][41] , \SUMB[6][40] , \SUMB[6][39] ,
         \SUMB[6][38] , \SUMB[6][37] , \SUMB[6][36] , \SUMB[6][35] ,
         \SUMB[6][34] , \SUMB[6][33] , \SUMB[6][32] , \SUMB[6][31] ,
         \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] ,
         \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] ,
         \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] ,
         \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][46] , \SUMB[5][45] , \SUMB[5][44] , \SUMB[5][43] ,
         \SUMB[5][42] , \SUMB[5][41] , \SUMB[5][40] , \SUMB[5][39] ,
         \SUMB[5][38] , \SUMB[5][37] , \SUMB[5][36] , \SUMB[5][35] ,
         \SUMB[5][34] , \SUMB[5][33] , \SUMB[5][32] , \SUMB[5][31] ,
         \SUMB[5][30] , \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] ,
         \SUMB[5][26] , \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] ,
         \SUMB[5][22] , \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] ,
         \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] , \CARRYB[26][31] ,
         \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][46] , \CARRYB[25][45] , \CARRYB[25][44] ,
         \CARRYB[25][43] , \CARRYB[25][42] , \CARRYB[25][41] ,
         \CARRYB[25][40] , \CARRYB[25][39] , \CARRYB[25][38] ,
         \CARRYB[25][37] , \CARRYB[25][36] , \CARRYB[25][35] ,
         \CARRYB[25][34] , \CARRYB[25][33] , \CARRYB[25][32] ,
         \CARRYB[25][31] , \CARRYB[25][30] , \CARRYB[25][29] ,
         \CARRYB[25][28] , \CARRYB[25][27] , \CARRYB[25][26] ,
         \CARRYB[25][25] , \CARRYB[25][24] , \CARRYB[25][23] ,
         \CARRYB[25][22] , \CARRYB[25][21] , \CARRYB[25][20] ,
         \CARRYB[25][19] , \CARRYB[25][18] , \CARRYB[25][17] ,
         \CARRYB[25][16] , \CARRYB[25][15] , \CARRYB[25][14] ,
         \CARRYB[25][13] , \CARRYB[25][12] , \CARRYB[25][11] ,
         \CARRYB[25][10] , \CARRYB[25][9] , \CARRYB[25][8] , \CARRYB[25][7] ,
         \CARRYB[25][6] , \CARRYB[25][5] , \CARRYB[25][4] , \CARRYB[25][3] ,
         \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] , \CARRYB[24][46] ,
         \CARRYB[24][45] , \CARRYB[24][44] , \CARRYB[24][43] ,
         \CARRYB[24][42] , \CARRYB[24][41] , \CARRYB[24][40] ,
         \CARRYB[24][39] , \CARRYB[24][38] , \CARRYB[24][37] ,
         \CARRYB[24][36] , \CARRYB[24][35] , \CARRYB[24][34] ,
         \CARRYB[24][33] , \CARRYB[24][32] , \CARRYB[24][31] ,
         \CARRYB[24][30] , \CARRYB[24][29] , \CARRYB[24][28] ,
         \CARRYB[24][27] , \CARRYB[24][26] , \CARRYB[24][25] ,
         \CARRYB[24][24] , \CARRYB[24][23] , \CARRYB[24][22] ,
         \CARRYB[24][21] , \CARRYB[24][20] , \CARRYB[24][19] ,
         \CARRYB[24][18] , \CARRYB[24][17] , \CARRYB[24][16] ,
         \CARRYB[24][15] , \CARRYB[24][14] , \CARRYB[24][13] ,
         \CARRYB[24][12] , \CARRYB[24][11] , \CARRYB[24][10] , \CARRYB[24][9] ,
         \CARRYB[24][8] , \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] ,
         \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] ,
         \CARRYB[24][0] , \CARRYB[23][46] , \CARRYB[23][45] , \CARRYB[23][44] ,
         \CARRYB[23][43] , \CARRYB[23][42] , \CARRYB[23][41] ,
         \CARRYB[23][40] , \CARRYB[23][39] , \CARRYB[23][38] ,
         \CARRYB[23][37] , \CARRYB[23][36] , \CARRYB[23][35] ,
         \CARRYB[23][34] , \CARRYB[23][33] , \CARRYB[23][32] ,
         \CARRYB[23][31] , \CARRYB[23][30] , \CARRYB[23][29] ,
         \CARRYB[23][28] , \CARRYB[23][27] , \CARRYB[23][26] ,
         \CARRYB[23][25] , \CARRYB[23][24] , \CARRYB[23][23] ,
         \CARRYB[23][22] , \CARRYB[23][21] , \CARRYB[23][20] ,
         \CARRYB[23][19] , \CARRYB[23][18] , \CARRYB[23][17] ,
         \CARRYB[23][16] , \CARRYB[23][15] , \CARRYB[23][14] ,
         \CARRYB[23][13] , \CARRYB[23][12] , \CARRYB[23][11] ,
         \CARRYB[23][10] , \CARRYB[23][9] , \CARRYB[23][8] , \CARRYB[23][7] ,
         \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] ,
         \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][46] ,
         \CARRYB[22][45] , \CARRYB[22][44] , \CARRYB[22][43] ,
         \CARRYB[22][42] , \CARRYB[22][41] , \CARRYB[22][40] ,
         \CARRYB[22][39] , \CARRYB[22][38] , \CARRYB[22][37] ,
         \CARRYB[22][36] , \CARRYB[22][35] , \CARRYB[22][34] ,
         \CARRYB[22][33] , \CARRYB[22][32] , \CARRYB[22][31] ,
         \CARRYB[22][30] , \CARRYB[22][29] , \CARRYB[22][28] ,
         \CARRYB[22][27] , \CARRYB[22][26] , \CARRYB[22][25] ,
         \CARRYB[22][24] , \CARRYB[22][23] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][12] , \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] ,
         \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][46] , \CARRYB[21][45] , \CARRYB[21][44] ,
         \CARRYB[21][43] , \CARRYB[21][42] , \CARRYB[21][41] ,
         \CARRYB[21][40] , \CARRYB[21][39] , \CARRYB[21][38] ,
         \CARRYB[21][37] , \CARRYB[21][36] , \CARRYB[21][35] ,
         \CARRYB[21][34] , \CARRYB[21][33] , \CARRYB[21][32] ,
         \CARRYB[21][31] , \CARRYB[21][30] , \CARRYB[21][29] ,
         \CARRYB[21][28] , \CARRYB[21][27] , \CARRYB[21][26] ,
         \CARRYB[21][25] , \CARRYB[21][24] , \CARRYB[21][23] ,
         \CARRYB[21][22] , \CARRYB[21][21] , \CARRYB[21][20] ,
         \CARRYB[21][19] , \CARRYB[21][18] , \CARRYB[21][17] ,
         \CARRYB[21][16] , \CARRYB[21][15] , \CARRYB[21][14] ,
         \CARRYB[21][13] , \CARRYB[21][12] , \CARRYB[21][11] ,
         \CARRYB[21][10] , \CARRYB[21][9] , \CARRYB[21][8] , \CARRYB[21][7] ,
         \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] , \CARRYB[21][3] ,
         \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] , \CARRYB[20][46] ,
         \CARRYB[20][45] , \CARRYB[20][44] , \CARRYB[20][43] ,
         \CARRYB[20][42] , \CARRYB[20][41] , \CARRYB[20][40] ,
         \CARRYB[20][39] , \CARRYB[20][38] , \CARRYB[20][37] ,
         \CARRYB[20][36] , \CARRYB[20][35] , \CARRYB[20][34] ,
         \CARRYB[20][33] , \CARRYB[20][32] , \CARRYB[20][31] ,
         \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][46] , \CARRYB[19][45] , \CARRYB[19][44] ,
         \CARRYB[19][43] , \CARRYB[19][42] , \CARRYB[19][41] ,
         \CARRYB[19][40] , \CARRYB[19][39] , \CARRYB[19][38] ,
         \CARRYB[19][37] , \CARRYB[19][36] , \CARRYB[19][35] ,
         \CARRYB[19][34] , \CARRYB[19][33] , \CARRYB[19][32] ,
         \CARRYB[19][31] , \CARRYB[19][30] , \CARRYB[19][29] ,
         \CARRYB[19][28] , \CARRYB[19][27] , \CARRYB[19][26] ,
         \CARRYB[19][25] , \CARRYB[19][24] , \CARRYB[19][23] ,
         \CARRYB[19][22] , \CARRYB[19][21] , \CARRYB[19][20] ,
         \CARRYB[19][19] , \CARRYB[19][18] , \CARRYB[19][17] ,
         \CARRYB[19][16] , \CARRYB[19][15] , \CARRYB[19][14] ,
         \CARRYB[19][13] , \CARRYB[19][12] , \CARRYB[19][11] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][46] ,
         \CARRYB[18][45] , \CARRYB[18][44] , \CARRYB[18][43] ,
         \CARRYB[18][42] , \CARRYB[18][41] , \CARRYB[18][40] ,
         \CARRYB[18][39] , \CARRYB[18][38] , \CARRYB[18][37] ,
         \CARRYB[18][36] , \CARRYB[18][35] , \CARRYB[18][34] ,
         \CARRYB[18][33] , \CARRYB[18][32] , \CARRYB[18][31] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][46] , \CARRYB[17][45] , \CARRYB[17][44] ,
         \CARRYB[17][43] , \CARRYB[17][42] , \CARRYB[17][41] ,
         \CARRYB[17][40] , \CARRYB[17][39] , \CARRYB[17][38] ,
         \CARRYB[17][37] , \CARRYB[17][36] , \CARRYB[17][35] ,
         \CARRYB[17][34] , \CARRYB[17][33] , \CARRYB[17][32] ,
         \CARRYB[17][31] , \CARRYB[17][30] , \CARRYB[17][29] ,
         \CARRYB[17][28] , \CARRYB[17][27] , \CARRYB[17][26] ,
         \CARRYB[17][25] , \CARRYB[17][24] , \CARRYB[17][23] ,
         \CARRYB[17][22] , \CARRYB[17][21] , \CARRYB[17][20] ,
         \CARRYB[17][19] , \CARRYB[17][18] , \CARRYB[17][17] ,
         \CARRYB[17][16] , \CARRYB[17][15] , \CARRYB[17][14] ,
         \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][46] ,
         \CARRYB[16][45] , \CARRYB[16][44] , \CARRYB[16][43] ,
         \CARRYB[16][42] , \CARRYB[16][41] , \CARRYB[16][40] ,
         \CARRYB[16][39] , \CARRYB[16][38] , \CARRYB[16][37] ,
         \CARRYB[16][36] , \CARRYB[16][35] , \CARRYB[16][34] ,
         \CARRYB[16][33] , \CARRYB[16][32] , \CARRYB[16][31] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \SUMB[26][31] , \SUMB[26][30] , \SUMB[26][29] ,
         \SUMB[26][28] , \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] ,
         \SUMB[26][24] , \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] ,
         \SUMB[26][20] , \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] ,
         \SUMB[26][16] , \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] ,
         \SUMB[26][12] , \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] ,
         \SUMB[26][8] , \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] ,
         \SUMB[26][4] , \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] ,
         \SUMB[25][46] , \SUMB[25][45] , \SUMB[25][44] , \SUMB[25][43] ,
         \SUMB[25][42] , \SUMB[25][41] , \SUMB[25][40] , \SUMB[25][39] ,
         \SUMB[25][38] , \SUMB[25][37] , \SUMB[25][36] , \SUMB[25][35] ,
         \SUMB[25][34] , \SUMB[25][33] , \SUMB[25][32] , \SUMB[25][31] ,
         \SUMB[25][30] , \SUMB[25][29] , \SUMB[25][28] , \SUMB[25][27] ,
         \SUMB[25][26] , \SUMB[25][25] , \SUMB[25][24] , \SUMB[25][23] ,
         \SUMB[25][22] , \SUMB[25][21] , \SUMB[25][20] , \SUMB[25][19] ,
         \SUMB[25][18] , \SUMB[25][17] , \SUMB[25][16] , \SUMB[25][15] ,
         \SUMB[25][14] , \SUMB[25][13] , \SUMB[25][12] , \SUMB[25][11] ,
         \SUMB[25][10] , \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] ,
         \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] ,
         \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][46] , \SUMB[24][45] ,
         \SUMB[24][44] , \SUMB[24][43] , \SUMB[24][42] , \SUMB[24][41] ,
         \SUMB[24][40] , \SUMB[24][39] , \SUMB[24][38] , \SUMB[24][37] ,
         \SUMB[24][36] , \SUMB[24][35] , \SUMB[24][34] , \SUMB[24][33] ,
         \SUMB[24][32] , \SUMB[24][31] , \SUMB[24][30] , \SUMB[24][29] ,
         \SUMB[24][28] , \SUMB[24][27] , \SUMB[24][26] , \SUMB[24][25] ,
         \SUMB[24][24] , \SUMB[24][23] , \SUMB[24][22] , \SUMB[24][21] ,
         \SUMB[24][20] , \SUMB[24][19] , \SUMB[24][18] , \SUMB[24][17] ,
         \SUMB[24][16] , \SUMB[24][15] , \SUMB[24][14] , \SUMB[24][13] ,
         \SUMB[24][12] , \SUMB[24][11] , \SUMB[24][10] , \SUMB[24][9] ,
         \SUMB[24][8] , \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] ,
         \SUMB[24][4] , \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] ,
         \SUMB[23][46] , \SUMB[23][45] , \SUMB[23][44] , \SUMB[23][43] ,
         \SUMB[23][42] , \SUMB[23][41] , \SUMB[23][40] , \SUMB[23][39] ,
         \SUMB[23][38] , \SUMB[23][37] , \SUMB[23][36] , \SUMB[23][35] ,
         \SUMB[23][34] , \SUMB[23][33] , \SUMB[23][32] , \SUMB[23][31] ,
         \SUMB[23][30] , \SUMB[23][29] , \SUMB[23][28] , \SUMB[23][27] ,
         \SUMB[23][26] , \SUMB[23][25] , \SUMB[23][24] , \SUMB[23][23] ,
         \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] ,
         \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] ,
         \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] ,
         \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] ,
         \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] ,
         \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][46] , \SUMB[22][45] ,
         \SUMB[22][44] , \SUMB[22][43] , \SUMB[22][42] , \SUMB[22][41] ,
         \SUMB[22][40] , \SUMB[22][39] , \SUMB[22][38] , \SUMB[22][37] ,
         \SUMB[22][36] , \SUMB[22][35] , \SUMB[22][34] , \SUMB[22][33] ,
         \SUMB[22][32] , \SUMB[22][31] , \SUMB[22][30] , \SUMB[22][29] ,
         \SUMB[22][28] , \SUMB[22][27] , \SUMB[22][26] , \SUMB[22][25] ,
         \SUMB[22][24] , \SUMB[22][23] , \SUMB[22][22] , \SUMB[22][21] ,
         \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] ,
         \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][13] ,
         \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] , \SUMB[22][9] ,
         \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] ,
         \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] ,
         \SUMB[21][46] , \SUMB[21][45] , \SUMB[21][44] , \SUMB[21][43] ,
         \SUMB[21][42] , \SUMB[21][41] , \SUMB[21][40] , \SUMB[21][39] ,
         \SUMB[21][38] , \SUMB[21][37] , \SUMB[21][36] , \SUMB[21][35] ,
         \SUMB[21][34] , \SUMB[21][33] , \SUMB[21][32] , \SUMB[21][31] ,
         \SUMB[21][30] , \SUMB[21][29] , \SUMB[21][28] , \SUMB[21][27] ,
         \SUMB[21][26] , \SUMB[21][25] , \SUMB[21][24] , \SUMB[21][23] ,
         \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] , \SUMB[21][19] ,
         \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] , \SUMB[21][15] ,
         \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] , \SUMB[21][11] ,
         \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] ,
         \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] ,
         \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][46] , \SUMB[20][45] ,
         \SUMB[20][44] , \SUMB[20][43] , \SUMB[20][42] , \SUMB[20][41] ,
         \SUMB[20][40] , \SUMB[20][39] , \SUMB[20][38] , \SUMB[20][37] ,
         \SUMB[20][36] , \SUMB[20][35] , \SUMB[20][34] , \SUMB[20][33] ,
         \SUMB[20][32] , \SUMB[20][31] , \SUMB[20][30] , \SUMB[20][29] ,
         \SUMB[20][28] , \SUMB[20][27] , \SUMB[20][26] , \SUMB[20][25] ,
         \SUMB[20][24] , \SUMB[20][23] , \SUMB[20][22] , \SUMB[20][21] ,
         \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] ,
         \SUMB[20][16] , \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] ,
         \SUMB[20][12] , \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] ,
         \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] ,
         \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] ,
         \SUMB[19][46] , \SUMB[19][45] , \SUMB[19][44] , \SUMB[19][43] ,
         \SUMB[19][42] , \SUMB[19][41] , \SUMB[19][40] , \SUMB[19][39] ,
         \SUMB[19][38] , \SUMB[19][37] , \SUMB[19][36] , \SUMB[19][35] ,
         \SUMB[19][34] , \SUMB[19][33] , \SUMB[19][32] , \SUMB[19][31] ,
         \SUMB[19][30] , \SUMB[19][29] , \SUMB[19][28] , \SUMB[19][27] ,
         \SUMB[19][26] , \SUMB[19][25] , \SUMB[19][24] , \SUMB[19][23] ,
         \SUMB[19][22] , \SUMB[19][21] , \SUMB[19][20] , \SUMB[19][19] ,
         \SUMB[19][18] , \SUMB[19][17] , \SUMB[19][16] , \SUMB[19][15] ,
         \SUMB[19][14] , \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] ,
         \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][46] , \SUMB[18][45] ,
         \SUMB[18][44] , \SUMB[18][43] , \SUMB[18][42] , \SUMB[18][41] ,
         \SUMB[18][40] , \SUMB[18][39] , \SUMB[18][38] , \SUMB[18][37] ,
         \SUMB[18][36] , \SUMB[18][35] , \SUMB[18][34] , \SUMB[18][33] ,
         \SUMB[18][32] , \SUMB[18][31] , \SUMB[18][30] , \SUMB[18][29] ,
         \SUMB[18][28] , \SUMB[18][27] , \SUMB[18][26] , \SUMB[18][25] ,
         \SUMB[18][24] , \SUMB[18][23] , \SUMB[18][22] , \SUMB[18][21] ,
         \SUMB[18][20] , \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][17] ,
         \SUMB[18][16] , \SUMB[18][15] , \SUMB[18][14] , \SUMB[18][13] ,
         \SUMB[18][12] , \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] ,
         \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] ,
         \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] ,
         \SUMB[17][46] , \SUMB[17][45] , \SUMB[17][44] , \SUMB[17][43] ,
         \SUMB[17][42] , \SUMB[17][41] , \SUMB[17][40] , \SUMB[17][39] ,
         \SUMB[17][38] , \SUMB[17][37] , \SUMB[17][36] , \SUMB[17][35] ,
         \SUMB[17][34] , \SUMB[17][33] , \SUMB[17][32] , \SUMB[17][31] ,
         \SUMB[17][30] , \SUMB[17][29] , \SUMB[17][28] , \SUMB[17][27] ,
         \SUMB[17][26] , \SUMB[17][25] , \SUMB[17][24] , \SUMB[17][23] ,
         \SUMB[17][22] , \SUMB[17][21] , \SUMB[17][20] , \SUMB[17][19] ,
         \SUMB[17][18] , \SUMB[17][17] , \SUMB[17][16] , \SUMB[17][15] ,
         \SUMB[17][14] , \SUMB[17][13] , \SUMB[17][12] , \SUMB[17][11] ,
         \SUMB[17][10] , \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] ,
         \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] ,
         \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][46] , \SUMB[16][45] ,
         \SUMB[16][44] , \SUMB[16][43] , \SUMB[16][42] , \SUMB[16][41] ,
         \SUMB[16][40] , \SUMB[16][39] , \SUMB[16][38] , \SUMB[16][37] ,
         \SUMB[16][36] , \SUMB[16][35] , \SUMB[16][34] , \SUMB[16][33] ,
         \SUMB[16][32] , \SUMB[16][31] , \SUMB[16][30] , \SUMB[16][29] ,
         \SUMB[16][28] , \SUMB[16][27] , \SUMB[16][26] , \SUMB[16][25] ,
         \SUMB[16][24] , \SUMB[16][23] , \SUMB[16][22] , \SUMB[16][21] ,
         \SUMB[16][20] , \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] ,
         \SUMB[16][16] , \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] ,
         \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] ,
         \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] ,
         \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] ,
         \CARRYB[37][15] , \CARRYB[37][14] , \CARRYB[37][13] ,
         \CARRYB[37][12] , \CARRYB[37][11] , \CARRYB[37][10] , \CARRYB[37][9] ,
         \CARRYB[37][8] , \CARRYB[37][7] , \CARRYB[37][6] , \CARRYB[37][5] ,
         \CARRYB[37][4] , \CARRYB[37][3] , \CARRYB[37][2] , \CARRYB[37][1] ,
         \CARRYB[37][0] , \CARRYB[36][46] , \CARRYB[36][45] , \CARRYB[36][44] ,
         \CARRYB[36][43] , \CARRYB[36][42] , \CARRYB[36][41] ,
         \CARRYB[36][40] , \CARRYB[36][39] , \CARRYB[36][38] ,
         \CARRYB[36][37] , \CARRYB[36][36] , \CARRYB[36][35] ,
         \CARRYB[36][34] , \CARRYB[36][33] , \CARRYB[36][32] ,
         \CARRYB[36][31] , \CARRYB[36][30] , \CARRYB[36][29] ,
         \CARRYB[36][28] , \CARRYB[36][27] , \CARRYB[36][26] ,
         \CARRYB[36][25] , \CARRYB[36][24] , \CARRYB[36][23] ,
         \CARRYB[36][22] , \CARRYB[36][21] , \CARRYB[36][20] ,
         \CARRYB[36][19] , \CARRYB[36][18] , \CARRYB[36][17] ,
         \CARRYB[36][16] , \CARRYB[36][15] , \CARRYB[36][14] ,
         \CARRYB[36][13] , \CARRYB[36][12] , \CARRYB[36][11] ,
         \CARRYB[36][10] , \CARRYB[36][9] , \CARRYB[36][8] , \CARRYB[36][7] ,
         \CARRYB[36][6] , \CARRYB[36][5] , \CARRYB[36][4] , \CARRYB[36][3] ,
         \CARRYB[36][2] , \CARRYB[36][1] , \CARRYB[36][0] , \CARRYB[35][46] ,
         \CARRYB[35][45] , \CARRYB[35][44] , \CARRYB[35][43] ,
         \CARRYB[35][42] , \CARRYB[35][41] , \CARRYB[35][40] ,
         \CARRYB[35][39] , \CARRYB[35][38] , \CARRYB[35][37] ,
         \CARRYB[35][36] , \CARRYB[35][35] , \CARRYB[35][34] ,
         \CARRYB[35][33] , \CARRYB[35][32] , \CARRYB[35][31] ,
         \CARRYB[35][30] , \CARRYB[35][29] , \CARRYB[35][28] ,
         \CARRYB[35][27] , \CARRYB[35][26] , \CARRYB[35][25] ,
         \CARRYB[35][24] , \CARRYB[35][23] , \CARRYB[35][22] ,
         \CARRYB[35][21] , \CARRYB[35][20] , \CARRYB[35][19] ,
         \CARRYB[35][18] , \CARRYB[35][17] , \CARRYB[35][16] ,
         \CARRYB[35][15] , \CARRYB[35][14] , \CARRYB[35][13] ,
         \CARRYB[35][12] , \CARRYB[35][11] , \CARRYB[35][10] , \CARRYB[35][9] ,
         \CARRYB[35][8] , \CARRYB[35][7] , \CARRYB[35][6] , \CARRYB[35][5] ,
         \CARRYB[35][4] , \CARRYB[35][3] , \CARRYB[35][2] , \CARRYB[35][1] ,
         \CARRYB[35][0] , \CARRYB[34][46] , \CARRYB[34][45] , \CARRYB[34][44] ,
         \CARRYB[34][43] , \CARRYB[34][42] , \CARRYB[34][41] ,
         \CARRYB[34][40] , \CARRYB[34][39] , \CARRYB[34][38] ,
         \CARRYB[34][37] , \CARRYB[34][36] , \CARRYB[34][35] ,
         \CARRYB[34][34] , \CARRYB[34][33] , \CARRYB[34][32] ,
         \CARRYB[34][31] , \CARRYB[34][30] , \CARRYB[34][29] ,
         \CARRYB[34][28] , \CARRYB[34][27] , \CARRYB[34][26] ,
         \CARRYB[34][25] , \CARRYB[34][24] , \CARRYB[34][23] ,
         \CARRYB[34][22] , \CARRYB[34][21] , \CARRYB[34][20] ,
         \CARRYB[34][19] , \CARRYB[34][18] , \CARRYB[34][17] ,
         \CARRYB[34][16] , \CARRYB[34][15] , \CARRYB[34][14] ,
         \CARRYB[34][13] , \CARRYB[34][12] , \CARRYB[34][11] ,
         \CARRYB[34][10] , \CARRYB[34][9] , \CARRYB[34][8] , \CARRYB[34][7] ,
         \CARRYB[34][6] , \CARRYB[34][5] , \CARRYB[34][4] , \CARRYB[34][3] ,
         \CARRYB[34][2] , \CARRYB[34][1] , \CARRYB[34][0] , \CARRYB[33][46] ,
         \CARRYB[33][45] , \CARRYB[33][44] , \CARRYB[33][43] ,
         \CARRYB[33][42] , \CARRYB[33][41] , \CARRYB[33][40] ,
         \CARRYB[33][39] , \CARRYB[33][38] , \CARRYB[33][37] ,
         \CARRYB[33][36] , \CARRYB[33][35] , \CARRYB[33][34] ,
         \CARRYB[33][33] , \CARRYB[33][32] , \CARRYB[33][31] ,
         \CARRYB[33][30] , \CARRYB[33][29] , \CARRYB[33][28] ,
         \CARRYB[33][27] , \CARRYB[33][26] , \CARRYB[33][25] ,
         \CARRYB[33][24] , \CARRYB[33][23] , \CARRYB[33][22] ,
         \CARRYB[33][21] , \CARRYB[33][20] , \CARRYB[33][19] ,
         \CARRYB[33][18] , \CARRYB[33][17] , \CARRYB[33][16] ,
         \CARRYB[33][15] , \CARRYB[33][14] , \CARRYB[33][13] ,
         \CARRYB[33][12] , \CARRYB[33][11] , \CARRYB[33][10] , \CARRYB[33][9] ,
         \CARRYB[33][8] , \CARRYB[33][7] , \CARRYB[33][6] , \CARRYB[33][5] ,
         \CARRYB[33][4] , \CARRYB[33][3] , \CARRYB[33][2] , \CARRYB[33][1] ,
         \CARRYB[33][0] , \CARRYB[32][46] , \CARRYB[32][45] , \CARRYB[32][44] ,
         \CARRYB[32][43] , \CARRYB[32][42] , \CARRYB[32][41] ,
         \CARRYB[32][40] , \CARRYB[32][39] , \CARRYB[32][38] ,
         \CARRYB[32][37] , \CARRYB[32][36] , \CARRYB[32][35] ,
         \CARRYB[32][34] , \CARRYB[32][33] , \CARRYB[32][32] ,
         \CARRYB[32][31] , \CARRYB[32][30] , \CARRYB[32][29] ,
         \CARRYB[32][28] , \CARRYB[32][27] , \CARRYB[32][26] ,
         \CARRYB[32][25] , \CARRYB[32][24] , \CARRYB[32][23] ,
         \CARRYB[32][22] , \CARRYB[32][21] , \CARRYB[32][20] ,
         \CARRYB[32][19] , \CARRYB[32][18] , \CARRYB[32][17] ,
         \CARRYB[32][16] , \CARRYB[32][15] , \CARRYB[32][14] ,
         \CARRYB[32][13] , \CARRYB[32][12] , \CARRYB[32][11] ,
         \CARRYB[32][10] , \CARRYB[32][9] , \CARRYB[32][8] , \CARRYB[32][7] ,
         \CARRYB[32][6] , \CARRYB[32][5] , \CARRYB[32][4] , \CARRYB[32][3] ,
         \CARRYB[32][2] , \CARRYB[32][1] , \CARRYB[32][0] , \CARRYB[31][46] ,
         \CARRYB[31][45] , \CARRYB[31][44] , \CARRYB[31][43] ,
         \CARRYB[31][42] , \CARRYB[31][41] , \CARRYB[31][40] ,
         \CARRYB[31][39] , \CARRYB[31][38] , \CARRYB[31][37] ,
         \CARRYB[31][36] , \CARRYB[31][35] , \CARRYB[31][34] ,
         \CARRYB[31][33] , \CARRYB[31][32] , \CARRYB[31][31] ,
         \CARRYB[31][30] , \CARRYB[31][29] , \CARRYB[31][28] ,
         \CARRYB[31][27] , \CARRYB[31][26] , \CARRYB[31][25] ,
         \CARRYB[31][24] , \CARRYB[31][23] , \CARRYB[31][22] ,
         \CARRYB[31][21] , \CARRYB[31][20] , \CARRYB[31][19] ,
         \CARRYB[31][18] , \CARRYB[31][17] , \CARRYB[31][16] ,
         \CARRYB[31][15] , \CARRYB[31][14] , \CARRYB[31][13] ,
         \CARRYB[31][12] , \CARRYB[31][11] , \CARRYB[31][10] , \CARRYB[31][9] ,
         \CARRYB[31][8] , \CARRYB[31][7] , \CARRYB[31][6] , \CARRYB[31][5] ,
         \CARRYB[31][4] , \CARRYB[31][3] , \CARRYB[31][2] , \CARRYB[31][1] ,
         \CARRYB[31][0] , \CARRYB[30][46] , \CARRYB[30][45] , \CARRYB[30][44] ,
         \CARRYB[30][43] , \CARRYB[30][42] , \CARRYB[30][41] ,
         \CARRYB[30][40] , \CARRYB[30][39] , \CARRYB[30][38] ,
         \CARRYB[30][37] , \CARRYB[30][36] , \CARRYB[30][35] ,
         \CARRYB[30][34] , \CARRYB[30][33] , \CARRYB[30][32] ,
         \CARRYB[30][31] , \CARRYB[30][30] , \CARRYB[30][29] ,
         \CARRYB[30][28] , \CARRYB[30][27] , \CARRYB[30][26] ,
         \CARRYB[30][25] , \CARRYB[30][24] , \CARRYB[30][23] ,
         \CARRYB[30][22] , \CARRYB[30][21] , \CARRYB[30][20] ,
         \CARRYB[30][19] , \CARRYB[30][18] , \CARRYB[30][17] ,
         \CARRYB[30][16] , \CARRYB[30][15] , \CARRYB[30][14] ,
         \CARRYB[30][13] , \CARRYB[30][12] , \CARRYB[30][11] ,
         \CARRYB[30][10] , \CARRYB[30][9] , \CARRYB[30][8] , \CARRYB[30][7] ,
         \CARRYB[30][6] , \CARRYB[30][5] , \CARRYB[30][4] , \CARRYB[30][3] ,
         \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] , \CARRYB[29][46] ,
         \CARRYB[29][45] , \CARRYB[29][44] , \CARRYB[29][43] ,
         \CARRYB[29][42] , \CARRYB[29][41] , \CARRYB[29][40] ,
         \CARRYB[29][39] , \CARRYB[29][38] , \CARRYB[29][37] ,
         \CARRYB[29][36] , \CARRYB[29][35] , \CARRYB[29][34] ,
         \CARRYB[29][33] , \CARRYB[29][32] , \CARRYB[29][31] ,
         \CARRYB[29][30] , \CARRYB[29][29] , \CARRYB[29][28] ,
         \CARRYB[29][27] , \CARRYB[29][26] , \CARRYB[29][25] ,
         \CARRYB[29][24] , \CARRYB[29][23] , \CARRYB[29][22] ,
         \CARRYB[29][21] , \CARRYB[29][20] , \CARRYB[29][19] ,
         \CARRYB[29][18] , \CARRYB[29][17] , \CARRYB[29][16] ,
         \CARRYB[29][15] , \CARRYB[29][14] , \CARRYB[29][13] ,
         \CARRYB[29][12] , \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] ,
         \CARRYB[29][4] , \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][46] , \CARRYB[28][45] , \CARRYB[28][44] ,
         \CARRYB[28][43] , \CARRYB[28][42] , \CARRYB[28][41] ,
         \CARRYB[28][40] , \CARRYB[28][39] , \CARRYB[28][38] ,
         \CARRYB[28][37] , \CARRYB[28][36] , \CARRYB[28][35] ,
         \CARRYB[28][34] , \CARRYB[28][33] , \CARRYB[28][32] ,
         \CARRYB[28][31] , \CARRYB[28][30] , \CARRYB[28][29] ,
         \CARRYB[28][28] , \CARRYB[28][27] , \CARRYB[28][26] ,
         \CARRYB[28][25] , \CARRYB[28][24] , \CARRYB[28][23] ,
         \CARRYB[28][22] , \CARRYB[28][21] , \CARRYB[28][20] ,
         \CARRYB[28][19] , \CARRYB[28][18] , \CARRYB[28][17] ,
         \CARRYB[28][16] , \CARRYB[28][15] , \CARRYB[28][14] ,
         \CARRYB[28][13] , \CARRYB[28][12] , \CARRYB[28][11] ,
         \CARRYB[28][10] , \CARRYB[28][9] , \CARRYB[28][8] , \CARRYB[28][7] ,
         \CARRYB[28][6] , \CARRYB[28][5] , \CARRYB[28][4] , \CARRYB[28][3] ,
         \CARRYB[28][2] , \CARRYB[28][1] , \CARRYB[28][0] , \CARRYB[27][46] ,
         \CARRYB[27][45] , \CARRYB[27][44] , \CARRYB[27][43] ,
         \CARRYB[27][42] , \CARRYB[27][41] , \CARRYB[27][40] ,
         \CARRYB[27][39] , \CARRYB[27][38] , \CARRYB[27][37] ,
         \CARRYB[27][36] , \CARRYB[27][35] , \CARRYB[27][34] ,
         \CARRYB[27][33] , \CARRYB[27][32] , \CARRYB[27][31] ,
         \CARRYB[27][30] , \CARRYB[27][29] , \CARRYB[27][28] ,
         \CARRYB[27][27] , \CARRYB[27][26] , \CARRYB[27][25] ,
         \CARRYB[27][24] , \CARRYB[27][23] , \CARRYB[27][22] ,
         \CARRYB[27][21] , \CARRYB[27][20] , \CARRYB[27][19] ,
         \CARRYB[27][18] , \CARRYB[27][17] , \CARRYB[27][16] ,
         \CARRYB[27][15] , \CARRYB[27][14] , \CARRYB[27][13] ,
         \CARRYB[27][12] , \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] ,
         \CARRYB[27][8] , \CARRYB[27][7] , \CARRYB[27][6] , \CARRYB[27][5] ,
         \CARRYB[27][4] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][46] , \CARRYB[26][45] , \CARRYB[26][44] ,
         \CARRYB[26][43] , \CARRYB[26][42] , \CARRYB[26][41] ,
         \CARRYB[26][40] , \CARRYB[26][39] , \CARRYB[26][38] ,
         \CARRYB[26][37] , \CARRYB[26][36] , \CARRYB[26][35] ,
         \CARRYB[26][34] , \CARRYB[26][33] , \CARRYB[26][32] , \SUMB[37][15] ,
         \SUMB[37][14] , \SUMB[37][13] , \SUMB[37][12] , \SUMB[37][11] ,
         \SUMB[37][10] , \SUMB[37][9] , \SUMB[37][8] , \SUMB[37][7] ,
         \SUMB[37][6] , \SUMB[37][5] , \SUMB[37][4] , \SUMB[37][3] ,
         \SUMB[37][2] , \SUMB[37][1] , \SUMB[36][46] , \SUMB[36][45] ,
         \SUMB[36][44] , \SUMB[36][43] , \SUMB[36][42] , \SUMB[36][41] ,
         \SUMB[36][40] , \SUMB[36][39] , \SUMB[36][38] , \SUMB[36][37] ,
         \SUMB[36][36] , \SUMB[36][35] , \SUMB[36][34] , \SUMB[36][33] ,
         \SUMB[36][32] , \SUMB[36][31] , \SUMB[36][30] , \SUMB[36][29] ,
         \SUMB[36][28] , \SUMB[36][27] , \SUMB[36][26] , \SUMB[36][25] ,
         \SUMB[36][24] , \SUMB[36][23] , \SUMB[36][22] , \SUMB[36][21] ,
         \SUMB[36][20] , \SUMB[36][19] , \SUMB[36][18] , \SUMB[36][17] ,
         \SUMB[36][16] , \SUMB[36][15] , \SUMB[36][14] , \SUMB[36][13] ,
         \SUMB[36][12] , \SUMB[36][11] , \SUMB[36][10] , \SUMB[36][9] ,
         \SUMB[36][8] , \SUMB[36][7] , \SUMB[36][6] , \SUMB[36][5] ,
         \SUMB[36][4] , \SUMB[36][3] , \SUMB[36][2] , \SUMB[36][1] ,
         \SUMB[35][46] , \SUMB[35][45] , \SUMB[35][44] , \SUMB[35][43] ,
         \SUMB[35][42] , \SUMB[35][41] , \SUMB[35][40] , \SUMB[35][39] ,
         \SUMB[35][38] , \SUMB[35][37] , \SUMB[35][36] , \SUMB[35][35] ,
         \SUMB[35][34] , \SUMB[35][33] , \SUMB[35][32] , \SUMB[35][31] ,
         \SUMB[35][30] , \SUMB[35][29] , \SUMB[35][28] , \SUMB[35][27] ,
         \SUMB[35][26] , \SUMB[35][25] , \SUMB[35][24] , \SUMB[35][23] ,
         \SUMB[35][22] , \SUMB[35][21] , \SUMB[35][20] , \SUMB[35][19] ,
         \SUMB[35][18] , \SUMB[35][17] , \SUMB[35][16] , \SUMB[35][15] ,
         \SUMB[35][14] , \SUMB[35][13] , \SUMB[35][12] , \SUMB[35][11] ,
         \SUMB[35][10] , \SUMB[35][9] , \SUMB[35][8] , \SUMB[35][7] ,
         \SUMB[35][6] , \SUMB[35][5] , \SUMB[35][4] , \SUMB[35][3] ,
         \SUMB[35][2] , \SUMB[35][1] , \SUMB[34][46] , \SUMB[34][45] ,
         \SUMB[34][44] , \SUMB[34][43] , \SUMB[34][42] , \SUMB[34][41] ,
         \SUMB[34][40] , \SUMB[34][39] , \SUMB[34][38] , \SUMB[34][37] ,
         \SUMB[34][36] , \SUMB[34][35] , \SUMB[34][34] , \SUMB[34][33] ,
         \SUMB[34][32] , \SUMB[34][31] , \SUMB[34][30] , \SUMB[34][29] ,
         \SUMB[34][28] , \SUMB[34][27] , \SUMB[34][26] , \SUMB[34][25] ,
         \SUMB[34][24] , \SUMB[34][23] , \SUMB[34][22] , \SUMB[34][21] ,
         \SUMB[34][20] , \SUMB[34][19] , \SUMB[34][18] , \SUMB[34][17] ,
         \SUMB[34][16] , \SUMB[34][15] , \SUMB[34][14] , \SUMB[34][13] ,
         \SUMB[34][12] , \SUMB[34][11] , \SUMB[34][10] , \SUMB[34][9] ,
         \SUMB[34][8] , \SUMB[34][7] , \SUMB[34][6] , \SUMB[34][5] ,
         \SUMB[34][4] , \SUMB[34][3] , \SUMB[34][2] , \SUMB[34][1] ,
         \SUMB[33][46] , \SUMB[33][45] , \SUMB[33][44] , \SUMB[33][43] ,
         \SUMB[33][42] , \SUMB[33][41] , \SUMB[33][40] , \SUMB[33][39] ,
         \SUMB[33][38] , \SUMB[33][37] , \SUMB[33][36] , \SUMB[33][35] ,
         \SUMB[33][34] , \SUMB[33][33] , \SUMB[33][32] , \SUMB[33][31] ,
         \SUMB[33][30] , \SUMB[33][29] , \SUMB[33][28] , \SUMB[33][27] ,
         \SUMB[33][26] , \SUMB[33][25] , \SUMB[33][24] , \SUMB[33][23] ,
         \SUMB[33][22] , \SUMB[33][21] , \SUMB[33][20] , \SUMB[33][19] ,
         \SUMB[33][18] , \SUMB[33][17] , \SUMB[33][16] , \SUMB[33][15] ,
         \SUMB[33][14] , \SUMB[33][13] , \SUMB[33][12] , \SUMB[33][11] ,
         \SUMB[33][10] , \SUMB[33][9] , \SUMB[33][8] , \SUMB[33][7] ,
         \SUMB[33][6] , \SUMB[33][5] , \SUMB[33][4] , \SUMB[33][3] ,
         \SUMB[33][2] , \SUMB[33][1] , \SUMB[32][46] , \SUMB[32][45] ,
         \SUMB[32][44] , \SUMB[32][43] , \SUMB[32][42] , \SUMB[32][41] ,
         \SUMB[32][40] , \SUMB[32][39] , \SUMB[32][38] , \SUMB[32][37] ,
         \SUMB[32][36] , \SUMB[32][35] , \SUMB[32][34] , \SUMB[32][33] ,
         \SUMB[32][32] , \SUMB[32][31] , \SUMB[32][30] , \SUMB[32][29] ,
         \SUMB[32][28] , \SUMB[32][27] , \SUMB[32][26] , \SUMB[32][25] ,
         \SUMB[32][24] , \SUMB[32][23] , \SUMB[32][22] , \SUMB[32][21] ,
         \SUMB[32][20] , \SUMB[32][19] , \SUMB[32][18] , \SUMB[32][17] ,
         \SUMB[32][16] , \SUMB[32][15] , \SUMB[32][14] , \SUMB[32][13] ,
         \SUMB[32][12] , \SUMB[32][11] , \SUMB[32][10] , \SUMB[32][9] ,
         \SUMB[32][8] , \SUMB[32][7] , \SUMB[32][6] , \SUMB[32][5] ,
         \SUMB[32][4] , \SUMB[32][3] , \SUMB[32][2] , \SUMB[32][1] ,
         \SUMB[31][46] , \SUMB[31][45] , \SUMB[31][44] , \SUMB[31][43] ,
         \SUMB[31][42] , \SUMB[31][41] , \SUMB[31][40] , \SUMB[31][39] ,
         \SUMB[31][38] , \SUMB[31][37] , \SUMB[31][36] , \SUMB[31][35] ,
         \SUMB[31][34] , \SUMB[31][33] , \SUMB[31][32] , \SUMB[31][31] ,
         \SUMB[31][30] , \SUMB[31][29] , \SUMB[31][28] , \SUMB[31][27] ,
         \SUMB[31][26] , \SUMB[31][25] , \SUMB[31][24] , \SUMB[31][23] ,
         \SUMB[31][22] , \SUMB[31][21] , \SUMB[31][20] , \SUMB[31][19] ,
         \SUMB[31][18] , \SUMB[31][17] , \SUMB[31][16] , \SUMB[31][15] ,
         \SUMB[31][14] , \SUMB[31][13] , \SUMB[31][12] , \SUMB[31][11] ,
         \SUMB[31][10] , \SUMB[31][9] , \SUMB[31][8] , \SUMB[31][7] ,
         \SUMB[31][6] , \SUMB[31][5] , \SUMB[31][4] , \SUMB[31][3] ,
         \SUMB[31][2] , \SUMB[31][1] , \SUMB[30][46] , \SUMB[30][45] ,
         \SUMB[30][44] , \SUMB[30][43] , \SUMB[30][42] , \SUMB[30][41] ,
         \SUMB[30][40] , \SUMB[30][39] , \SUMB[30][38] , \SUMB[30][37] ,
         \SUMB[30][36] , \SUMB[30][35] , \SUMB[30][34] , \SUMB[30][33] ,
         \SUMB[30][32] , \SUMB[30][31] , \SUMB[30][30] , \SUMB[30][29] ,
         \SUMB[30][28] , \SUMB[30][27] , \SUMB[30][26] , \SUMB[30][25] ,
         \SUMB[30][24] , \SUMB[30][23] , \SUMB[30][22] , \SUMB[30][21] ,
         \SUMB[30][20] , \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] ,
         \SUMB[30][16] , \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] ,
         \SUMB[30][12] , \SUMB[30][11] , \SUMB[30][9] , \SUMB[30][8] ,
         \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] , \SUMB[30][4] ,
         \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] , \SUMB[29][46] ,
         \SUMB[29][45] , \SUMB[29][44] , \SUMB[29][43] , \SUMB[29][42] ,
         \SUMB[29][41] , \SUMB[29][40] , \SUMB[29][39] , \SUMB[29][38] ,
         \SUMB[29][37] , \SUMB[29][36] , \SUMB[29][35] , \SUMB[29][34] ,
         \SUMB[29][33] , \SUMB[29][32] , \SUMB[29][31] , \SUMB[29][30] ,
         \SUMB[29][29] , \SUMB[29][28] , \SUMB[29][27] , \SUMB[29][26] ,
         \SUMB[29][25] , \SUMB[29][24] , \SUMB[29][23] , \SUMB[29][22] ,
         \SUMB[29][21] , \SUMB[29][20] , \SUMB[29][19] , \SUMB[29][18] ,
         \SUMB[29][17] , \SUMB[29][16] , \SUMB[29][15] , \SUMB[29][14] ,
         \SUMB[29][13] , \SUMB[29][12] , \SUMB[29][11] , \SUMB[29][10] ,
         \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] , \SUMB[29][6] ,
         \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] , \SUMB[29][2] ,
         \SUMB[29][1] , \SUMB[28][46] , \SUMB[28][45] , \SUMB[28][44] ,
         \SUMB[28][43] , \SUMB[28][42] , \SUMB[28][41] , \SUMB[28][40] ,
         \SUMB[28][39] , \SUMB[28][38] , \SUMB[28][37] , \SUMB[28][36] ,
         \SUMB[28][35] , \SUMB[28][34] , \SUMB[28][33] , \SUMB[28][32] ,
         \SUMB[28][31] , \SUMB[28][30] , \SUMB[28][29] , \SUMB[28][28] ,
         \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] , \SUMB[28][24] ,
         \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] , \SUMB[28][20] ,
         \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] , \SUMB[28][16] ,
         \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] , \SUMB[28][12] ,
         \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] , \SUMB[28][8] ,
         \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] , \SUMB[28][4] ,
         \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][46] ,
         \SUMB[27][45] , \SUMB[27][44] , \SUMB[27][43] , \SUMB[27][42] ,
         \SUMB[27][41] , \SUMB[27][40] , \SUMB[27][39] , \SUMB[27][38] ,
         \SUMB[27][37] , \SUMB[27][36] , \SUMB[27][35] , \SUMB[27][34] ,
         \SUMB[27][33] , \SUMB[27][32] , \SUMB[27][31] , \SUMB[27][30] ,
         \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] , \SUMB[27][26] ,
         \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] , \SUMB[27][22] ,
         \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] , \SUMB[27][18] ,
         \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] , \SUMB[27][14] ,
         \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] , \SUMB[27][10] ,
         \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] , \SUMB[27][6] ,
         \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] , \SUMB[27][2] ,
         \SUMB[27][1] , \SUMB[26][46] , \SUMB[26][45] , \SUMB[26][44] ,
         \SUMB[26][43] , \SUMB[26][42] , \SUMB[26][41] , \SUMB[26][40] ,
         \SUMB[26][39] , \SUMB[26][38] , \SUMB[26][37] , \SUMB[26][36] ,
         \SUMB[26][35] , \SUMB[26][34] , \SUMB[26][33] , \SUMB[26][32] ,
         \CARRYB[47][46] , \CARRYB[47][45] , \CARRYB[47][44] ,
         \CARRYB[47][43] , \CARRYB[47][42] , \CARRYB[47][41] ,
         \CARRYB[47][40] , \CARRYB[47][39] , \CARRYB[47][38] ,
         \CARRYB[47][37] , \CARRYB[47][36] , \CARRYB[47][35] ,
         \CARRYB[47][34] , \CARRYB[47][33] , \CARRYB[47][32] ,
         \CARRYB[47][31] , \CARRYB[47][30] , \CARRYB[47][29] ,
         \CARRYB[47][28] , \CARRYB[47][27] , \CARRYB[47][26] ,
         \CARRYB[47][25] , \CARRYB[47][24] , \CARRYB[47][23] ,
         \CARRYB[47][22] , \CARRYB[47][21] , \CARRYB[47][20] ,
         \CARRYB[47][19] , \CARRYB[47][18] , \CARRYB[47][17] ,
         \CARRYB[47][16] , \CARRYB[47][15] , \CARRYB[47][14] ,
         \CARRYB[47][13] , \CARRYB[47][12] , \CARRYB[47][11] ,
         \CARRYB[47][10] , \CARRYB[47][9] , \CARRYB[47][8] , \CARRYB[47][7] ,
         \CARRYB[47][6] , \CARRYB[47][5] , \CARRYB[47][4] , \CARRYB[47][3] ,
         \CARRYB[47][2] , \CARRYB[47][1] , \CARRYB[47][0] , \CARRYB[46][46] ,
         \CARRYB[46][45] , \CARRYB[46][44] , \CARRYB[46][43] ,
         \CARRYB[46][42] , \CARRYB[46][41] , \CARRYB[46][40] ,
         \CARRYB[46][39] , \CARRYB[46][38] , \CARRYB[46][37] ,
         \CARRYB[46][36] , \CARRYB[46][35] , \CARRYB[46][34] ,
         \CARRYB[46][33] , \CARRYB[46][32] , \CARRYB[46][31] ,
         \CARRYB[46][30] , \CARRYB[46][29] , \CARRYB[46][28] ,
         \CARRYB[46][27] , \CARRYB[46][26] , \CARRYB[46][25] ,
         \CARRYB[46][24] , \CARRYB[46][23] , \CARRYB[46][22] ,
         \CARRYB[46][21] , \CARRYB[46][20] , \CARRYB[46][19] ,
         \CARRYB[46][18] , \CARRYB[46][17] , \CARRYB[46][16] ,
         \CARRYB[46][15] , \CARRYB[46][14] , \CARRYB[46][13] ,
         \CARRYB[46][12] , \CARRYB[46][11] , \CARRYB[46][10] , \CARRYB[46][9] ,
         \CARRYB[46][8] , \CARRYB[46][7] , \CARRYB[46][6] , \CARRYB[46][5] ,
         \CARRYB[46][4] , \CARRYB[46][3] , \CARRYB[46][2] , \CARRYB[46][1] ,
         \CARRYB[46][0] , \CARRYB[45][46] , \CARRYB[45][45] , \CARRYB[45][44] ,
         \CARRYB[45][43] , \CARRYB[45][42] , \CARRYB[45][41] ,
         \CARRYB[45][40] , \CARRYB[45][39] , \CARRYB[45][38] ,
         \CARRYB[45][37] , \CARRYB[45][36] , \CARRYB[45][35] ,
         \CARRYB[45][34] , \CARRYB[45][33] , \CARRYB[45][32] ,
         \CARRYB[45][31] , \CARRYB[45][30] , \CARRYB[45][29] ,
         \CARRYB[45][28] , \CARRYB[45][27] , \CARRYB[45][26] ,
         \CARRYB[45][25] , \CARRYB[45][24] , \CARRYB[45][23] ,
         \CARRYB[45][22] , \CARRYB[45][21] , \CARRYB[45][20] ,
         \CARRYB[45][19] , \CARRYB[45][18] , \CARRYB[45][17] ,
         \CARRYB[45][16] , \CARRYB[45][15] , \CARRYB[45][14] ,
         \CARRYB[45][13] , \CARRYB[45][12] , \CARRYB[45][11] ,
         \CARRYB[45][10] , \CARRYB[45][9] , \CARRYB[45][8] , \CARRYB[45][7] ,
         \CARRYB[45][6] , \CARRYB[45][5] , \CARRYB[45][4] , \CARRYB[45][3] ,
         \CARRYB[45][2] , \CARRYB[45][1] , \CARRYB[45][0] , \CARRYB[44][46] ,
         \CARRYB[44][45] , \CARRYB[44][44] , \CARRYB[44][43] ,
         \CARRYB[44][42] , \CARRYB[44][41] , \CARRYB[44][40] ,
         \CARRYB[44][39] , \CARRYB[44][38] , \CARRYB[44][37] ,
         \CARRYB[44][36] , \CARRYB[44][35] , \CARRYB[44][34] ,
         \CARRYB[44][33] , \CARRYB[44][32] , \CARRYB[44][31] ,
         \CARRYB[44][30] , \CARRYB[44][29] , \CARRYB[44][28] ,
         \CARRYB[44][27] , \CARRYB[44][26] , \CARRYB[44][25] ,
         \CARRYB[44][24] , \CARRYB[44][23] , \CARRYB[44][22] ,
         \CARRYB[44][21] , \CARRYB[44][20] , \CARRYB[44][19] ,
         \CARRYB[44][18] , \CARRYB[44][17] , \CARRYB[44][16] ,
         \CARRYB[44][15] , \CARRYB[44][14] , \CARRYB[44][13] ,
         \CARRYB[44][12] , \CARRYB[44][11] , \CARRYB[44][10] , \CARRYB[44][9] ,
         \CARRYB[44][8] , \CARRYB[44][7] , \CARRYB[44][6] , \CARRYB[44][5] ,
         \CARRYB[44][4] , \CARRYB[44][3] , \CARRYB[44][2] , \CARRYB[44][1] ,
         \CARRYB[44][0] , \CARRYB[43][46] , \CARRYB[43][45] , \CARRYB[43][44] ,
         \CARRYB[43][43] , \CARRYB[43][42] , \CARRYB[43][41] ,
         \CARRYB[43][40] , \CARRYB[43][39] , \CARRYB[43][38] ,
         \CARRYB[43][37] , \CARRYB[43][36] , \CARRYB[43][35] ,
         \CARRYB[43][34] , \CARRYB[43][33] , \CARRYB[43][32] ,
         \CARRYB[43][31] , \CARRYB[43][30] , \CARRYB[43][29] ,
         \CARRYB[43][28] , \CARRYB[43][27] , \CARRYB[43][26] ,
         \CARRYB[43][25] , \CARRYB[43][24] , \CARRYB[43][23] ,
         \CARRYB[43][22] , \CARRYB[43][21] , \CARRYB[43][20] ,
         \CARRYB[43][19] , \CARRYB[43][18] , \CARRYB[43][17] ,
         \CARRYB[43][16] , \CARRYB[43][15] , \CARRYB[43][14] ,
         \CARRYB[43][13] , \CARRYB[43][12] , \CARRYB[43][11] ,
         \CARRYB[43][10] , \CARRYB[43][9] , \CARRYB[43][8] , \CARRYB[43][7] ,
         \CARRYB[43][6] , \CARRYB[43][5] , \CARRYB[43][4] , \CARRYB[43][3] ,
         \CARRYB[43][2] , \CARRYB[43][1] , \CARRYB[43][0] , \CARRYB[42][46] ,
         \CARRYB[42][45] , \CARRYB[42][44] , \CARRYB[42][43] ,
         \CARRYB[42][42] , \CARRYB[42][41] , \CARRYB[42][40] ,
         \CARRYB[42][39] , \CARRYB[42][38] , \CARRYB[42][37] ,
         \CARRYB[42][36] , \CARRYB[42][35] , \CARRYB[42][34] ,
         \CARRYB[42][33] , \CARRYB[42][32] , \CARRYB[42][31] ,
         \CARRYB[42][30] , \CARRYB[42][29] , \CARRYB[42][28] ,
         \CARRYB[42][27] , \CARRYB[42][26] , \CARRYB[42][25] ,
         \CARRYB[42][24] , \CARRYB[42][23] , \CARRYB[42][22] ,
         \CARRYB[42][21] , \CARRYB[42][20] , \CARRYB[42][19] ,
         \CARRYB[42][18] , \CARRYB[42][17] , \CARRYB[42][16] ,
         \CARRYB[42][15] , \CARRYB[42][14] , \CARRYB[42][13] ,
         \CARRYB[42][12] , \CARRYB[42][11] , \CARRYB[42][10] , \CARRYB[42][9] ,
         \CARRYB[42][8] , \CARRYB[42][7] , \CARRYB[42][6] , \CARRYB[42][5] ,
         \CARRYB[42][4] , \CARRYB[42][3] , \CARRYB[42][2] , \CARRYB[42][1] ,
         \CARRYB[42][0] , \CARRYB[41][46] , \CARRYB[41][45] , \CARRYB[41][44] ,
         \CARRYB[41][43] , \CARRYB[41][42] , \CARRYB[41][41] ,
         \CARRYB[41][40] , \CARRYB[41][39] , \CARRYB[41][38] ,
         \CARRYB[41][37] , \CARRYB[41][36] , \CARRYB[41][35] ,
         \CARRYB[41][34] , \CARRYB[41][33] , \CARRYB[41][32] ,
         \CARRYB[41][31] , \CARRYB[41][30] , \CARRYB[41][29] ,
         \CARRYB[41][28] , \CARRYB[41][27] , \CARRYB[41][26] ,
         \CARRYB[41][25] , \CARRYB[41][24] , \CARRYB[41][23] ,
         \CARRYB[41][22] , \CARRYB[41][21] , \CARRYB[41][20] ,
         \CARRYB[41][19] , \CARRYB[41][18] , \CARRYB[41][17] ,
         \CARRYB[41][16] , \CARRYB[41][15] , \CARRYB[41][14] ,
         \CARRYB[41][13] , \CARRYB[41][12] , \CARRYB[41][11] ,
         \CARRYB[41][10] , \CARRYB[41][9] , \CARRYB[41][8] , \CARRYB[41][7] ,
         \CARRYB[41][6] , \CARRYB[41][5] , \CARRYB[41][4] , \CARRYB[41][3] ,
         \CARRYB[41][2] , \CARRYB[41][1] , \CARRYB[41][0] , \CARRYB[40][46] ,
         \CARRYB[40][45] , \CARRYB[40][44] , \CARRYB[40][43] ,
         \CARRYB[40][42] , \CARRYB[40][41] , \CARRYB[40][40] ,
         \CARRYB[40][39] , \CARRYB[40][38] , \CARRYB[40][37] ,
         \CARRYB[40][36] , \CARRYB[40][35] , \CARRYB[40][34] ,
         \CARRYB[40][33] , \CARRYB[40][32] , \CARRYB[40][31] ,
         \CARRYB[40][30] , \CARRYB[40][29] , \CARRYB[40][28] ,
         \CARRYB[40][27] , \CARRYB[40][26] , \CARRYB[40][25] ,
         \CARRYB[40][24] , \CARRYB[40][23] , \CARRYB[40][22] ,
         \CARRYB[40][21] , \CARRYB[40][20] , \CARRYB[40][19] ,
         \CARRYB[40][18] , \CARRYB[40][17] , \CARRYB[40][16] ,
         \CARRYB[40][15] , \CARRYB[40][14] , \CARRYB[40][13] ,
         \CARRYB[40][12] , \CARRYB[40][11] , \CARRYB[40][10] , \CARRYB[40][9] ,
         \CARRYB[40][8] , \CARRYB[40][7] , \CARRYB[40][6] , \CARRYB[40][5] ,
         \CARRYB[40][4] , \CARRYB[40][3] , \CARRYB[40][2] , \CARRYB[40][1] ,
         \CARRYB[40][0] , \CARRYB[39][46] , \CARRYB[39][45] , \CARRYB[39][44] ,
         \CARRYB[39][43] , \CARRYB[39][42] , \CARRYB[39][41] ,
         \CARRYB[39][40] , \CARRYB[39][39] , \CARRYB[39][38] ,
         \CARRYB[39][37] , \CARRYB[39][36] , \CARRYB[39][35] ,
         \CARRYB[39][34] , \CARRYB[39][33] , \CARRYB[39][32] ,
         \CARRYB[39][31] , \CARRYB[39][30] , \CARRYB[39][29] ,
         \CARRYB[39][28] , \CARRYB[39][27] , \CARRYB[39][26] ,
         \CARRYB[39][25] , \CARRYB[39][24] , \CARRYB[39][23] ,
         \CARRYB[39][22] , \CARRYB[39][21] , \CARRYB[39][20] ,
         \CARRYB[39][19] , \CARRYB[39][18] , \CARRYB[39][17] ,
         \CARRYB[39][16] , \CARRYB[39][15] , \CARRYB[39][14] ,
         \CARRYB[39][13] , \CARRYB[39][12] , \CARRYB[39][11] ,
         \CARRYB[39][10] , \CARRYB[39][9] , \CARRYB[39][8] , \CARRYB[39][7] ,
         \CARRYB[39][6] , \CARRYB[39][5] , \CARRYB[39][4] , \CARRYB[39][3] ,
         \CARRYB[39][2] , \CARRYB[39][1] , \CARRYB[39][0] , \CARRYB[38][46] ,
         \CARRYB[38][45] , \CARRYB[38][44] , \CARRYB[38][43] ,
         \CARRYB[38][42] , \CARRYB[38][41] , \CARRYB[38][40] ,
         \CARRYB[38][39] , \CARRYB[38][38] , \CARRYB[38][37] ,
         \CARRYB[38][36] , \CARRYB[38][35] , \CARRYB[38][34] ,
         \CARRYB[38][33] , \CARRYB[38][32] , \CARRYB[38][31] ,
         \CARRYB[38][30] , \CARRYB[38][29] , \CARRYB[38][28] ,
         \CARRYB[38][27] , \CARRYB[38][26] , \CARRYB[38][25] ,
         \CARRYB[38][24] , \CARRYB[38][23] , \CARRYB[38][22] ,
         \CARRYB[38][21] , \CARRYB[38][20] , \CARRYB[38][19] ,
         \CARRYB[38][18] , \CARRYB[38][17] , \CARRYB[38][16] ,
         \CARRYB[38][15] , \CARRYB[38][14] , \CARRYB[38][13] ,
         \CARRYB[38][12] , \CARRYB[38][11] , \CARRYB[38][10] , \CARRYB[38][9] ,
         \CARRYB[38][8] , \CARRYB[38][7] , \CARRYB[38][6] , \CARRYB[38][5] ,
         \CARRYB[38][4] , \CARRYB[38][3] , \CARRYB[38][2] , \CARRYB[38][1] ,
         \CARRYB[38][0] , \CARRYB[37][46] , \CARRYB[37][45] , \CARRYB[37][44] ,
         \CARRYB[37][43] , \CARRYB[37][42] , \CARRYB[37][41] ,
         \CARRYB[37][40] , \CARRYB[37][39] , \CARRYB[37][38] ,
         \CARRYB[37][37] , \CARRYB[37][36] , \CARRYB[37][35] ,
         \CARRYB[37][34] , \CARRYB[37][33] , \CARRYB[37][32] ,
         \CARRYB[37][31] , \CARRYB[37][30] , \CARRYB[37][29] ,
         \CARRYB[37][28] , \CARRYB[37][27] , \CARRYB[37][26] ,
         \CARRYB[37][25] , \CARRYB[37][24] , \CARRYB[37][23] ,
         \CARRYB[37][22] , \CARRYB[37][21] , \CARRYB[37][20] ,
         \CARRYB[37][19] , \CARRYB[37][18] , \CARRYB[37][17] ,
         \CARRYB[37][16] , \SUMB[47][45] , \SUMB[47][44] , \SUMB[47][43] ,
         \SUMB[47][42] , \SUMB[47][41] , \SUMB[47][40] , \SUMB[47][39] ,
         \SUMB[47][38] , \SUMB[47][37] , \SUMB[47][36] , \SUMB[47][35] ,
         \SUMB[47][34] , \SUMB[47][33] , \SUMB[47][32] , \SUMB[47][31] ,
         \SUMB[47][30] , \SUMB[47][29] , \SUMB[47][28] , \SUMB[47][27] ,
         \SUMB[47][26] , \SUMB[47][25] , \SUMB[47][24] , \SUMB[47][23] ,
         \SUMB[47][22] , \SUMB[47][21] , \SUMB[47][20] , \SUMB[47][19] ,
         \SUMB[47][18] , \SUMB[47][17] , \SUMB[47][16] , \SUMB[47][15] ,
         \SUMB[47][14] , \SUMB[47][13] , \SUMB[47][12] , \SUMB[47][11] ,
         \SUMB[47][10] , \SUMB[47][9] , \SUMB[47][8] , \SUMB[47][7] ,
         \SUMB[47][6] , \SUMB[47][5] , \SUMB[47][4] , \SUMB[47][3] ,
         \SUMB[47][2] , \SUMB[47][1] , \SUMB[47][0] , \SUMB[46][46] ,
         \SUMB[46][45] , \SUMB[46][44] , \SUMB[46][43] , \SUMB[46][42] ,
         \SUMB[46][41] , \SUMB[46][40] , \SUMB[46][39] , \SUMB[46][38] ,
         \SUMB[46][37] , \SUMB[46][36] , \SUMB[46][35] , \SUMB[46][34] ,
         \SUMB[46][33] , \SUMB[46][32] , \SUMB[46][31] , \SUMB[46][30] ,
         \SUMB[46][29] , \SUMB[46][28] , \SUMB[46][27] , \SUMB[46][26] ,
         \SUMB[46][25] , \SUMB[46][24] , \SUMB[46][23] , \SUMB[46][22] ,
         \SUMB[46][21] , \SUMB[46][20] , \SUMB[46][19] , \SUMB[46][18] ,
         \SUMB[46][17] , \SUMB[46][16] , \SUMB[46][15] , \SUMB[46][14] ,
         \SUMB[46][13] , \SUMB[46][12] , \SUMB[46][11] , \SUMB[46][10] ,
         \SUMB[46][9] , \SUMB[46][8] , \SUMB[46][7] , \SUMB[46][6] ,
         \SUMB[46][5] , \SUMB[46][4] , \SUMB[46][3] , \SUMB[46][2] ,
         \SUMB[46][1] , \SUMB[45][46] , \SUMB[45][45] , \SUMB[45][44] ,
         \SUMB[45][43] , \SUMB[45][42] , \SUMB[45][41] , \SUMB[45][40] ,
         \SUMB[45][39] , \SUMB[45][38] , \SUMB[45][37] , \SUMB[45][36] ,
         \SUMB[45][35] , \SUMB[45][34] , \SUMB[45][33] , \SUMB[45][32] ,
         \SUMB[45][31] , \SUMB[45][30] , \SUMB[45][29] , \SUMB[45][28] ,
         \SUMB[45][27] , \SUMB[45][26] , \SUMB[45][25] , \SUMB[45][24] ,
         \SUMB[45][23] , \SUMB[45][22] , \SUMB[45][21] , \SUMB[45][20] ,
         \SUMB[45][19] , \SUMB[45][18] , \SUMB[45][17] , \SUMB[45][16] ,
         \SUMB[45][15] , \SUMB[45][14] , \SUMB[45][13] , \SUMB[45][12] ,
         \SUMB[45][11] , \SUMB[45][10] , \SUMB[45][9] , \SUMB[45][8] ,
         \SUMB[45][7] , \SUMB[45][6] , \SUMB[45][5] , \SUMB[45][4] ,
         \SUMB[45][3] , \SUMB[45][2] , \SUMB[45][1] , \SUMB[44][46] ,
         \SUMB[44][45] , \SUMB[44][44] , \SUMB[44][43] , \SUMB[44][42] ,
         \SUMB[44][41] , \SUMB[44][40] , \SUMB[44][39] , \SUMB[44][38] ,
         \SUMB[44][37] , \SUMB[44][36] , \SUMB[44][35] , \SUMB[44][34] ,
         \SUMB[44][33] , \SUMB[44][32] , \SUMB[44][31] , \SUMB[44][30] ,
         \SUMB[44][29] , \SUMB[44][28] , \SUMB[44][27] , \SUMB[44][26] ,
         \SUMB[44][25] , \SUMB[44][24] , \SUMB[44][23] , \SUMB[44][22] ,
         \SUMB[44][21] , \SUMB[44][20] , \SUMB[44][19] , \SUMB[44][18] ,
         \SUMB[44][17] , \SUMB[44][16] , \SUMB[44][15] , \SUMB[44][14] ,
         \SUMB[44][13] , \SUMB[44][12] , \SUMB[44][11] , \SUMB[44][10] ,
         \SUMB[44][9] , \SUMB[44][8] , \SUMB[44][7] , \SUMB[44][6] ,
         \SUMB[44][5] , \SUMB[44][4] , \SUMB[44][3] , \SUMB[44][2] ,
         \SUMB[44][1] , \SUMB[43][46] , \SUMB[43][45] , \SUMB[43][44] ,
         \SUMB[43][43] , \SUMB[43][42] , \SUMB[43][41] , \SUMB[43][40] ,
         \SUMB[43][39] , \SUMB[43][38] , \SUMB[43][37] , \SUMB[43][36] ,
         \SUMB[43][35] , \SUMB[43][34] , \SUMB[43][33] , \SUMB[43][32] ,
         \SUMB[43][31] , \SUMB[43][30] , \SUMB[43][29] , \SUMB[43][28] ,
         \SUMB[43][27] , \SUMB[43][26] , \SUMB[43][25] , \SUMB[43][24] ,
         \SUMB[43][23] , \SUMB[43][22] , \SUMB[43][21] , \SUMB[43][20] ,
         \SUMB[43][19] , \SUMB[43][18] , \SUMB[43][17] , \SUMB[43][16] ,
         \SUMB[43][15] , \SUMB[43][14] , \SUMB[43][13] , \SUMB[43][12] ,
         \SUMB[43][11] , \SUMB[43][10] , \SUMB[43][9] , \SUMB[43][8] ,
         \SUMB[43][7] , \SUMB[43][6] , \SUMB[43][5] , \SUMB[43][4] ,
         \SUMB[43][3] , \SUMB[43][2] , \SUMB[43][1] , \SUMB[42][46] ,
         \SUMB[42][45] , \SUMB[42][44] , \SUMB[42][43] , \SUMB[42][42] ,
         \SUMB[42][41] , \SUMB[42][40] , \SUMB[42][39] , \SUMB[42][38] ,
         \SUMB[42][37] , \SUMB[42][36] , \SUMB[42][35] , \SUMB[42][34] ,
         \SUMB[42][33] , \SUMB[42][32] , \SUMB[42][31] , \SUMB[42][30] ,
         \SUMB[42][29] , \SUMB[42][28] , \SUMB[42][27] , \SUMB[42][26] ,
         \SUMB[42][25] , \SUMB[42][24] , \SUMB[42][23] , \SUMB[42][22] ,
         \SUMB[42][21] , \SUMB[42][20] , \SUMB[42][19] , \SUMB[42][18] ,
         \SUMB[42][17] , \SUMB[42][16] , \SUMB[42][15] , \SUMB[42][14] ,
         \SUMB[42][13] , \SUMB[42][12] , \SUMB[42][11] , \SUMB[42][10] ,
         \SUMB[42][9] , \SUMB[42][8] , \SUMB[42][7] , \SUMB[42][6] ,
         \SUMB[42][5] , \SUMB[42][4] , \SUMB[42][3] , \SUMB[42][2] ,
         \SUMB[42][1] , \SUMB[41][46] , \SUMB[41][45] , \SUMB[41][44] ,
         \SUMB[41][43] , \SUMB[41][42] , \SUMB[41][41] , \SUMB[41][40] ,
         \SUMB[41][39] , \SUMB[41][38] , \SUMB[41][37] , \SUMB[41][36] ,
         \SUMB[41][35] , \SUMB[41][34] , \SUMB[41][33] , \SUMB[41][32] ,
         \SUMB[41][31] , \SUMB[41][30] , \SUMB[41][29] , \SUMB[41][28] ,
         \SUMB[41][27] , \SUMB[41][26] , \SUMB[41][25] , \SUMB[41][24] ,
         \SUMB[41][23] , \SUMB[41][22] , \SUMB[41][21] , \SUMB[41][20] ,
         \SUMB[41][19] , \SUMB[41][18] , \SUMB[41][17] , \SUMB[41][16] ,
         \SUMB[41][15] , \SUMB[41][14] , \SUMB[41][13] , \SUMB[41][12] ,
         \SUMB[41][11] , \SUMB[41][10] , \SUMB[41][9] , \SUMB[41][8] ,
         \SUMB[41][7] , \SUMB[41][6] , \SUMB[41][5] , \SUMB[41][4] ,
         \SUMB[41][3] , \SUMB[41][2] , \SUMB[41][1] , \SUMB[40][46] ,
         \SUMB[40][45] , \SUMB[40][44] , \SUMB[40][43] , \SUMB[40][42] ,
         \SUMB[40][41] , \SUMB[40][40] , \SUMB[40][39] , \SUMB[40][38] ,
         \SUMB[40][37] , \SUMB[40][36] , \SUMB[40][35] , \SUMB[40][34] ,
         \SUMB[40][33] , \SUMB[40][32] , \SUMB[40][31] , \SUMB[40][30] ,
         \SUMB[40][29] , \SUMB[40][28] , \SUMB[40][27] , \SUMB[40][26] ,
         \SUMB[40][25] , \SUMB[40][24] , \SUMB[40][23] , \SUMB[40][22] ,
         \SUMB[40][21] , \SUMB[40][20] , \SUMB[40][19] , \SUMB[40][18] ,
         \SUMB[40][17] , \SUMB[40][16] , \SUMB[40][15] , \SUMB[40][14] ,
         \SUMB[40][13] , \SUMB[40][12] , \SUMB[40][11] , \SUMB[40][10] ,
         \SUMB[40][9] , \SUMB[40][8] , \SUMB[40][7] , \SUMB[40][6] ,
         \SUMB[40][5] , \SUMB[40][4] , \SUMB[40][3] , \SUMB[40][2] ,
         \SUMB[40][1] , \SUMB[39][46] , \SUMB[39][45] , \SUMB[39][44] ,
         \SUMB[39][43] , \SUMB[39][42] , \SUMB[39][41] , \SUMB[39][40] ,
         \SUMB[39][39] , \SUMB[39][38] , \SUMB[39][37] , \SUMB[39][36] ,
         \SUMB[39][35] , \SUMB[39][34] , \SUMB[39][33] , \SUMB[39][32] ,
         \SUMB[39][31] , \SUMB[39][30] , \SUMB[39][29] , \SUMB[39][28] ,
         \SUMB[39][27] , \SUMB[39][26] , \SUMB[39][25] , \SUMB[39][24] ,
         \SUMB[39][23] , \SUMB[39][22] , \SUMB[39][21] , \SUMB[39][20] ,
         \SUMB[39][19] , \SUMB[39][18] , \SUMB[39][17] , \SUMB[39][16] ,
         \SUMB[39][15] , \SUMB[39][14] , \SUMB[39][13] , \SUMB[39][12] ,
         \SUMB[39][11] , \SUMB[39][10] , \SUMB[39][9] , \SUMB[39][8] ,
         \SUMB[39][7] , \SUMB[39][6] , \SUMB[39][5] , \SUMB[39][4] ,
         \SUMB[39][3] , \SUMB[39][2] , \SUMB[39][1] , \SUMB[38][46] ,
         \SUMB[38][45] , \SUMB[38][44] , \SUMB[38][43] , \SUMB[38][42] ,
         \SUMB[38][41] , \SUMB[38][40] , \SUMB[38][39] , \SUMB[38][38] ,
         \SUMB[38][37] , \SUMB[38][36] , \SUMB[38][35] , \SUMB[38][34] ,
         \SUMB[38][33] , \SUMB[38][32] , \SUMB[38][31] , \SUMB[38][30] ,
         \SUMB[38][29] , \SUMB[38][28] , \SUMB[38][27] , \SUMB[38][26] ,
         \SUMB[38][25] , \SUMB[38][24] , \SUMB[38][23] , \SUMB[38][22] ,
         \SUMB[38][21] , \SUMB[38][20] , \SUMB[38][19] , \SUMB[38][18] ,
         \SUMB[38][17] , \SUMB[38][16] , \SUMB[38][15] , \SUMB[38][14] ,
         \SUMB[38][13] , \SUMB[38][12] , \SUMB[38][11] , \SUMB[38][10] ,
         \SUMB[38][9] , \SUMB[38][8] , \SUMB[38][7] , \SUMB[38][6] ,
         \SUMB[38][5] , \SUMB[38][4] , \SUMB[38][3] , \SUMB[38][2] ,
         \SUMB[38][1] , \SUMB[37][46] , \SUMB[37][45] , \SUMB[37][44] ,
         \SUMB[37][43] , \SUMB[37][42] , \SUMB[37][41] , \SUMB[37][40] ,
         \SUMB[37][39] , \SUMB[37][38] , \SUMB[37][37] , \SUMB[37][36] ,
         \SUMB[37][35] , \SUMB[37][34] , \SUMB[37][33] , \SUMB[37][32] ,
         \SUMB[37][31] , \SUMB[37][30] , \SUMB[37][29] , \SUMB[37][28] ,
         \SUMB[37][27] , \SUMB[37][26] , \SUMB[37][25] , \SUMB[37][24] ,
         \SUMB[37][23] , \SUMB[37][22] , \SUMB[37][21] , \SUMB[37][20] ,
         \SUMB[37][19] , \SUMB[37][18] , \SUMB[37][17] , \SUMB[37][16] ,
         \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] ,
         \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] ,
         \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] ,
         \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] ,
         \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] ,
         \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] ,
         \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[44] , \A1[43] ,
         \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] ,
         \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] ,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] ,
         \A2[87] , \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] ,
         \A2[80] , \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] ,
         \A2[73] , \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] ,
         \A2[66] , \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] ,
         \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] ,
         \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n249, n250, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n269, n270, n277,
         n278, n279, n280, n284, n285, n286, n287, n289, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n312, n316, n318, n319, n320,
         n321, n322, n323, n324, n326, n327, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430;
  assign \ab[47][47]  = B[47];
  assign \ab[46][46]  = B[46];
  assign \ab[45][45]  = B[45];
  assign \ab[44][44]  = B[44];
  assign \ab[43][43]  = B[43];
  assign \ab[42][42]  = B[42];
  assign \ab[41][41]  = B[41];
  assign \ab[40][40]  = B[40];
  assign \ab[39][39]  = B[39];
  assign \ab[38][38]  = B[38];
  assign \ab[37][37]  = B[37];
  assign \ab[36][36]  = B[36];
  assign \ab[35][35]  = B[35];
  assign \ab[34][34]  = B[34];
  assign \ab[33][33]  = B[33];
  assign \ab[32][32]  = B[32];
  assign \ab[31][31]  = B[31];
  assign \ab[30][30]  = B[30];
  assign \ab[29][29]  = B[29];
  assign \ab[28][28]  = B[28];
  assign \ab[27][27]  = B[27];
  assign \ab[26][26]  = B[26];
  assign \ab[25][25]  = B[25];
  assign \ab[24][24]  = B[24];
  assign \ab[23][23]  = B[23];
  assign \ab[22][22]  = B[22];
  assign \ab[21][21]  = B[21];
  assign \ab[20][20]  = B[20];
  assign \ab[19][19]  = B[19];
  assign \ab[18][18]  = B[18];
  assign \ab[17][17]  = B[17];
  assign \ab[16][16]  = B[16];
  assign \ab[15][15]  = B[15];
  assign \ab[14][14]  = B[14];
  assign \ab[13][13]  = B[13];
  assign \ab[12][12]  = B[12];
  assign \ab[11][11]  = B[11];
  assign \ab[10][10]  = B[10];
  assign \ab[9][9]  = B[9];
  assign \ab[8][8]  = B[8];
  assign \ab[7][7]  = B[7];
  assign \ab[6][6]  = B[6];
  assign \ab[5][5]  = B[5];
  assign \ab[4][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[1][1]  = B[1];

  FA1AP S2_43_19 ( .A(\ab[43][19] ), .B(\CARRYB[42][19] ), .CI(\SUMB[42][20] ), 
        .CO(\CARRYB[43][19] ), .S(\SUMB[43][19] ) );
  FA1AP S2_23_32 ( .A(\ab[32][23] ), .B(\CARRYB[22][32] ), .CI(\SUMB[22][33] ), 
        .CO(\CARRYB[23][32] ), .S(\SUMB[23][32] ) );
  FA1AP S2_20_25 ( .A(\ab[25][20] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA1AP S2_11_20 ( .A(\CARRYB[10][20] ), .B(n627), .CI(\SUMB[10][21] ), .CO(
        \CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1AP S2_9_36 ( .A(\CARRYB[8][36] ), .B(n567), .CI(\SUMB[8][37] ), .CO(
        \CARRYB[9][36] ), .S(\SUMB[9][36] ) );
  FA1AP S2_2_35 ( .A(n2214), .B(\CARRYB[1][35] ), .CI(\SUMB[1][36] ), .CO(
        \CARRYB[2][35] ), .S(\SUMB[2][35] ) );
  LOG_POLY_DW01_add_5 FS_1 ( .A({1'b0, \A1[92] , \A1[91] , \A1[90] , \A1[89] , 
        \A1[88] , \A1[87] , \A1[86] , \A1[85] , \A1[84] , \A1[83] , \A1[82] , 
        \A1[81] , \A1[80] , \A1[79] , \A1[78] , \A1[77] , \A1[76] , \A1[75] , 
        \A1[74] , \A1[73] , \A1[72] , \A1[71] , \A1[70] , \A1[69] , \A1[68] , 
        \A1[67] , \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] , \A1[61] , 
        \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , 
        \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , 
        \A1[46] , \SUMB[47][0] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , 
        \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[93] , 
        \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] , \A2[86] , 
        \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] , \A2[79] , 
        \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] , \A2[72] , 
        \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] , \A2[65] , 
        \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , 
        \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , 
        \A2[50] , \A2[49] , \A2[48] , \A2[47] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[95:2])
         );
  FA1A S2_8_2 ( .A(n336), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1P S2_19_5 ( .A(n420), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), .CO(
        \CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1P S2_34_34 ( .A(\CARRYB[33][34] ), .B(n735), .CI(\SUMB[33][35] ), .CO(
        \CARRYB[34][34] ), .S(\SUMB[34][34] ) );
  FA1P S2_21_4 ( .A(n366), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), .CO(
        \CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1P S2_19_4 ( .A(n2301), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), .CO(
        \CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1P S2_20_4 ( .A(n2302), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), .CO(
        \CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA1P S2_19_19 ( .A(\CARRYB[18][19] ), .B(n2358), .CI(\SUMB[18][20] ), .CO(
        \CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA1P S2_12_18 ( .A(n664), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), .CO(
        \CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA1P S2_13_18 ( .A(\SUMB[12][19] ), .B(\CARRYB[12][18] ), .CI(n695), .CO(
        \CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA1P S2_24_18 ( .A(\CARRYB[23][18] ), .B(\ab[24][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA1P S2_32_18 ( .A(\CARRYB[31][18] ), .B(\ab[32][18] ), .CI(\SUMB[31][19] ), 
        .CO(\CARRYB[32][18] ), .S(\SUMB[32][18] ) );
  FA1P S2_33_18 ( .A(\CARRYB[32][18] ), .B(\ab[33][18] ), .CI(\SUMB[32][19] ), 
        .CO(\CARRYB[33][18] ), .S(\SUMB[33][18] ) );
  FA1P S2_40_1 ( .A(n2195), .B(\CARRYB[39][1] ), .CI(\SUMB[39][2] ), .CO(
        \CARRYB[40][1] ), .S(\SUMB[40][1] ) );
  FA1P S2_41_1 ( .A(n2222), .B(\CARRYB[40][1] ), .CI(\SUMB[40][2] ), .CO(
        \CARRYB[41][1] ), .S(\SUMB[41][1] ) );
  FA1P S2_26_25 ( .A(\CARRYB[25][25] ), .B(\ab[26][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA1P S2_34_24 ( .A(\ab[34][24] ), .B(\CARRYB[33][24] ), .CI(\SUMB[33][25] ), 
        .CO(\CARRYB[34][24] ), .S(\SUMB[34][24] ) );
  FA1P S2_35_3 ( .A(n2291), .B(\CARRYB[34][3] ), .CI(\SUMB[34][4] ), .CO(
        \CARRYB[35][3] ), .S(\SUMB[35][3] ) );
  FA1P S2_23_3 ( .A(n2271), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), .CO(
        \CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA1P S2_33_3 ( .A(n2275), .B(\CARRYB[32][3] ), .CI(\SUMB[32][4] ), .CO(
        \CARRYB[33][3] ), .S(\SUMB[33][3] ) );
  FA1P S2_34_3 ( .A(n2276), .B(\CARRYB[33][3] ), .CI(\SUMB[33][4] ), .CO(
        \CARRYB[34][3] ), .S(\SUMB[34][3] ) );
  FA1P S2_12_40 ( .A(\ab[40][12] ), .B(\CARRYB[11][40] ), .CI(\SUMB[11][41] ), 
        .CO(\CARRYB[12][40] ), .S(\SUMB[12][40] ) );
  FA1P S2_13_40 ( .A(\ab[40][13] ), .B(\CARRYB[12][40] ), .CI(\SUMB[12][41] ), 
        .CO(\CARRYB[13][40] ), .S(\SUMB[13][40] ) );
  FA1P S2_22_40 ( .A(\ab[40][22] ), .B(\CARRYB[21][40] ), .CI(\SUMB[21][41] ), 
        .CO(\CARRYB[22][40] ), .S(\SUMB[22][40] ) );
  FA1P S2_10_10 ( .A(n2339), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), .CO(
        \CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1P S2_23_35 ( .A(\ab[35][23] ), .B(\CARRYB[22][35] ), .CI(\SUMB[22][36] ), 
        .CO(\CARRYB[23][35] ), .S(\SUMB[23][35] ) );
  FA1P S2_24_35 ( .A(\ab[35][24] ), .B(\CARRYB[23][35] ), .CI(\SUMB[23][36] ), 
        .CO(\CARRYB[24][35] ), .S(\SUMB[24][35] ) );
  FA1P S2_12_7 ( .A(n508), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), .CO(
        \CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1P S2_22_7 ( .A(n506), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), .CO(
        \CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA1P S2_23_7 ( .A(n495), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), .CO(
        \CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA1P S2_42_7 ( .A(n505), .B(\CARRYB[41][7] ), .CI(\SUMB[41][8] ), .CO(
        \CARRYB[42][7] ), .S(\SUMB[42][7] ) );
  FA1P S2_24_7 ( .A(\SUMB[23][8] ), .B(\CARRYB[23][7] ), .CI(n500), .CO(
        \CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA1P S2_25_12 ( .A(n661), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), .CO(
        \CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA1P S2_24_6 ( .A(n462), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), .CO(
        \CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA1P S2_25_6 ( .A(n430), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), .CO(
        \CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA1P S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA1P S2_27_17 ( .A(\CARRYB[26][17] ), .B(\ab[27][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA1P S4_32 ( .A(\ab[47][32] ), .B(\CARRYB[46][32] ), .CI(\SUMB[46][33] ), 
        .CO(\CARRYB[47][32] ), .S(\SUMB[47][32] ) );
  FA1P S2_41_32 ( .A(\ab[41][32] ), .B(\CARRYB[40][32] ), .CI(\SUMB[40][33] ), 
        .CO(\CARRYB[41][32] ), .S(\SUMB[41][32] ) );
  FA1P S2_34_31 ( .A(\CARRYB[33][31] ), .B(\ab[34][31] ), .CI(\SUMB[33][32] ), 
        .CO(\CARRYB[34][31] ), .S(\SUMB[34][31] ) );
  FA1A S4_42 ( .A(\ab[47][42] ), .B(\CARRYB[46][42] ), .CI(\SUMB[46][43] ), 
        .CO(\CARRYB[47][42] ), .S(\SUMB[47][42] ) );
  FA1P S2_20_37 ( .A(\ab[37][20] ), .B(\CARRYB[19][37] ), .CI(\SUMB[19][38] ), 
        .CO(\CARRYB[20][37] ), .S(\SUMB[20][37] ) );
  FA1P S2_30_37 ( .A(\ab[37][30] ), .B(\CARRYB[29][37] ), .CI(\SUMB[29][38] ), 
        .CO(\CARRYB[30][37] ), .S(\SUMB[30][37] ) );
  FA1P S3_17_46 ( .A(\ab[46][17] ), .B(\CARRYB[16][46] ), .CI(\ab[47][16] ), 
        .CO(\CARRYB[17][46] ), .S(\SUMB[17][46] ) );
  FA1P S2_17_2 ( .A(n2262), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), .CO(
        \CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1P S2_22_36 ( .A(\ab[36][22] ), .B(\CARRYB[21][36] ), .CI(\SUMB[21][37] ), 
        .CO(\CARRYB[22][36] ), .S(\SUMB[22][36] ) );
  FA1 S4_34 ( .A(\ab[47][34] ), .B(\CARRYB[46][34] ), .CI(\SUMB[46][35] ), 
        .CO(\CARRYB[47][34] ), .S(\SUMB[47][34] ) );
  FA1P S2_34_39 ( .A(\ab[39][34] ), .B(\CARRYB[33][39] ), .CI(\SUMB[33][40] ), 
        .CO(\CARRYB[34][39] ), .S(\SUMB[34][39] ) );
  FA1P S2_13_39 ( .A(\ab[39][13] ), .B(\CARRYB[12][39] ), .CI(\SUMB[12][40] ), 
        .CO(\CARRYB[13][39] ), .S(\SUMB[13][39] ) );
  FA1P S2_23_39 ( .A(\ab[39][23] ), .B(\CARRYB[22][39] ), .CI(\SUMB[22][40] ), 
        .CO(\CARRYB[23][39] ), .S(\SUMB[23][39] ) );
  FA1P S2_24_39 ( .A(\ab[39][24] ), .B(\CARRYB[23][39] ), .CI(\SUMB[23][40] ), 
        .CO(\CARRYB[24][39] ), .S(\SUMB[24][39] ) );
  FA1P S2_7_5 ( .A(n304), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1P S2_17_5 ( .A(n398), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), .CO(
        \CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1P S2_18_5 ( .A(n415), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), .CO(
        \CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1P S2_28_5 ( .A(n412), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), .CO(
        \CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA1P S2_29_5 ( .A(n411), .B(\CARRYB[28][5] ), .CI(\SUMB[28][6] ), .CO(
        \CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA1A S2_10_5 ( .A(n424), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1P S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA1P S2_25_27 ( .A(\ab[27][25] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA1P S2_25_38 ( .A(\ab[38][25] ), .B(\CARRYB[24][38] ), .CI(\SUMB[24][39] ), 
        .CO(\CARRYB[25][38] ), .S(\SUMB[25][38] ) );
  FA1P S2_31_37 ( .A(\ab[37][31] ), .B(\CARRYB[30][37] ), .CI(\SUMB[30][38] ), 
        .CO(\CARRYB[31][37] ), .S(\SUMB[31][37] ) );
  FA1P S2_15_38 ( .A(\ab[38][15] ), .B(\CARRYB[14][38] ), .CI(\SUMB[14][39] ), 
        .CO(\CARRYB[15][38] ), .S(\SUMB[15][38] ) );
  FA1P S2_14_12 ( .A(\CARRYB[13][12] ), .B(n659), .CI(\SUMB[13][13] ), .CO(
        \CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1P S2_42_42 ( .A(n2413), .B(\CARRYB[41][42] ), .CI(\SUMB[41][43] ), .CO(
        \CARRYB[42][42] ), .S(\SUMB[42][42] ) );
  FA1P S2_27_1 ( .A(n2166), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), .CO(
        \CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA1P S4_2 ( .A(n339), .B(\CARRYB[46][2] ), .CI(\SUMB[46][3] ), .CO(
        \CARRYB[47][2] ), .S(\SUMB[47][2] ) );
  FA1P S2_8_22 ( .A(\CARRYB[7][22] ), .B(n539), .CI(\SUMB[7][23] ), .CO(
        \CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1P S2_23_36 ( .A(\ab[36][23] ), .B(\CARRYB[22][36] ), .CI(\SUMB[22][37] ), 
        .CO(\CARRYB[23][36] ), .S(\SUMB[23][36] ) );
  FA1P S2_35_30 ( .A(\ab[35][30] ), .B(\CARRYB[34][30] ), .CI(\SUMB[34][31] ), 
        .CO(\CARRYB[35][30] ), .S(\SUMB[35][30] ) );
  FA1P S2_36_30 ( .A(\ab[36][30] ), .B(\CARRYB[35][30] ), .CI(\SUMB[35][31] ), 
        .CO(\CARRYB[36][30] ), .S(\SUMB[36][30] ) );
  FA1P S2_10_43 ( .A(\ab[43][10] ), .B(\CARRYB[9][43] ), .CI(\SUMB[9][44] ), 
        .CO(\CARRYB[10][43] ), .S(\SUMB[10][43] ) );
  FA1A S2_45_39 ( .A(\ab[45][39] ), .B(\CARRYB[44][39] ), .CI(\SUMB[44][40] ), 
        .CO(\CARRYB[45][39] ), .S(\SUMB[45][39] ) );
  FA1P S2_14_17 ( .A(n710), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), .CO(
        \CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA1 S2_15_37 ( .A(\ab[37][15] ), .B(\CARRYB[14][37] ), .CI(\SUMB[14][38] ), 
        .CO(\CARRYB[15][37] ), .S(\SUMB[15][37] ) );
  FA1P S2_38_20 ( .A(\ab[38][20] ), .B(\CARRYB[37][20] ), .CI(\SUMB[37][21] ), 
        .CO(\CARRYB[38][20] ), .S(\SUMB[38][20] ) );
  FA1P S2_26_11 ( .A(n630), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), .CO(
        \CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA1P S2_27_6 ( .A(\SUMB[26][7] ), .B(\CARRYB[26][6] ), .CI(n442), .CO(
        \CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA1P S2_28_6 ( .A(n447), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), .CO(
        \CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA1P S2_21_5 ( .A(n395), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), .CO(
        \CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1P S2_37_38 ( .A(\ab[38][37] ), .B(\CARRYB[36][38] ), .CI(\SUMB[36][39] ), 
        .CO(\CARRYB[37][38] ), .S(\SUMB[37][38] ) );
  FA1P S2_21_40 ( .A(\ab[40][21] ), .B(\CARRYB[20][40] ), .CI(\SUMB[20][41] ), 
        .CO(\CARRYB[21][40] ), .S(\SUMB[21][40] ) );
  FA1P S2_35_13 ( .A(\CARRYB[34][13] ), .B(\ab[35][13] ), .CI(\SUMB[34][14] ), 
        .CO(\CARRYB[35][13] ), .S(\SUMB[35][13] ) );
  FA1P S2_43_42 ( .A(\ab[43][42] ), .B(\CARRYB[42][42] ), .CI(\SUMB[42][43] ), 
        .CO(\CARRYB[43][42] ), .S(\SUMB[43][42] ) );
  FA1P S2_44_42 ( .A(\ab[44][42] ), .B(\CARRYB[43][42] ), .CI(\SUMB[43][43] ), 
        .CO(\CARRYB[44][42] ), .S(\SUMB[44][42] ) );
  FA1P S2_13_13 ( .A(\CARRYB[12][13] ), .B(n2346), .CI(\SUMB[12][14] ), .CO(
        \CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1P S2_39_8 ( .A(n547), .B(\CARRYB[38][8] ), .CI(\SUMB[38][9] ), .CO(
        \CARRYB[39][8] ), .S(\SUMB[39][8] ) );
  FA1P S2_28_23 ( .A(\CARRYB[27][23] ), .B(\ab[28][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA1A S2_38_27 ( .A(\ab[38][27] ), .B(\CARRYB[37][27] ), .CI(\SUMB[37][28] ), 
        .CO(\CARRYB[38][27] ), .S(\SUMB[38][27] ) );
  FA1P S2_16_16 ( .A(\CARRYB[15][16] ), .B(n2352), .CI(\SUMB[15][17] ), .CO(
        \CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA1P S2_17_16 ( .A(\SUMB[16][17] ), .B(\ab[17][16] ), .CI(\CARRYB[16][16] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA1P S2_39_22 ( .A(\ab[39][22] ), .B(\CARRYB[38][22] ), .CI(\SUMB[38][23] ), 
        .CO(\CARRYB[39][22] ), .S(\SUMB[39][22] ) );
  FA1P S2_41_30 ( .A(\ab[41][30] ), .B(\CARRYB[40][30] ), .CI(\SUMB[40][31] ), 
        .CO(\CARRYB[41][30] ), .S(\SUMB[41][30] ) );
  FA1P S2_45_2 ( .A(n2247), .B(\CARRYB[44][2] ), .CI(\SUMB[44][3] ), .CO(
        \CARRYB[45][2] ), .S(\SUMB[45][2] ) );
  FA1P S2_46_2 ( .A(n2257), .B(\CARRYB[45][2] ), .CI(\SUMB[45][3] ), .CO(
        \CARRYB[46][2] ), .S(\SUMB[46][2] ) );
  FA1P S2_18_2 ( .A(n2216), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), .CO(
        \CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1 S4_40 ( .A(\ab[47][40] ), .B(\CARRYB[46][40] ), .CI(\SUMB[46][41] ), 
        .CO(\CARRYB[47][40] ), .S(\SUMB[47][40] ) );
  FA1P S2_33_22 ( .A(\ab[33][22] ), .B(\CARRYB[32][22] ), .CI(\SUMB[32][23] ), 
        .CO(\CARRYB[33][22] ), .S(\SUMB[33][22] ) );
  FA1P S2_32_21 ( .A(\ab[32][21] ), .B(\CARRYB[31][21] ), .CI(\SUMB[31][22] ), 
        .CO(\CARRYB[32][21] ), .S(\SUMB[32][21] ) );
  FA1P S2_14_40 ( .A(\CARRYB[13][40] ), .B(\ab[40][14] ), .CI(\SUMB[13][41] ), 
        .CO(\CARRYB[14][40] ), .S(\SUMB[14][40] ) );
  FA1P S2_29_39 ( .A(\ab[39][29] ), .B(\CARRYB[28][39] ), .CI(\SUMB[28][40] ), 
        .CO(\CARRYB[29][39] ), .S(\SUMB[29][39] ) );
  FA1P S2_12_39 ( .A(\ab[39][12] ), .B(\CARRYB[11][39] ), .CI(\SUMB[11][40] ), 
        .CO(\CARRYB[12][39] ), .S(\SUMB[12][39] ) );
  FA1A S2_8_9 ( .A(n552), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1P S2_17_20 ( .A(\ab[20][17] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA1P S2_18_20 ( .A(\CARRYB[17][20] ), .B(\ab[20][18] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA1P S2_42_18 ( .A(\CARRYB[41][18] ), .B(\ab[42][18] ), .CI(\SUMB[41][19] ), 
        .CO(\CARRYB[42][18] ), .S(\SUMB[42][18] ) );
  FA1P S2_43_18 ( .A(\CARRYB[42][18] ), .B(\ab[43][18] ), .CI(\SUMB[42][19] ), 
        .CO(\CARRYB[43][18] ), .S(\SUMB[43][18] ) );
  FA1P S3_16_46 ( .A(\ab[46][16] ), .B(\CARRYB[15][46] ), .CI(\ab[47][15] ), 
        .CO(\CARRYB[16][46] ), .S(\SUMB[16][46] ) );
  FA1P S2_43_20 ( .A(\ab[43][20] ), .B(\CARRYB[42][20] ), .CI(\SUMB[42][21] ), 
        .CO(\CARRYB[43][20] ), .S(\SUMB[43][20] ) );
  FA1A S2_10_34 ( .A(\CARRYB[9][34] ), .B(n590), .CI(\SUMB[9][35] ), .CO(
        \CARRYB[10][34] ), .S(\SUMB[10][34] ) );
  FA1P S2_8_41 ( .A(n546), .B(\CARRYB[7][41] ), .CI(\SUMB[7][42] ), .CO(
        \CARRYB[8][41] ), .S(\SUMB[8][41] ) );
  FA1P S2_9_41 ( .A(n612), .B(\CARRYB[8][41] ), .CI(\SUMB[8][42] ), .CO(
        \CARRYB[9][41] ), .S(\SUMB[9][41] ) );
  FA1P S2_21_8 ( .A(n526), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), .CO(
        \CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1P S2_36_38 ( .A(\ab[38][36] ), .B(\CARRYB[35][38] ), .CI(\SUMB[35][39] ), 
        .CO(\CARRYB[36][38] ), .S(\SUMB[36][38] ) );
  FA1P S2_15_3 ( .A(n340), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1P S2_39_33 ( .A(\ab[39][33] ), .B(\CARRYB[38][33] ), .CI(\SUMB[38][34] ), 
        .CO(\CARRYB[39][33] ), .S(\SUMB[39][33] ) );
  FA1P S2_40_33 ( .A(\ab[40][33] ), .B(\CARRYB[39][33] ), .CI(\SUMB[39][34] ), 
        .CO(\CARRYB[40][33] ), .S(\SUMB[40][33] ) );
  FA1A S2_46_39 ( .A(\ab[46][39] ), .B(\CARRYB[45][39] ), .CI(\SUMB[45][40] ), 
        .CO(\CARRYB[46][39] ), .S(\SUMB[46][39] ) );
  FA1P S2_9_44 ( .A(\ab[9][44] ), .B(\CARRYB[8][44] ), .CI(\SUMB[8][45] ), 
        .CO(\CARRYB[9][44] ), .S(\SUMB[9][44] ) );
  FA1P S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA1P S1_32_0 ( .A(n332), .B(\CARRYB[31][0] ), .CI(\SUMB[31][1] ), .CO(
        \CARRYB[32][0] ), .S(\A1[30] ) );
  FA1P S1_42_0 ( .A(n2225), .B(\CARRYB[41][0] ), .CI(\SUMB[41][1] ), .CO(
        \CARRYB[42][0] ), .S(\A1[40] ) );
  FA1P S2_27_12 ( .A(\CARRYB[26][12] ), .B(n663), .CI(\SUMB[26][13] ), .CO(
        \CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA1P S2_15_16 ( .A(n722), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), .CO(
        \CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA1P S2_14_38 ( .A(\ab[38][14] ), .B(\CARRYB[13][38] ), .CI(\SUMB[13][39] ), 
        .CO(\CARRYB[14][38] ), .S(\SUMB[14][38] ) );
  FA1P S2_32_37 ( .A(\ab[37][32] ), .B(\CARRYB[31][37] ), .CI(\SUMB[31][38] ), 
        .CO(\CARRYB[32][37] ), .S(\SUMB[32][37] ) );
  FA1A S2_39_13 ( .A(\ab[39][13] ), .B(\CARRYB[38][13] ), .CI(\SUMB[38][14] ), 
        .CO(\CARRYB[39][13] ), .S(\SUMB[39][13] ) );
  FA1P S2_24_4 ( .A(n365), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), .CO(
        \CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA1P S2_25_4 ( .A(n364), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), .CO(
        \CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA1P S2_43_2 ( .A(n2252), .B(\CARRYB[42][2] ), .CI(\SUMB[42][3] ), .CO(
        \CARRYB[43][2] ), .S(\SUMB[43][2] ) );
  FA1P S2_44_2 ( .A(n2248), .B(\CARRYB[43][2] ), .CI(\SUMB[43][3] ), .CO(
        \CARRYB[44][2] ), .S(\SUMB[44][2] ) );
  FA1P S2_10_19 ( .A(n608), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), .CO(
        \CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1P S2_25_8 ( .A(n538), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), .CO(
        \CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA1A S2_39_40 ( .A(\ab[40][39] ), .B(\CARRYB[38][40] ), .CI(\SUMB[38][41] ), 
        .CO(\CARRYB[39][40] ), .S(\SUMB[39][40] ) );
  FA1P S2_44_17 ( .A(\SUMB[43][18] ), .B(\CARRYB[43][17] ), .CI(\ab[44][17] ), 
        .CO(\CARRYB[44][17] ), .S(\SUMB[44][17] ) );
  FA1P S2_11_18 ( .A(n638), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), .CO(
        \CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1P S2_22_8 ( .A(n539), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), .CO(
        \CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA1P S2_46_34 ( .A(\ab[46][34] ), .B(\CARRYB[45][34] ), .CI(\SUMB[45][35] ), 
        .CO(\CARRYB[46][34] ), .S(\SUMB[46][34] ) );
  FA1P S2_43_34 ( .A(\ab[43][34] ), .B(\CARRYB[42][34] ), .CI(\SUMB[42][35] ), 
        .CO(\CARRYB[43][34] ), .S(\SUMB[43][34] ) );
  FA1A S2_13_41 ( .A(\CARRYB[12][41] ), .B(\ab[41][13] ), .CI(\SUMB[12][42] ), 
        .CO(\CARRYB[13][41] ), .S(\SUMB[13][41] ) );
  FA1 S2_36_40 ( .A(\ab[40][36] ), .B(\CARRYB[35][40] ), .CI(\SUMB[35][41] ), 
        .CO(\CARRYB[36][40] ), .S(\SUMB[36][40] ) );
  FA1P S2_28_24 ( .A(\CARRYB[27][24] ), .B(\ab[28][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA1P S2_7_41 ( .A(n499), .B(\CARRYB[6][41] ), .CI(\SUMB[6][42] ), .CO(
        \CARRYB[7][41] ), .S(\SUMB[7][41] ) );
  FA1P S2_27_7 ( .A(n498), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), .CO(
        \CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA1A S2_10_2 ( .A(n345), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1P S2_41_17 ( .A(\ab[41][17] ), .B(\CARRYB[40][17] ), .CI(\SUMB[40][18] ), 
        .CO(\CARRYB[41][17] ), .S(\SUMB[41][17] ) );
  FA1P S2_26_5 ( .A(n410), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), .CO(
        \CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA1P S2_20_15 ( .A(\CARRYB[19][15] ), .B(n724), .CI(\SUMB[19][16] ), .CO(
        \CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA1P S2_23_40 ( .A(\ab[40][23] ), .B(\CARRYB[22][40] ), .CI(\SUMB[22][41] ), 
        .CO(\CARRYB[23][40] ), .S(\SUMB[23][40] ) );
  FA1P S2_24_40 ( .A(\ab[40][24] ), .B(\CARRYB[23][40] ), .CI(\SUMB[23][41] ), 
        .CO(\CARRYB[24][40] ), .S(\SUMB[24][40] ) );
  FA1P S2_31_40 ( .A(\ab[40][31] ), .B(\CARRYB[30][40] ), .CI(\SUMB[30][41] ), 
        .CO(\CARRYB[31][40] ), .S(\SUMB[31][40] ) );
  FA1P S2_13_4 ( .A(n372), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), .CO(
        \CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_22_4 ( .A(n356), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), .CO(
        \CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA1P S2_31_31 ( .A(n2386), .B(\CARRYB[30][31] ), .CI(\SUMB[30][32] ), .CO(
        \CARRYB[31][31] ), .S(\SUMB[31][31] ) );
  FA1P S2_39_36 ( .A(\ab[39][36] ), .B(\CARRYB[38][36] ), .CI(\SUMB[38][37] ), 
        .CO(\CARRYB[39][36] ), .S(\SUMB[39][36] ) );
  FA1P S2_11_40 ( .A(\ab[40][11] ), .B(\CARRYB[10][40] ), .CI(\SUMB[10][41] ), 
        .CO(\CARRYB[11][40] ), .S(\SUMB[11][40] ) );
  FA1P S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA1P S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA1P S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA1P S2_30_31 ( .A(\ab[31][30] ), .B(\CARRYB[29][31] ), .CI(\SUMB[29][32] ), 
        .CO(\CARRYB[30][31] ), .S(\SUMB[30][31] ) );
  FA1 S2_8_37 ( .A(n551), .B(\CARRYB[7][37] ), .CI(\SUMB[7][38] ), .CO(
        \CARRYB[8][37] ), .S(\SUMB[8][37] ) );
  FA1P S2_45_42 ( .A(\ab[45][42] ), .B(\CARRYB[44][42] ), .CI(\SUMB[44][43] ), 
        .CO(\CARRYB[45][42] ), .S(\SUMB[45][42] ) );
  FA1P S2_46_42 ( .A(\ab[46][42] ), .B(\CARRYB[45][42] ), .CI(\SUMB[45][43] ), 
        .CO(\CARRYB[46][42] ), .S(\SUMB[46][42] ) );
  FA1P S3_11_46 ( .A(\ab[46][11] ), .B(\CARRYB[10][46] ), .CI(\ab[47][10] ), 
        .CO(\CARRYB[11][46] ), .S(\SUMB[11][46] ) );
  FA1P S3_12_46 ( .A(\ab[46][12] ), .B(\CARRYB[11][46] ), .CI(\ab[47][11] ), 
        .CO(\CARRYB[12][46] ), .S(\SUMB[12][46] ) );
  FA1P S2_35_16 ( .A(\ab[35][16] ), .B(\CARRYB[34][16] ), .CI(\SUMB[34][17] ), 
        .CO(\CARRYB[35][16] ), .S(\SUMB[35][16] ) );
  FA1P S2_30_23 ( .A(\CARRYB[29][23] ), .B(\ab[30][23] ), .CI(\SUMB[29][24] ), 
        .CO(\CARRYB[30][23] ), .S(\SUMB[30][23] ) );
  FA1P S2_10_44 ( .A(\ab[44][10] ), .B(\CARRYB[9][44] ), .CI(\SUMB[9][45] ), 
        .CO(\CARRYB[10][44] ), .S(\SUMB[10][44] ) );
  FA1P S2_11_44 ( .A(\ab[44][11] ), .B(\CARRYB[10][44] ), .CI(\SUMB[10][45] ), 
        .CO(\CARRYB[11][44] ), .S(\SUMB[11][44] ) );
  FA1P S2_8_34 ( .A(\CARRYB[7][34] ), .B(n522), .CI(\SUMB[7][35] ), .CO(
        \CARRYB[8][34] ), .S(\SUMB[8][34] ) );
  FA1P S2_15_11 ( .A(\CARRYB[14][11] ), .B(n626), .CI(\SUMB[14][12] ), .CO(
        \CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA1AP S2_14_41 ( .A(\CARRYB[13][41] ), .B(\ab[41][14] ), .CI(\SUMB[13][42] ), 
        .CO(\CARRYB[14][41] ), .S(\SUMB[14][41] ) );
  FA1P S2_28_15 ( .A(\CARRYB[27][15] ), .B(n721), .CI(\SUMB[27][16] ), .CO(
        \CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA1A S2_44_21 ( .A(\CARRYB[43][21] ), .B(\ab[44][21] ), .CI(\SUMB[43][22] ), 
        .CO(\CARRYB[44][21] ), .S(\SUMB[44][21] ) );
  FA1P S2_35_1 ( .A(n2188), .B(\CARRYB[34][1] ), .CI(\SUMB[34][2] ), .CO(
        \CARRYB[35][1] ), .S(\SUMB[35][1] ) );
  FA1P S2_43_1 ( .A(n2202), .B(\CARRYB[42][1] ), .CI(\SUMB[42][2] ), .CO(
        \CARRYB[43][1] ), .S(\SUMB[43][1] ) );
  FA1P S2_22_29 ( .A(\ab[29][22] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA1P S2_26_39 ( .A(\ab[39][26] ), .B(\CARRYB[25][39] ), .CI(\SUMB[25][40] ), 
        .CO(\CARRYB[26][39] ), .S(\SUMB[26][39] ) );
  FA1P S2_8_44 ( .A(n516), .B(\CARRYB[7][44] ), .CI(\SUMB[7][45] ), .CO(
        \CARRYB[8][44] ), .S(\SUMB[8][44] ) );
  FA1A S2_43_4 ( .A(\CARRYB[42][4] ), .B(n389), .CI(\SUMB[42][5] ), .CO(
        \CARRYB[43][4] ), .S(\SUMB[43][4] ) );
  FA1P S2_30_5 ( .A(n392), .B(\CARRYB[29][5] ), .CI(\SUMB[29][6] ), .CO(
        \CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA1P S2_31_2 ( .A(n2198), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), .CO(
        \CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FA1 S2_21_24 ( .A(\CARRYB[20][24] ), .B(\ab[24][21] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA1P S2_42_9 ( .A(\SUMB[41][10] ), .B(\CARRYB[41][9] ), .CI(n583), .CO(
        \CARRYB[42][9] ), .S(\SUMB[42][9] ) );
  FA1P S2_25_39 ( .A(\ab[39][25] ), .B(\CARRYB[24][39] ), .CI(\SUMB[24][40] ), 
        .CO(\CARRYB[25][39] ), .S(\SUMB[25][39] ) );
  FA1P S2_11_24 ( .A(\CARRYB[10][24] ), .B(n621), .CI(\SUMB[10][25] ), .CO(
        \CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1P S2_18_42 ( .A(\ab[42][18] ), .B(\CARRYB[17][42] ), .CI(\SUMB[17][43] ), 
        .CO(\CARRYB[18][42] ), .S(\SUMB[18][42] ) );
  FA1P S2_18_15 ( .A(n713), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), .CO(
        \CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA1P S2_19_15 ( .A(\CARRYB[18][15] ), .B(n725), .CI(\SUMB[18][16] ), .CO(
        \CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA1P S2_45_11 ( .A(\CARRYB[44][11] ), .B(\ab[45][11] ), .CI(\SUMB[44][12] ), 
        .CO(\CARRYB[45][11] ), .S(\SUMB[45][11] ) );
  FA1P S2_9_31 ( .A(n562), .B(\CARRYB[8][31] ), .CI(\SUMB[8][32] ), .CO(
        \CARRYB[9][31] ), .S(\SUMB[9][31] ) );
  FA1P S2_35_23 ( .A(\ab[35][23] ), .B(\CARRYB[34][23] ), .CI(\SUMB[34][24] ), 
        .CO(\CARRYB[35][23] ), .S(\SUMB[35][23] ) );
  FA1P S2_30_7 ( .A(n489), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), .CO(
        \CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA1P S2_44_5 ( .A(n439), .B(\CARRYB[43][5] ), .CI(\SUMB[43][6] ), .CO(
        \CARRYB[44][5] ), .S(\SUMB[44][5] ) );
  FA1P S2_20_14 ( .A(n709), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), .CO(
        \CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA1P S2_21_14 ( .A(\CARRYB[20][14] ), .B(n704), .CI(\SUMB[20][15] ), .CO(
        \CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA1 S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA1P S2_4_14 ( .A(n385), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), .CO(
        \CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1P S2_5_14 ( .A(n417), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1 S2_39_24 ( .A(\ab[39][24] ), .B(\CARRYB[38][24] ), .CI(\SUMB[38][25] ), 
        .CO(\CARRYB[39][24] ), .S(\SUMB[39][24] ) );
  FA1P S2_23_13 ( .A(\SUMB[22][14] ), .B(\CARRYB[22][13] ), .CI(n684), .CO(
        \CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA1P S2_28_12 ( .A(\CARRYB[27][12] ), .B(n668), .CI(\SUMB[27][13] ), .CO(
        \CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA1P S2_30_15 ( .A(\ab[30][15] ), .B(\CARRYB[29][15] ), .CI(\SUMB[29][16] ), 
        .CO(\CARRYB[30][15] ), .S(\SUMB[30][15] ) );
  FA1P S2_6_23 ( .A(n438), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), .CO(
        \CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1P S2_45_19 ( .A(\ab[45][19] ), .B(\CARRYB[44][19] ), .CI(\SUMB[44][20] ), 
        .CO(\CARRYB[45][19] ), .S(\SUMB[45][19] ) );
  FA1P S2_14_11 ( .A(n625), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), .CO(
        \CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1P S2_9_9 ( .A(n2337), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1P S3_15_46 ( .A(\ab[46][15] ), .B(\CARRYB[14][46] ), .CI(\ab[47][14] ), 
        .CO(\CARRYB[15][46] ), .S(\SUMB[15][46] ) );
  FA1P S2_16_35 ( .A(\ab[35][16] ), .B(\CARRYB[15][35] ), .CI(\SUMB[15][36] ), 
        .CO(\CARRYB[16][35] ), .S(\SUMB[16][35] ) );
  FA1P S2_8_29 ( .A(\CARRYB[7][29] ), .B(n549), .CI(\SUMB[7][30] ), .CO(
        \CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1P S2_29_16 ( .A(\CARRYB[28][16] ), .B(\ab[29][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA1P S2_29_6 ( .A(n455), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), .CO(
        \CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA1P S2_21_37 ( .A(\ab[37][21] ), .B(\CARRYB[20][37] ), .CI(\SUMB[20][38] ), 
        .CO(\CARRYB[21][37] ), .S(\SUMB[21][37] ) );
  FA1P S2_35_19 ( .A(\ab[35][19] ), .B(\CARRYB[34][19] ), .CI(\SUMB[34][20] ), 
        .CO(\CARRYB[35][19] ), .S(\SUMB[35][19] ) );
  FA1A S2_46_27 ( .A(\ab[46][27] ), .B(\CARRYB[45][27] ), .CI(\SUMB[45][28] ), 
        .CO(\CARRYB[46][27] ), .S(\SUMB[46][27] ) );
  FA1P S2_42_14 ( .A(\SUMB[41][15] ), .B(\ab[42][14] ), .CI(\CARRYB[41][14] ), 
        .CO(\CARRYB[42][14] ), .S(\SUMB[42][14] ) );
  FA1P S2_16_10 ( .A(n607), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), .CO(
        \CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1P S2_16_5 ( .A(n400), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), .CO(
        \CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1A S2_27_30 ( .A(\CARRYB[26][30] ), .B(\ab[30][27] ), .CI(\SUMB[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA1P S2_32_30 ( .A(\ab[32][30] ), .B(\CARRYB[31][30] ), .CI(\SUMB[31][31] ), 
        .CO(\CARRYB[32][30] ), .S(\SUMB[32][30] ) );
  FA1P S2_20_19 ( .A(\CARRYB[19][19] ), .B(\ab[20][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA1 S2_32_16 ( .A(\ab[32][16] ), .B(\CARRYB[31][16] ), .CI(\SUMB[31][17] ), 
        .CO(\CARRYB[32][16] ), .S(\SUMB[32][16] ) );
  FA1P S2_31_5 ( .A(n416), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), .CO(
        \CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FA1P S2_10_40 ( .A(n637), .B(\CARRYB[9][40] ), .CI(\SUMB[9][41] ), .CO(
        \CARRYB[10][40] ), .S(\SUMB[10][40] ) );
  FA1P S2_10_25 ( .A(\CARRYB[9][25] ), .B(n591), .CI(\SUMB[9][26] ), .CO(
        \CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1 S2_19_13 ( .A(n679), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), .CO(
        \CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA1P S2_3_19 ( .A(\CARRYB[2][19] ), .B(n2272), .CI(\SUMB[2][20] ), .CO(
        \CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1 S2_10_16 ( .A(\CARRYB[9][16] ), .B(n607), .CI(\SUMB[9][17] ), .CO(
        \CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1P S2_11_30 ( .A(n623), .B(\CARRYB[10][30] ), .CI(\SUMB[10][31] ), .CO(
        \CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA1P S2_7_43 ( .A(\CARRYB[6][43] ), .B(n474), .CI(\SUMB[6][44] ), .CO(
        \CARRYB[7][43] ), .S(\SUMB[7][43] ) );
  FA1 S2_41_37 ( .A(\ab[41][37] ), .B(\CARRYB[40][37] ), .CI(\SUMB[40][38] ), 
        .CO(\CARRYB[41][37] ), .S(\SUMB[41][37] ) );
  FA1P S2_11_43 ( .A(\ab[43][11] ), .B(\CARRYB[10][43] ), .CI(\SUMB[10][44] ), 
        .CO(\CARRYB[11][43] ), .S(\SUMB[11][43] ) );
  FA1P S2_12_43 ( .A(\ab[43][12] ), .B(\CARRYB[11][43] ), .CI(\SUMB[11][44] ), 
        .CO(\CARRYB[12][43] ), .S(\SUMB[12][43] ) );
  FA1P S2_22_42 ( .A(\ab[42][22] ), .B(\CARRYB[21][42] ), .CI(\SUMB[21][43] ), 
        .CO(\CARRYB[22][42] ), .S(\SUMB[22][42] ) );
  FA1P S2_23_42 ( .A(\ab[42][23] ), .B(\CARRYB[22][42] ), .CI(\SUMB[22][43] ), 
        .CO(\CARRYB[23][42] ), .S(\SUMB[23][42] ) );
  FA1P S2_45_33 ( .A(\ab[45][33] ), .B(\CARRYB[44][33] ), .CI(\SUMB[44][34] ), 
        .CO(\CARRYB[45][33] ), .S(\SUMB[45][33] ) );
  FA1P S2_15_10 ( .A(n588), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), .CO(
        \CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1P S2_33_39 ( .A(\ab[39][33] ), .B(\CARRYB[32][39] ), .CI(\SUMB[32][40] ), 
        .CO(\CARRYB[33][39] ), .S(\SUMB[33][39] ) );
  FA1 S2_45_27 ( .A(\SUMB[44][28] ), .B(\CARRYB[44][27] ), .CI(\ab[45][27] ), 
        .CO(\CARRYB[45][27] ), .S(\SUMB[45][27] ) );
  FA1P S2_3_43 ( .A(\SUMB[2][44] ), .B(\CARRYB[2][43] ), .CI(n2297), .CO(
        \CARRYB[3][43] ), .S(\SUMB[3][43] ) );
  FA1P S2_44_20 ( .A(\ab[44][20] ), .B(\CARRYB[43][20] ), .CI(\SUMB[43][21] ), 
        .CO(\CARRYB[44][20] ), .S(\SUMB[44][20] ) );
  FA1P S2_45_20 ( .A(\ab[45][20] ), .B(\CARRYB[44][20] ), .CI(\SUMB[44][21] ), 
        .CO(\CARRYB[45][20] ), .S(\SUMB[45][20] ) );
  FA1P S2_34_29 ( .A(\ab[34][29] ), .B(\CARRYB[33][29] ), .CI(\SUMB[33][30] ), 
        .CO(\CARRYB[34][29] ), .S(\SUMB[34][29] ) );
  FA1P S2_17_7 ( .A(n488), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), .CO(
        \CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1P S2_21_27 ( .A(\CARRYB[20][27] ), .B(\ab[27][21] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA1P S2_38_37 ( .A(\ab[38][37] ), .B(\CARRYB[37][37] ), .CI(\SUMB[37][38] ), 
        .CO(\CARRYB[38][37] ), .S(\SUMB[38][37] ) );
  FA1AP S2_26_29 ( .A(\ab[29][26] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA1P S2_4_37 ( .A(\CARRYB[3][37] ), .B(n361), .CI(\SUMB[3][38] ), .CO(
        \CARRYB[4][37] ), .S(\SUMB[4][37] ) );
  FA1A S2_35_28 ( .A(\ab[35][28] ), .B(\CARRYB[34][28] ), .CI(\SUMB[34][29] ), 
        .CO(\CARRYB[35][28] ), .S(\SUMB[35][28] ) );
  FA1P S2_19_20 ( .A(\CARRYB[18][20] ), .B(\ab[20][19] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA1P S2_9_24 ( .A(n571), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), .CO(
        \CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1P S2_10_24 ( .A(\CARRYB[9][24] ), .B(n597), .CI(\SUMB[9][25] ), .CO(
        \CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1 S2_46_17 ( .A(\ab[46][17] ), .B(\CARRYB[45][17] ), .CI(\SUMB[45][18] ), 
        .CO(\CARRYB[46][17] ), .S(\SUMB[46][17] ) );
  FA1P S2_32_39 ( .A(\ab[39][32] ), .B(\CARRYB[31][39] ), .CI(\SUMB[31][40] ), 
        .CO(\CARRYB[32][39] ), .S(\SUMB[32][39] ) );
  FA1 S2_34_28 ( .A(\SUMB[33][29] ), .B(\CARRYB[33][28] ), .CI(\ab[34][28] ), 
        .CO(\CARRYB[34][28] ), .S(\SUMB[34][28] ) );
  FA1A S2_18_35 ( .A(\ab[35][18] ), .B(\CARRYB[17][35] ), .CI(\SUMB[17][36] ), 
        .CO(\CARRYB[18][35] ), .S(\SUMB[18][35] ) );
  FA1A S2_4_18 ( .A(\CARRYB[3][18] ), .B(n2308), .CI(\SUMB[3][19] ), .CO(
        \CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1P S2_8_25 ( .A(\CARRYB[7][25] ), .B(n538), .CI(\SUMB[7][26] ), .CO(
        \CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1P S2_35_4 ( .A(n363), .B(\CARRYB[34][4] ), .CI(\SUMB[34][5] ), .CO(
        \CARRYB[35][4] ), .S(\SUMB[35][4] ) );
  FA1P S2_9_5 ( .A(n437), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1P S2_5_32 ( .A(n407), .B(\CARRYB[4][32] ), .CI(\SUMB[4][33] ), .CO(
        \CARRYB[5][32] ), .S(\SUMB[5][32] ) );
  FA1AP S2_3_31 ( .A(\CARRYB[2][31] ), .B(n2268), .CI(\SUMB[2][32] ), .CO(
        \CARRYB[3][31] ), .S(\SUMB[3][31] ) );
  FA1P S2_9_19 ( .A(\CARRYB[8][19] ), .B(n556), .CI(\SUMB[8][20] ), .CO(
        \CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1P S2_3_14 ( .A(n341), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), .CO(
        \CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1AP S2_21_31 ( .A(\ab[31][21] ), .B(\CARRYB[20][31] ), .CI(\SUMB[20][32] ), 
        .CO(\CARRYB[21][31] ), .S(\SUMB[21][31] ) );
  FA1P S2_5_26 ( .A(n410), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), .CO(
        \CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1P S2_3_27 ( .A(\CARRYB[2][27] ), .B(n2274), .CI(\SUMB[2][28] ), .CO(
        \CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1P S2_9_25 ( .A(\CARRYB[8][25] ), .B(n557), .CI(\SUMB[8][26] ), .CO(
        \CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1P S2_21_13 ( .A(n696), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), .CO(
        \CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA1A S2_36_45 ( .A(\ab[45][36] ), .B(\CARRYB[35][45] ), .CI(\SUMB[35][46] ), 
        .CO(\CARRYB[36][45] ), .S(\SUMB[36][45] ) );
  FA1A S2_46_44 ( .A(\ab[46][44] ), .B(\CARRYB[45][44] ), .CI(\SUMB[45][45] ), 
        .CO(\CARRYB[46][44] ), .S(\SUMB[46][44] ) );
  FA1P S3_14_46 ( .A(\ab[46][14] ), .B(\CARRYB[13][46] ), .CI(\ab[47][13] ), 
        .CO(\CARRYB[14][46] ), .S(\SUMB[14][46] ) );
  FA1P S3_10_46 ( .A(\ab[46][10] ), .B(\CARRYB[9][46] ), .CI(\ab[9][47] ), 
        .CO(\CARRYB[10][46] ), .S(\SUMB[10][46] ) );
  FA1A S2_2_11 ( .A(n335), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), .CO(
        \CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1 S2_46_20 ( .A(\ab[46][20] ), .B(\CARRYB[45][20] ), .CI(\SUMB[45][21] ), 
        .CO(\CARRYB[46][20] ), .S(\SUMB[46][20] ) );
  FA1P S2_45_4 ( .A(\CARRYB[44][4] ), .B(n360), .CI(\SUMB[44][5] ), .CO(
        \CARRYB[45][4] ), .S(\SUMB[45][4] ) );
  FA1P S2_33_24 ( .A(\ab[33][24] ), .B(\CARRYB[32][24] ), .CI(\SUMB[32][25] ), 
        .CO(\CARRYB[33][24] ), .S(\SUMB[33][24] ) );
  FA1P S2_40_8 ( .A(n545), .B(\CARRYB[39][8] ), .CI(\SUMB[39][9] ), .CO(
        \CARRYB[40][8] ), .S(\SUMB[40][8] ) );
  FA1P S2_2_36 ( .A(n2260), .B(\CARRYB[1][36] ), .CI(\SUMB[1][37] ), .CO(
        \CARRYB[2][36] ), .S(\SUMB[2][36] ) );
  FA1P S2_44_34 ( .A(\ab[44][34] ), .B(\CARRYB[43][34] ), .CI(\SUMB[43][35] ), 
        .CO(\CARRYB[44][34] ), .S(\SUMB[44][34] ) );
  FA1AP S2_8_35 ( .A(n507), .B(\CARRYB[7][35] ), .CI(\SUMB[7][36] ), .CO(
        \CARRYB[8][35] ), .S(\SUMB[8][35] ) );
  FA1A S2_42_19 ( .A(\CARRYB[41][19] ), .B(\ab[42][19] ), .CI(\SUMB[41][20] ), 
        .CO(\CARRYB[42][19] ), .S(\SUMB[42][19] ) );
  FA1A S1_2_0 ( .A(n2428), .B(\ab[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S2_2_1 ( .A(n2430), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_2_2 ( .A(n2319), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S2_4_4 ( .A(n2329), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_7_7 ( .A(n2335), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S1_3_0 ( .A(n2425), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S3_42_46 ( .A(\ab[46][42] ), .B(\CARRYB[41][46] ), .CI(\ab[47][41] ), 
        .CO(\CARRYB[42][46] ), .S(\SUMB[42][46] ) );
  FA1A S3_40_46 ( .A(\ab[46][40] ), .B(\CARRYB[39][46] ), .CI(\ab[47][39] ), 
        .CO(\CARRYB[40][46] ), .S(\SUMB[40][46] ) );
  FA1A S3_39_46 ( .A(\ab[46][39] ), .B(\CARRYB[38][46] ), .CI(\ab[47][38] ), 
        .CO(\CARRYB[39][46] ), .S(\SUMB[39][46] ) );
  FA1A S3_44_46 ( .A(\ab[46][44] ), .B(\CARRYB[43][46] ), .CI(\ab[47][43] ), 
        .CO(\CARRYB[44][46] ), .S(\SUMB[44][46] ) );
  FA1A S2_37_42 ( .A(\ab[42][37] ), .B(\CARRYB[36][42] ), .CI(\SUMB[36][43] ), 
        .CO(\CARRYB[37][42] ), .S(\SUMB[37][42] ) );
  FA1A S2_43_40 ( .A(\ab[43][40] ), .B(\CARRYB[42][40] ), .CI(\SUMB[42][41] ), 
        .CO(\CARRYB[43][40] ), .S(\SUMB[43][40] ) );
  FA1A S2_38_42 ( .A(\ab[42][38] ), .B(\CARRYB[37][42] ), .CI(\SUMB[37][43] ), 
        .CO(\CARRYB[38][42] ), .S(\SUMB[38][42] ) );
  FA1A S2_36_43 ( .A(\ab[43][36] ), .B(\CARRYB[35][43] ), .CI(\SUMB[35][44] ), 
        .CO(\CARRYB[36][43] ), .S(\SUMB[36][43] ) );
  FA1A S2_44_40 ( .A(\ab[44][40] ), .B(\CARRYB[43][40] ), .CI(\SUMB[43][41] ), 
        .CO(\CARRYB[44][40] ), .S(\SUMB[44][40] ) );
  FA1A S3_34_46 ( .A(\ab[46][34] ), .B(\CARRYB[33][46] ), .CI(\ab[47][33] ), 
        .CO(\CARRYB[34][46] ), .S(\SUMB[34][46] ) );
  FA1A S2_3_4 ( .A(n344), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_11_2 ( .A(n335), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(
        \CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_6_4 ( .A(n393), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_43_45 ( .A(\ab[45][43] ), .B(\CARRYB[42][45] ), .CI(\SUMB[42][46] ), 
        .CO(\CARRYB[43][45] ), .S(\SUMB[43][45] ) );
  FA1A S2_40_45 ( .A(\ab[45][40] ), .B(\CARRYB[39][45] ), .CI(\SUMB[39][46] ), 
        .CO(\CARRYB[40][45] ), .S(\SUMB[40][45] ) );
  FA1A S2_39_45 ( .A(\ab[45][39] ), .B(\CARRYB[38][45] ), .CI(\SUMB[38][46] ), 
        .CO(\CARRYB[39][45] ), .S(\SUMB[39][45] ) );
  FA1A S2_6_2 ( .A(n343), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_8_4 ( .A(n391), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_5_7 ( .A(n304), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_15_2 ( .A(n324), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_10_6 ( .A(n496), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_37_41 ( .A(\ab[41][37] ), .B(\CARRYB[36][41] ), .CI(\SUMB[36][42] ), 
        .CO(\CARRYB[37][41] ), .S(\SUMB[37][41] ) );
  FA1A S2_2_5 ( .A(n2267), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_4_5 ( .A(n390), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_13_1 ( .A(n2194), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), .CO(
        \CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_21_1 ( .A(n2179), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), .CO(
        \CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_5_8 ( .A(n419), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_45_44 ( .A(\ab[45][44] ), .B(\CARRYB[44][44] ), .CI(\SUMB[44][45] ), 
        .CO(\CARRYB[45][44] ), .S(\SUMB[45][44] ) );
  FA1A S2_33_45 ( .A(\ab[45][33] ), .B(\CARRYB[32][45] ), .CI(\SUMB[32][46] ), 
        .CO(\CARRYB[33][45] ), .S(\SUMB[33][45] ) );
  FA1AP S4_24 ( .A(\CARRYB[46][24] ), .B(\ab[47][24] ), .CI(\SUMB[46][25] ), 
        .CO(\CARRYB[47][24] ), .S(\SUMB[47][24] ) );
  FA1AP S4_9 ( .A(\CARRYB[46][9] ), .B(\ab[9][47] ), .CI(\SUMB[46][10] ), .CO(
        \CARRYB[47][9] ), .S(\SUMB[47][9] ) );
  FA1A S2_6_5 ( .A(n448), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_10_8 ( .A(n577), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_26_2 ( .A(n2258), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), .CO(
        \CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA1A S2_31_44 ( .A(\ab[44][31] ), .B(\CARRYB[30][44] ), .CI(\SUMB[30][45] ), 
        .CO(\CARRYB[31][44] ), .S(\SUMB[31][44] ) );
  FA1A S2_34_44 ( .A(\ab[44][34] ), .B(\CARRYB[33][44] ), .CI(\SUMB[33][45] ), 
        .CO(\CARRYB[34][44] ), .S(\SUMB[34][44] ) );
  FA1A S2_42_34 ( .A(\ab[42][34] ), .B(\CARRYB[41][34] ), .CI(\SUMB[41][35] ), 
        .CO(\CARRYB[42][34] ), .S(\SUMB[42][34] ) );
  FA1A S2_46_9 ( .A(\CARRYB[45][9] ), .B(\ab[9][46] ), .CI(\SUMB[45][10] ), 
        .CO(\CARRYB[46][9] ), .S(\SUMB[46][9] ) );
  FA1A S2_7_3 ( .A(n352), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_28_2 ( .A(n2210), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), .CO(
        \CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA1AP S2_19_39 ( .A(\ab[39][19] ), .B(\CARRYB[18][39] ), .CI(\SUMB[18][40] ), 
        .CO(\CARRYB[19][39] ), .S(\SUMB[19][39] ) );
  FA1A S2_36_44 ( .A(\ab[44][36] ), .B(\CARRYB[35][44] ), .CI(\SUMB[35][45] ), 
        .CO(\CARRYB[36][44] ), .S(\SUMB[36][44] ) );
  FA1A S2_35_45 ( .A(\ab[45][35] ), .B(\CARRYB[34][45] ), .CI(\SUMB[34][46] ), 
        .CO(\CARRYB[35][45] ), .S(\SUMB[35][45] ) );
  FA1A S1_23_0 ( .A(n2227), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), .CO(
        \CARRYB[23][0] ), .S(\A1[21] ) );
  FA1A S1_8_0 ( .A(n327), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_5_0 ( .A(n2256), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_4_0 ( .A(n326), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S2_3_11 ( .A(n354), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), .CO(
        \CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_16_8 ( .A(n525), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), .CO(
        \CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1A S2_22_11 ( .A(\CARRYB[21][11] ), .B(n641), .CI(\SUMB[21][12] ), .CO(
        \CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA1AP S4_6 ( .A(n487), .B(\CARRYB[46][6] ), .CI(\SUMB[46][7] ), .CO(
        \CARRYB[47][6] ), .S(\SUMB[47][6] ) );
  FA1A S2_11_9 ( .A(n594), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), .CO(
        \CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_14_9 ( .A(n576), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), .CO(
        \CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_44_22 ( .A(\ab[44][22] ), .B(\CARRYB[43][22] ), .CI(\SUMB[43][23] ), 
        .CO(\CARRYB[44][22] ), .S(\SUMB[44][22] ) );
  FA1A S2_27_10 ( .A(n611), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), .CO(
        \CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA1A S1_17_0 ( .A(n2193), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), .CO(
        \CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S1_11_0 ( .A(n289), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(
        \CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S2_21_10 ( .A(\CARRYB[20][10] ), .B(n616), .CI(\SUMB[20][11] ), .CO(
        \CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1AP S4_21 ( .A(\ab[47][21] ), .B(\CARRYB[46][21] ), .CI(\SUMB[46][22] ), 
        .CO(\CARRYB[47][21] ), .S(\SUMB[47][21] ) );
  FA1AP S4_16 ( .A(\ab[47][16] ), .B(\CARRYB[46][16] ), .CI(\SUMB[46][17] ), 
        .CO(\CARRYB[47][16] ), .S(\SUMB[47][16] ) );
  FA1AP S4_3 ( .A(\CARRYB[46][3] ), .B(n368), .CI(\SUMB[46][4] ), .CO(
        \CARRYB[47][3] ), .S(\SUMB[47][3] ) );
  FA1AP S4_4 ( .A(\CARRYB[46][4] ), .B(n406), .CI(\SUMB[46][5] ), .CO(
        \CARRYB[47][4] ), .S(\SUMB[47][4] ) );
  FA1A S1_21_0 ( .A(n331), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), .CO(
        \CARRYB[21][0] ), .S(\A1[19] ) );
  FA1A S2_6_6 ( .A(n2333), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_4_6 ( .A(n393), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S4_30 ( .A(\ab[47][30] ), .B(\CARRYB[46][30] ), .CI(\SUMB[46][31] ), 
        .CO(\CARRYB[47][30] ), .S(\SUMB[47][30] ) );
  FA1P S2_4_20 ( .A(n2302), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), .CO(
        \CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1P S2_45_34 ( .A(\ab[45][34] ), .B(\CARRYB[44][34] ), .CI(\SUMB[44][35] ), 
        .CO(\CARRYB[45][34] ), .S(\SUMB[45][34] ) );
  FA1AP S2_4_38 ( .A(n370), .B(\CARRYB[3][38] ), .CI(\SUMB[3][39] ), .CO(
        \CARRYB[4][38] ), .S(\SUMB[4][38] ) );
  FA1A S2_24_19 ( .A(\CARRYB[23][19] ), .B(\ab[24][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA1 S2_46_13 ( .A(\ab[46][13] ), .B(\CARRYB[45][13] ), .CI(\SUMB[45][14] ), 
        .CO(\CARRYB[46][13] ), .S(\SUMB[46][13] ) );
  FA1P S2_34_23 ( .A(\ab[34][23] ), .B(\CARRYB[33][23] ), .CI(\SUMB[33][24] ), 
        .CO(\CARRYB[34][23] ), .S(\SUMB[34][23] ) );
  FA1 S2_6_14 ( .A(\CARRYB[5][14] ), .B(n452), .CI(\SUMB[5][15] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1P S2_6_43 ( .A(\CARRYB[5][43] ), .B(n473), .CI(\SUMB[5][44] ), .CO(
        \CARRYB[6][43] ), .S(\SUMB[6][43] ) );
  FA1 S2_2_4 ( .A(n323), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1P S2_10_12 ( .A(\CARRYB[9][12] ), .B(n615), .CI(\SUMB[9][13] ), .CO(
        \CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1P S3_7_46 ( .A(n306), .B(\CARRYB[6][46] ), .CI(n487), .CO(\CARRYB[7][46] ), .S(\SUMB[7][46] ) );
  FA1P S2_16_2 ( .A(n319), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), .CO(
        \CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1 S2_10_9 ( .A(n587), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1 S2_38_3 ( .A(n2294), .B(\CARRYB[37][3] ), .CI(\SUMB[37][4] ), .CO(
        \CARRYB[38][3] ), .S(\SUMB[38][3] ) );
  FA1 S2_5_9 ( .A(n437), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1 S2_29_9 ( .A(n575), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), .CO(
        \CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA1P S2_17_6 ( .A(n436), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), .CO(
        \CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1P S2_34_4 ( .A(n2303), .B(\CARRYB[33][4] ), .CI(\SUMB[33][5] ), .CO(
        \CARRYB[34][4] ), .S(\SUMB[34][4] ) );
  FA1P S2_12_3 ( .A(n351), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), .CO(
        \CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1AP S4_8 ( .A(\ab[8][47] ), .B(\CARRYB[46][8] ), .CI(\SUMB[46][9] ), .CO(
        \CARRYB[47][8] ), .S(\SUMB[47][8] ) );
  FA1A S2_3_3 ( .A(n2327), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1AP S4_28 ( .A(\CARRYB[46][28] ), .B(\ab[47][28] ), .CI(\SUMB[46][29] ), 
        .CO(\CARRYB[47][28] ), .S(\SUMB[47][28] ) );
  FA1A S2_44_45 ( .A(\ab[45][44] ), .B(\CARRYB[43][45] ), .CI(\SUMB[43][46] ), 
        .CO(\CARRYB[44][45] ), .S(\SUMB[44][45] ) );
  FA1AP S4_18 ( .A(\ab[47][18] ), .B(\CARRYB[46][18] ), .CI(\SUMB[46][19] ), 
        .CO(\CARRYB[47][18] ), .S(\SUMB[47][18] ) );
  FA1P S2_4_26 ( .A(n362), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), .CO(
        \CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1P S2_37_15 ( .A(\ab[37][15] ), .B(\CARRYB[36][15] ), .CI(\SUMB[36][16] ), 
        .CO(\CARRYB[37][15] ), .S(\SUMB[37][15] ) );
  FA1 S2_8_13 ( .A(n544), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), .CO(
        \CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_5_13 ( .A(n422), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), .CO(
        \CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1P S2_2_17 ( .A(n2262), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), .CO(
        \CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1P S2_14_4 ( .A(n385), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(
        \CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_4_2 ( .A(n323), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S3_33_46 ( .A(\ab[46][33] ), .B(\CARRYB[32][46] ), .CI(\ab[47][32] ), 
        .CO(\CARRYB[33][46] ), .S(\SUMB[33][46] ) );
  FA1A S2_11_6 ( .A(n491), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(
        \CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1 S2_7_10 ( .A(n528), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), .CO(
        \CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_6_10 ( .A(n496), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), .CO(
        \CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1 S2_14_2 ( .A(n284), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), .CO(
        \CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1 S2_12_2 ( .A(n287), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), .CO(
        \CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1P S2_11_3 ( .A(n354), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(
        \CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_9_1 ( .A(n2217), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1P S2_4_12 ( .A(n386), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), .CO(
        \CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1P S2_5_12 ( .A(n405), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), .CO(
        \CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_3_6 ( .A(n357), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1P S2_6_11 ( .A(n491), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), .CO(
        \CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1 S2_2_6 ( .A(n343), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_39_38 ( .A(\ab[39][38] ), .B(\CARRYB[38][38] ), .CI(\SUMB[38][39] ), 
        .CO(\CARRYB[39][38] ), .S(\SUMB[39][38] ) );
  FA1P S2_8_10 ( .A(n577), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), .CO(
        \CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1AP S2_9_12 ( .A(\CARRYB[8][12] ), .B(n566), .CI(\SUMB[8][13] ), .CO(
        \CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1P S2_6_9 ( .A(n484), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_4_7 ( .A(n369), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1 S2_17_8 ( .A(n517), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), .CO(
        \CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1 S2_6_8 ( .A(n483), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1 S2_15_8 ( .A(n527), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1 S2_13_8 ( .A(n544), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), .CO(
        \CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1P S2_36_3 ( .A(n2277), .B(\CARRYB[35][3] ), .CI(\SUMB[35][4] ), .CO(
        \CARRYB[36][3] ), .S(\SUMB[36][3] ) );
  FA1P S2_41_9 ( .A(n612), .B(\CARRYB[40][9] ), .CI(\SUMB[40][10] ), .CO(
        \CARRYB[41][9] ), .S(\SUMB[41][9] ) );
  FA1AP S2_2_14 ( .A(\CARRYB[1][14] ), .B(n284), .CI(\SUMB[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1P S2_30_4 ( .A(n2281), .B(\CARRYB[29][4] ), .CI(\SUMB[29][5] ), .CO(
        \CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA1P S2_20_9 ( .A(n535), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), .CO(
        \CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1P S2_8_24 ( .A(n534), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), .CO(
        \CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1AP S2_23_11 ( .A(\CARRYB[22][11] ), .B(n642), .CI(\SUMB[22][12] ), .CO(
        \CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA1P S2_41_7 ( .A(\CARRYB[40][7] ), .B(n499), .CI(\SUMB[40][8] ), .CO(
        \CARRYB[41][7] ), .S(\SUMB[41][7] ) );
  FA1P S2_42_6 ( .A(\CARRYB[41][6] ), .B(n478), .CI(\SUMB[41][7] ), .CO(
        \CARRYB[42][6] ), .S(\SUMB[42][6] ) );
  FA1P S2_43_6 ( .A(\CARRYB[42][6] ), .B(n473), .CI(\SUMB[42][7] ), .CO(
        \CARRYB[43][6] ), .S(\SUMB[43][6] ) );
  FA1P S1_41_0 ( .A(n2239), .B(\CARRYB[40][0] ), .CI(\SUMB[40][1] ), .CO(
        \CARRYB[41][0] ), .S(\A1[39] ) );
  FA1P S2_32_6 ( .A(n435), .B(\CARRYB[31][6] ), .CI(\SUMB[31][7] ), .CO(
        \CARRYB[32][6] ), .S(\SUMB[32][6] ) );
  FA1P S2_32_2 ( .A(n2211), .B(\CARRYB[31][2] ), .CI(\SUMB[31][3] ), .CO(
        \CARRYB[32][2] ), .S(\SUMB[32][2] ) );
  FA1P S2_21_7 ( .A(n477), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), .CO(
        \CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA1P S2_21_9 ( .A(n561), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), .CO(
        \CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1P S2_27_40 ( .A(\ab[40][27] ), .B(\CARRYB[26][40] ), .CI(\SUMB[26][41] ), 
        .CO(\CARRYB[27][40] ), .S(\SUMB[27][40] ) );
  FA1 S2_26_10 ( .A(n604), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), .CO(
        \CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA1P S2_34_38 ( .A(\ab[38][34] ), .B(\CARRYB[33][38] ), .CI(\SUMB[33][39] ), 
        .CO(\CARRYB[34][38] ), .S(\SUMB[34][38] ) );
  FA1P S2_35_38 ( .A(\ab[38][35] ), .B(\CARRYB[34][38] ), .CI(\SUMB[34][39] ), 
        .CO(\CARRYB[35][38] ), .S(\SUMB[35][38] ) );
  FA1AP S2_25_11 ( .A(n633), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), .CO(
        \CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA1P S2_27_5 ( .A(n381), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), .CO(
        \CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA1P S2_2_15 ( .A(n324), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1P S2_12_22 ( .A(\CARRYB[11][22] ), .B(n678), .CI(\SUMB[11][23] ), .CO(
        \CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA1P S2_13_22 ( .A(n681), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), .CO(
        \CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA1P S2_3_15 ( .A(n340), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), .CO(
        \CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1P S2_23_6 ( .A(n438), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), .CO(
        \CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA1A S2_42_24 ( .A(\CARRYB[41][24] ), .B(\ab[42][24] ), .CI(\SUMB[41][25] ), 
        .CO(\CARRYB[42][24] ), .S(\SUMB[42][24] ) );
  FA1A S2_8_27 ( .A(\CARRYB[7][27] ), .B(n524), .CI(\SUMB[7][28] ), .CO(
        \CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1P S2_12_44 ( .A(\ab[44][12] ), .B(\CARRYB[11][44] ), .CI(\SUMB[11][45] ), 
        .CO(\CARRYB[12][44] ), .S(\SUMB[12][44] ) );
  FA1P S2_13_44 ( .A(\ab[44][13] ), .B(\CARRYB[12][44] ), .CI(\SUMB[12][45] ), 
        .CO(\CARRYB[13][44] ), .S(\SUMB[13][44] ) );
  FA1P S2_25_5 ( .A(n404), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), .CO(
        \CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA1P S3_8_46 ( .A(n503), .B(\CARRYB[7][46] ), .CI(\ab[7][47] ), .CO(
        \CARRYB[8][46] ), .S(\SUMB[8][46] ) );
  FA1P S3_9_46 ( .A(\ab[9][46] ), .B(\CARRYB[8][46] ), .CI(\ab[8][47] ), .CO(
        \CARRYB[9][46] ), .S(\SUMB[9][46] ) );
  FA1P S2_10_23 ( .A(n603), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), .CO(
        \CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA1P S2_3_35 ( .A(n2291), .B(\CARRYB[2][35] ), .CI(\SUMB[2][36] ), .CO(
        \CARRYB[3][35] ), .S(\SUMB[3][35] ) );
  FA1P S2_4_35 ( .A(n363), .B(\CARRYB[3][35] ), .CI(\SUMB[3][36] ), .CO(
        \CARRYB[4][35] ), .S(\SUMB[4][35] ) );
  FA1P S2_11_10 ( .A(n606), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), .CO(
        \CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1P S2_30_40 ( .A(\ab[40][30] ), .B(\CARRYB[29][40] ), .CI(\SUMB[29][41] ), 
        .CO(\CARRYB[30][40] ), .S(\SUMB[30][40] ) );
  FA1P S2_21_18 ( .A(\CARRYB[20][18] ), .B(\ab[21][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA1AP S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA1P S2_20_23 ( .A(\CARRYB[19][23] ), .B(\ab[23][20] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA1P S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA1A S2_4_13 ( .A(n372), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), .CO(
        \CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1 S2_26_9 ( .A(\CARRYB[25][9] ), .B(n564), .CI(\SUMB[25][10] ), .CO(
        \CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA1P S2_39_10 ( .A(n640), .B(\CARRYB[38][10] ), .CI(\SUMB[38][11] ), .CO(
        \CARRYB[39][10] ), .S(\SUMB[39][10] ) );
  FA1P S2_22_25 ( .A(\ab[25][22] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA1P S2_29_3 ( .A(n2270), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), .CO(
        \CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA1 S2_13_6 ( .A(n461), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), .CO(
        \CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1P S2_17_9 ( .A(n574), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), .CO(
        \CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1AP S2_19_43 ( .A(\ab[43][19] ), .B(\CARRYB[18][43] ), .CI(\SUMB[18][44] ), 
        .CO(\CARRYB[19][43] ), .S(\SUMB[19][43] ) );
  FA1 S2_3_42 ( .A(n2296), .B(\CARRYB[2][42] ), .CI(\SUMB[2][43] ), .CO(
        \CARRYB[3][42] ), .S(\SUMB[3][42] ) );
  FA1P S2_45_17 ( .A(\ab[45][17] ), .B(\CARRYB[44][17] ), .CI(\SUMB[44][18] ), 
        .CO(\CARRYB[45][17] ), .S(\SUMB[45][17] ) );
  FA1P S2_19_28 ( .A(\ab[28][19] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA1P S2_20_7 ( .A(n470), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), .CO(
        \CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1P S2_18_7 ( .A(n512), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), .CO(
        \CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1 S2_46_30 ( .A(\ab[46][30] ), .B(\CARRYB[45][30] ), .CI(\SUMB[45][31] ), 
        .CO(\CARRYB[46][30] ), .S(\SUMB[46][30] ) );
  FA1AP S2_46_26 ( .A(\ab[46][26] ), .B(\CARRYB[45][26] ), .CI(\SUMB[45][27] ), 
        .CO(\CARRYB[46][26] ), .S(\SUMB[46][26] ) );
  FA1P S2_3_36 ( .A(n2277), .B(\CARRYB[2][36] ), .CI(\SUMB[2][37] ), .CO(
        \CARRYB[3][36] ), .S(\SUMB[3][36] ) );
  FA1P S2_40_36 ( .A(\ab[40][36] ), .B(\CARRYB[39][36] ), .CI(\SUMB[39][37] ), 
        .CO(\CARRYB[40][36] ), .S(\SUMB[40][36] ) );
  FA1AP S2_45_22 ( .A(\ab[45][22] ), .B(\CARRYB[44][22] ), .CI(\SUMB[44][23] ), 
        .CO(\CARRYB[45][22] ), .S(\SUMB[45][22] ) );
  FA1P S2_38_33 ( .A(\ab[38][33] ), .B(\CARRYB[37][33] ), .CI(\SUMB[37][34] ), 
        .CO(\CARRYB[38][33] ), .S(\SUMB[38][33] ) );
  FA1P S2_36_34 ( .A(\ab[36][34] ), .B(\CARRYB[35][34] ), .CI(\SUMB[35][35] ), 
        .CO(\CARRYB[36][34] ), .S(\SUMB[36][34] ) );
  FA1 S2_44_14 ( .A(\ab[44][14] ), .B(\CARRYB[43][14] ), .CI(\SUMB[43][15] ), 
        .CO(\CARRYB[44][14] ), .S(\SUMB[44][14] ) );
  FA1P S2_20_30 ( .A(\ab[30][20] ), .B(\CARRYB[19][30] ), .CI(\SUMB[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA1P S2_9_10 ( .A(n587), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), .CO(
        \CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1P S2_2_23 ( .A(\CARRYB[1][23] ), .B(n2199), .CI(\SUMB[1][24] ), .CO(
        \CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1 S2_3_29 ( .A(\CARRYB[2][29] ), .B(n2270), .CI(\SUMB[2][30] ), .CO(
        \CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1 S2_21_12 ( .A(\CARRYB[20][12] ), .B(n667), .CI(\SUMB[20][13] ), .CO(
        \CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA1P S2_43_14 ( .A(\CARRYB[42][14] ), .B(\ab[43][14] ), .CI(\SUMB[42][15] ), 
        .CO(\CARRYB[43][14] ), .S(\SUMB[43][14] ) );
  FA1P S2_28_4 ( .A(n2307), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), .CO(
        \CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA1P S2_29_4 ( .A(n2299), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), .CO(
        \CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA1P S2_18_4 ( .A(n2308), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), .CO(
        \CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA1P S2_41_34 ( .A(\ab[41][34] ), .B(\CARRYB[40][34] ), .CI(\SUMB[40][35] ), 
        .CO(\CARRYB[41][34] ), .S(\SUMB[41][34] ) );
  FA1P S2_11_29 ( .A(n639), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), .CO(
        \CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1AP S2_43_16 ( .A(\ab[43][16] ), .B(\CARRYB[42][16] ), .CI(\SUMB[42][17] ), 
        .CO(\CARRYB[43][16] ), .S(\SUMB[43][16] ) );
  FA1AP S2_15_15 ( .A(n2349), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), .CO(
        \CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA1P S2_9_23 ( .A(\CARRYB[8][23] ), .B(n584), .CI(\SUMB[8][24] ), .CO(
        \CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1P S2_13_17 ( .A(n687), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), .CO(
        \CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA1P S2_12_17 ( .A(\CARRYB[11][17] ), .B(n677), .CI(\SUMB[11][18] ), .CO(
        \CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA1P S2_19_6 ( .A(n460), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), .CO(
        \CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1P S2_20_6 ( .A(n429), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), .CO(
        \CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1 S2_37_5 ( .A(n397), .B(\CARRYB[36][5] ), .CI(\SUMB[36][6] ), .CO(
        \CARRYB[37][5] ), .S(\SUMB[37][5] ) );
  FA1AP S2_21_34 ( .A(\CARRYB[20][34] ), .B(\ab[34][21] ), .CI(\SUMB[20][35] ), 
        .CO(\CARRYB[21][34] ), .S(\SUMB[21][34] ) );
  FA1P S2_4_33 ( .A(n2306), .B(\CARRYB[3][33] ), .CI(\SUMB[3][34] ), .CO(
        \CARRYB[4][33] ), .S(\SUMB[4][33] ) );
  FA1P S2_36_27 ( .A(\ab[36][27] ), .B(\CARRYB[35][27] ), .CI(\SUMB[35][28] ), 
        .CO(\CARRYB[36][27] ), .S(\SUMB[36][27] ) );
  FA1P S2_31_1 ( .A(n2185), .B(\CARRYB[30][1] ), .CI(\SUMB[30][2] ), .CO(
        \CARRYB[31][1] ), .S(\SUMB[31][1] ) );
  FA1P S2_32_1 ( .A(n2311), .B(\CARRYB[31][1] ), .CI(\SUMB[31][2] ), .CO(
        \CARRYB[32][1] ), .S(\SUMB[32][1] ) );
  FA1P S2_8_1 ( .A(n2232), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1P S2_8_43 ( .A(\CARRYB[7][43] ), .B(n520), .CI(\SUMB[7][44] ), .CO(
        \CARRYB[8][43] ), .S(\SUMB[8][43] ) );
  FA1P S2_31_29 ( .A(\ab[31][29] ), .B(\CARRYB[30][29] ), .CI(\SUMB[30][30] ), 
        .CO(\CARRYB[31][29] ), .S(\SUMB[31][29] ) );
  FA1A S2_23_1 ( .A(n2315), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), .CO(
        \CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA1 S2_43_22 ( .A(\ab[43][22] ), .B(\CARRYB[42][22] ), .CI(\SUMB[42][23] ), 
        .CO(\CARRYB[43][22] ), .S(\SUMB[43][22] ) );
  FA1P S2_32_22 ( .A(\CARRYB[31][22] ), .B(\ab[32][22] ), .CI(\SUMB[31][23] ), 
        .CO(\CARRYB[32][22] ), .S(\SUMB[32][22] ) );
  FA1A S2_32_7 ( .A(\CARRYB[31][7] ), .B(n476), .CI(\SUMB[31][8] ), .CO(
        \CARRYB[32][7] ), .S(\SUMB[32][7] ) );
  FA1AP S2_41_5 ( .A(n444), .B(\CARRYB[40][5] ), .CI(\SUMB[40][6] ), .CO(
        \CARRYB[41][5] ), .S(\SUMB[41][5] ) );
  FA1P S2_33_21 ( .A(\ab[33][21] ), .B(\CARRYB[32][21] ), .CI(\SUMB[32][22] ), 
        .CO(\CARRYB[33][21] ), .S(\SUMB[33][21] ) );
  FA1P S2_34_21 ( .A(\ab[34][21] ), .B(\CARRYB[33][21] ), .CI(\SUMB[33][22] ), 
        .CO(\CARRYB[34][21] ), .S(\SUMB[34][21] ) );
  FA1P S2_6_19 ( .A(n460), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), .CO(
        \CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1P S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA1P S2_5_34 ( .A(n403), .B(\CARRYB[4][34] ), .CI(\SUMB[4][35] ), .CO(
        \CARRYB[5][34] ), .S(\SUMB[5][34] ) );
  FA1P S2_19_38 ( .A(\ab[38][19] ), .B(\CARRYB[18][38] ), .CI(\SUMB[18][39] ), 
        .CO(\CARRYB[19][38] ), .S(\SUMB[19][38] ) );
  FA1 S2_20_38 ( .A(\ab[38][20] ), .B(\CARRYB[19][38] ), .CI(\SUMB[19][39] ), 
        .CO(\CARRYB[20][38] ), .S(\SUMB[20][38] ) );
  FA1P S2_2_27 ( .A(\CARRYB[1][27] ), .B(n2209), .CI(\SUMB[1][28] ), .CO(
        \CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1AP S2_27_9 ( .A(\CARRYB[26][9] ), .B(n573), .CI(\SUMB[26][10] ), .CO(
        \CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA1P S2_17_42 ( .A(\ab[42][17] ), .B(\CARRYB[16][42] ), .CI(\SUMB[16][43] ), 
        .CO(\CARRYB[17][42] ), .S(\SUMB[17][42] ) );
  FA1P S2_33_38 ( .A(\ab[38][33] ), .B(\CARRYB[32][38] ), .CI(\SUMB[32][39] ), 
        .CO(\CARRYB[33][38] ), .S(\SUMB[33][38] ) );
  FA1 S2_37_37 ( .A(n2400), .B(\CARRYB[36][37] ), .CI(\SUMB[36][38] ), .CO(
        \CARRYB[37][37] ), .S(\SUMB[37][37] ) );
  FA1P S2_35_37 ( .A(\ab[37][35] ), .B(\CARRYB[34][37] ), .CI(\SUMB[34][38] ), 
        .CO(\CARRYB[35][37] ), .S(\SUMB[35][37] ) );
  FA1P S2_36_37 ( .A(\ab[37][36] ), .B(\CARRYB[35][37] ), .CI(\SUMB[35][38] ), 
        .CO(\CARRYB[36][37] ), .S(\SUMB[36][37] ) );
  FA1P S2_21_3 ( .A(n2293), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), .CO(
        \CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1P S2_22_3 ( .A(n2292), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), .CO(
        \CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA1P S2_28_3 ( .A(n2284), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), .CO(
        \CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA1P S2_40_2 ( .A(n2250), .B(\CARRYB[39][2] ), .CI(\SUMB[39][3] ), .CO(
        \CARRYB[40][2] ), .S(\SUMB[40][2] ) );
  FA1A S2_6_3 ( .A(n357), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1P S2_16_3 ( .A(n337), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), .CO(
        \CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1 S2_3_23 ( .A(\CARRYB[2][23] ), .B(n2271), .CI(\SUMB[2][24] ), .CO(
        \CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA1P S2_5_20 ( .A(n402), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), .CO(
        \CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1P S2_13_29 ( .A(n689), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), .CO(
        \CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA1 S2_41_23 ( .A(\SUMB[40][24] ), .B(\CARRYB[40][23] ), .CI(\ab[41][23] ), 
        .CO(\CARRYB[41][23] ), .S(\SUMB[41][23] ) );
  FA1P S2_2_38 ( .A(\CARRYB[1][38] ), .B(n2249), .CI(\SUMB[1][39] ), .CO(
        \CARRYB[2][38] ), .S(\SUMB[2][38] ) );
  FA1P S2_4_21 ( .A(n366), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), .CO(
        \CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1AP S2_4_34 ( .A(n2303), .B(\CARRYB[3][34] ), .CI(\SUMB[3][35] ), .CO(
        \CARRYB[4][34] ), .S(\SUMB[4][34] ) );
  FA1P S2_18_31 ( .A(\ab[31][18] ), .B(\CARRYB[17][31] ), .CI(\SUMB[17][32] ), 
        .CO(\CARRYB[18][31] ), .S(\SUMB[18][31] ) );
  FA1AP S2_5_19 ( .A(n420), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), .CO(
        \CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1AP S2_5_18 ( .A(\CARRYB[4][18] ), .B(n415), .CI(\SUMB[4][19] ), .CO(
        \CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1P S2_19_14 ( .A(\CARRYB[18][14] ), .B(n699), .CI(\SUMB[18][15] ), .CO(
        \CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA1P S2_4_27 ( .A(n2309), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), .CO(
        \CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1P S2_20_11 ( .A(\CARRYB[19][11] ), .B(n627), .CI(\SUMB[19][12] ), .CO(
        \CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA1P S2_3_17 ( .A(n2279), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), .CO(
        \CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1P S2_4_17 ( .A(n371), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), .CO(
        \CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1P S2_39_31 ( .A(\ab[39][31] ), .B(\CARRYB[38][31] ), .CI(\SUMB[38][32] ), 
        .CO(\CARRYB[39][31] ), .S(\SUMB[39][31] ) );
  FA1AP S2_4_28 ( .A(\CARRYB[3][28] ), .B(n2307), .CI(\SUMB[3][29] ), .CO(
        \CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1A S2_29_8 ( .A(n549), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), .CO(
        \CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA1 S1_20_0 ( .A(n892), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), .CO(
        \CARRYB[20][0] ), .S(\A1[18] ) );
  FA1P S1_34_0 ( .A(n2189), .B(\CARRYB[33][0] ), .CI(\SUMB[33][1] ), .CO(
        \CARRYB[34][0] ), .S(\A1[32] ) );
  FA1P S2_34_30 ( .A(\ab[34][30] ), .B(\CARRYB[33][30] ), .CI(\SUMB[33][31] ), 
        .CO(\CARRYB[34][30] ), .S(\SUMB[34][30] ) );
  FA1A S2_29_13 ( .A(n689), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), .CO(
        \CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA1AP S2_25_15 ( .A(n723), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), .CO(
        \CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA1P S2_7_19 ( .A(n497), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), .CO(
        \CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S2_8_32 ( .A(n529), .B(\CARRYB[7][32] ), .CI(\SUMB[7][33] ), .CO(
        \CARRYB[8][32] ), .S(\SUMB[8][32] ) );
  FA1P S2_31_21 ( .A(\ab[31][21] ), .B(\CARRYB[30][21] ), .CI(\SUMB[30][22] ), 
        .CO(\CARRYB[31][21] ), .S(\SUMB[31][21] ) );
  FA1A S2_34_27 ( .A(\CARRYB[33][27] ), .B(\ab[34][27] ), .CI(\SUMB[33][28] ), 
        .CO(\CARRYB[34][27] ), .S(\SUMB[34][27] ) );
  FA1P S2_36_8 ( .A(n543), .B(\CARRYB[35][8] ), .CI(\SUMB[35][9] ), .CO(
        \CARRYB[36][8] ), .S(\SUMB[36][8] ) );
  FA1P S1_44_0 ( .A(n2204), .B(\CARRYB[43][0] ), .CI(\SUMB[43][1] ), .CO(
        \CARRYB[44][0] ), .S(\A1[42] ) );
  FA1P S1_45_0 ( .A(n2243), .B(\CARRYB[44][0] ), .CI(\SUMB[44][1] ), .CO(
        \CARRYB[45][0] ), .S(\A1[43] ) );
  FA1P S1_27_0 ( .A(n2224), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), .CO(
        \CARRYB[27][0] ), .S(\A1[25] ) );
  FA1P S1_33_0 ( .A(n2313), .B(\CARRYB[32][0] ), .CI(\SUMB[32][1] ), .CO(
        \CARRYB[33][0] ), .S(\A1[31] ) );
  FA1P S1_9_0 ( .A(n2229), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1 S1_10_0 ( .A(n2230), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1 S2_7_21 ( .A(\CARRYB[6][21] ), .B(n477), .CI(\SUMB[6][22] ), .CO(
        \CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA1P S2_31_23 ( .A(\ab[31][23] ), .B(\CARRYB[30][23] ), .CI(\SUMB[30][24] ), 
        .CO(\CARRYB[31][23] ), .S(\SUMB[31][23] ) );
  FA1P S2_32_23 ( .A(\CARRYB[31][23] ), .B(\ab[32][23] ), .CI(\SUMB[31][24] ), 
        .CO(\CARRYB[32][23] ), .S(\SUMB[32][23] ) );
  FA1 S2_24_16 ( .A(\CARRYB[23][16] ), .B(\ab[24][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA1A S2_30_13 ( .A(\CARRYB[29][13] ), .B(n692), .CI(\SUMB[29][14] ), .CO(
        \CARRYB[30][13] ), .S(\SUMB[30][13] ) );
  FA1AP S2_31_27 ( .A(\CARRYB[30][27] ), .B(\ab[31][27] ), .CI(\SUMB[30][28] ), 
        .CO(\CARRYB[31][27] ), .S(\SUMB[31][27] ) );
  FA1P S2_44_13 ( .A(\CARRYB[43][13] ), .B(\ab[44][13] ), .CI(\SUMB[43][14] ), 
        .CO(\CARRYB[44][13] ), .S(\SUMB[44][13] ) );
  FA1AP S2_20_12 ( .A(\CARRYB[19][12] ), .B(n665), .CI(\SUMB[19][13] ), .CO(
        \CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA1P S2_31_34 ( .A(\ab[34][31] ), .B(\CARRYB[30][34] ), .CI(\SUMB[30][35] ), 
        .CO(\CARRYB[31][34] ), .S(\SUMB[31][34] ) );
  FA1AP S2_11_15 ( .A(\CARRYB[10][15] ), .B(n626), .CI(\SUMB[10][16] ), .CO(
        \CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1 S2_23_19 ( .A(\CARRYB[22][19] ), .B(\ab[23][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA1P S2_29_12 ( .A(\CARRYB[28][12] ), .B(n676), .CI(\SUMB[28][13] ), .CO(
        \CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA1 S2_20_29 ( .A(\ab[29][20] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA1 S2_9_20 ( .A(\CARRYB[8][20] ), .B(n535), .CI(\SUMB[8][21] ), .CO(
        \CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1 S2_34_6 ( .A(n459), .B(\CARRYB[33][6] ), .CI(\SUMB[33][7] ), .CO(
        \CARRYB[34][6] ), .S(\SUMB[34][6] ) );
  FA1AP S2_40_25 ( .A(\ab[40][25] ), .B(\CARRYB[39][25] ), .CI(\SUMB[39][26] ), 
        .CO(\CARRYB[40][25] ), .S(\SUMB[40][25] ) );
  FA1P S2_14_28 ( .A(n706), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), .CO(
        \CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA1P S2_15_28 ( .A(n721), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), .CO(
        \CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA1A S2_17_13 ( .A(\CARRYB[16][13] ), .B(n687), .CI(\SUMB[16][14] ), .CO(
        \CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA1AP S2_35_22 ( .A(\CARRYB[34][22] ), .B(\ab[35][22] ), .CI(\SUMB[34][23] ), 
        .CO(\CARRYB[35][22] ), .S(\SUMB[35][22] ) );
  FA1P S2_36_5 ( .A(n399), .B(\CARRYB[35][5] ), .CI(\SUMB[35][6] ), .CO(
        \CARRYB[36][5] ), .S(\SUMB[36][5] ) );
  FA1P S2_12_24 ( .A(\CARRYB[11][24] ), .B(n660), .CI(\SUMB[11][25] ), .CO(
        \CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA1 S2_18_21 ( .A(\CARRYB[17][21] ), .B(\ab[21][18] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA1AP S2_13_35 ( .A(\CARRYB[12][35] ), .B(\ab[35][13] ), .CI(\SUMB[12][36] ), 
        .CO(\CARRYB[13][35] ), .S(\SUMB[13][35] ) );
  FA1AP S2_7_18 ( .A(n512), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), .CO(
        \CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1AP S2_18_17 ( .A(\CARRYB[17][17] ), .B(\ab[18][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA1 S2_3_39 ( .A(n2305), .B(\CARRYB[2][39] ), .CI(\SUMB[2][40] ), .CO(
        \CARRYB[3][39] ), .S(\SUMB[3][39] ) );
  FA1A S1_31_0 ( .A(n2170), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), .CO(
        \CARRYB[31][0] ), .S(\A1[29] ) );
  FA1AP S2_11_16 ( .A(n624), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), .CO(
        \CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1A S2_32_8 ( .A(n529), .B(\CARRYB[31][8] ), .CI(\SUMB[31][9] ), .CO(
        \CARRYB[32][8] ), .S(\SUMB[32][8] ) );
  FA1AP S2_23_12 ( .A(\CARRYB[22][12] ), .B(n666), .CI(\SUMB[22][13] ), .CO(
        \CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA1P S2_28_9 ( .A(n563), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), .CO(
        \CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA1AP S2_28_25 ( .A(\CARRYB[27][25] ), .B(\ab[28][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA1AP S2_6_33 ( .A(n433), .B(\CARRYB[5][33] ), .CI(\SUMB[5][34] ), .CO(
        \CARRYB[6][33] ), .S(\SUMB[6][33] ) );
  FA1AP S2_6_16 ( .A(n445), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), .CO(
        \CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1AP S2_28_21 ( .A(\CARRYB[27][21] ), .B(\ab[28][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA1AP S2_26_21 ( .A(\ab[26][21] ), .B(\CARRYB[25][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA1P S2_16_27 ( .A(\ab[27][16] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA1AP S2_12_28 ( .A(n668), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), .CO(
        \CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA1P S2_39_12 ( .A(\ab[39][12] ), .B(\CARRYB[38][12] ), .CI(\SUMB[38][13] ), 
        .CO(\CARRYB[39][12] ), .S(\SUMB[39][12] ) );
  FA1AP S2_11_34 ( .A(\CARRYB[10][34] ), .B(n632), .CI(\SUMB[10][35] ), .CO(
        \CARRYB[11][34] ), .S(\SUMB[11][34] ) );
  FA1AP S2_26_28 ( .A(\ab[28][26] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), 
        .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FA1P S2_26_20 ( .A(\CARRYB[25][20] ), .B(\ab[26][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA1P S2_18_13 ( .A(\CARRYB[17][13] ), .B(n695), .CI(\SUMB[17][14] ), .CO(
        \CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA1 S2_16_13 ( .A(\CARRYB[15][13] ), .B(n686), .CI(\SUMB[15][14] ), .CO(
        \CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA1 S2_8_12 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .CI(n532), .CO(
        \CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1P S3_13_46 ( .A(\ab[46][13] ), .B(\CARRYB[12][46] ), .CI(\ab[47][12] ), 
        .CO(\CARRYB[13][46] ), .S(\SUMB[13][46] ) );
  FA1P S3_4_46 ( .A(n302), .B(\CARRYB[3][46] ), .CI(n368), .CO(\CARRYB[4][46] ), .S(\SUMB[4][46] ) );
  FA1 S2_41_38 ( .A(\ab[41][38] ), .B(\CARRYB[40][38] ), .CI(\SUMB[40][39] ), 
        .CO(\CARRYB[41][38] ), .S(\SUMB[41][38] ) );
  FA1P S2_19_30 ( .A(\ab[30][19] ), .B(\CARRYB[18][30] ), .CI(\SUMB[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA1AP S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA1P S2_42_31 ( .A(\ab[42][31] ), .B(\CARRYB[41][31] ), .CI(\SUMB[41][32] ), 
        .CO(\CARRYB[42][31] ), .S(\SUMB[42][31] ) );
  FA1P S2_5_23 ( .A(n408), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), .CO(
        \CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S2_37_26 ( .A(\CARRYB[36][26] ), .B(\ab[37][26] ), .CI(\SUMB[36][27] ), 
        .CO(\CARRYB[37][26] ), .S(\SUMB[37][26] ) );
  FA1 S2_4_11 ( .A(n388), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), .CO(
        \CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1P S2_7_11 ( .A(n504), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), .CO(
        \CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1P S2_40_7 ( .A(n492), .B(\CARRYB[39][7] ), .CI(\SUMB[39][8] ), .CO(
        \CARRYB[40][7] ), .S(\SUMB[40][7] ) );
  FA1P S2_12_30 ( .A(n662), .B(\CARRYB[11][30] ), .CI(\SUMB[11][31] ), .CO(
        \CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA1P S2_19_23 ( .A(\CARRYB[18][23] ), .B(\ab[23][19] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA1AP S2_18_14 ( .A(n698), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), .CO(
        \CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA1P S2_37_7 ( .A(\CARRYB[36][7] ), .B(n472), .CI(\SUMB[36][8] ), .CO(
        \CARRYB[37][7] ), .S(\SUMB[37][7] ) );
  FA1AP S2_40_24 ( .A(\ab[40][24] ), .B(\CARRYB[39][24] ), .CI(\SUMB[39][25] ), 
        .CO(\CARRYB[40][24] ), .S(\SUMB[40][24] ) );
  FA1P S2_3_26 ( .A(n2288), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), .CO(
        \CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1AP S2_23_37 ( .A(\ab[37][23] ), .B(\CARRYB[22][37] ), .CI(\SUMB[22][38] ), 
        .CO(\CARRYB[23][37] ), .S(\SUMB[23][37] ) );
  FA1 S2_14_14 ( .A(\CARRYB[13][14] ), .B(n261), .CI(\SUMB[13][15] ), .CO(
        \CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_22_12 ( .A(\CARRYB[21][12] ), .B(n678), .CI(\SUMB[21][13] ), .CO(
        \CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA1A S2_36_18 ( .A(\CARRYB[35][18] ), .B(\ab[36][18] ), .CI(\SUMB[35][19] ), 
        .CO(\CARRYB[36][18] ), .S(\SUMB[36][18] ) );
  FA1 S2_46_12 ( .A(\CARRYB[45][12] ), .B(\ab[46][12] ), .CI(\SUMB[45][13] ), 
        .CO(\CARRYB[46][12] ), .S(\SUMB[46][12] ) );
  FA1AP S4_12 ( .A(\CARRYB[46][12] ), .B(\ab[47][12] ), .CI(\SUMB[46][13] ), 
        .CO(\CARRYB[47][12] ), .S(\SUMB[47][12] ) );
  FA1P S2_16_42 ( .A(\ab[42][16] ), .B(\CARRYB[15][42] ), .CI(\SUMB[15][43] ), 
        .CO(\CARRYB[16][42] ), .S(\SUMB[16][42] ) );
  FA1P S2_24_42 ( .A(\ab[42][24] ), .B(\CARRYB[23][42] ), .CI(\SUMB[23][43] ), 
        .CO(\CARRYB[24][42] ), .S(\SUMB[24][42] ) );
  FA1P S2_13_42 ( .A(\ab[42][13] ), .B(\CARRYB[12][42] ), .CI(\SUMB[12][43] ), 
        .CO(\CARRYB[13][42] ), .S(\SUMB[13][42] ) );
  FA1P S4_19 ( .A(\ab[47][19] ), .B(\CARRYB[46][19] ), .CI(\SUMB[46][20] ), 
        .CO(\CARRYB[47][19] ), .S(\SUMB[47][19] ) );
  FA1P S2_13_9 ( .A(n572), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), .CO(
        \CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1P S2_16_9 ( .A(n548), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), .CO(
        \CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1A S2_14_10 ( .A(n595), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), .CO(
        \CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1P S2_15_9 ( .A(n559), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), .CO(
        \CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1P S2_39_11 ( .A(\CARRYB[38][11] ), .B(\ab[39][11] ), .CI(\SUMB[38][12] ), 
        .CO(\CARRYB[39][11] ), .S(\SUMB[39][11] ) );
  FA1P S2_9_33 ( .A(n558), .B(\CARRYB[8][33] ), .CI(\SUMB[8][34] ), .CO(
        \CARRYB[9][33] ), .S(\SUMB[9][33] ) );
  FA1P S2_12_26 ( .A(\CARRYB[11][26] ), .B(n657), .CI(\SUMB[11][27] ), .CO(
        \CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA1AP S2_13_15 ( .A(n691), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), .CO(
        \CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_15_14 ( .A(n707), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), .CO(
        \CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA1P S2_11_14 ( .A(n625), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), .CO(
        \CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1AP S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA1AP S2_42_12 ( .A(\ab[42][12] ), .B(\CARRYB[41][12] ), .CI(\SUMB[41][13] ), 
        .CO(\CARRYB[42][12] ), .S(\SUMB[42][12] ) );
  FA1AP S2_29_27 ( .A(\SUMB[28][28] ), .B(\ab[29][27] ), .CI(\CARRYB[28][27] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA1AP S4_23 ( .A(\ab[47][23] ), .B(\CARRYB[46][23] ), .CI(\SUMB[46][24] ), 
        .CO(\CARRYB[47][23] ), .S(\SUMB[47][23] ) );
  FA1 S2_8_16 ( .A(\CARRYB[7][16] ), .B(n525), .CI(\SUMB[7][17] ), .CO(
        \CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1 S2_17_39 ( .A(\ab[39][17] ), .B(\CARRYB[16][39] ), .CI(\SUMB[16][40] ), 
        .CO(\CARRYB[17][39] ), .S(\SUMB[17][39] ) );
  FA1A S2_33_25 ( .A(\ab[33][25] ), .B(\CARRYB[32][25] ), .CI(\SUMB[32][26] ), 
        .CO(\CARRYB[33][25] ), .S(\SUMB[33][25] ) );
  FA1P S2_9_40 ( .A(n593), .B(\CARRYB[8][40] ), .CI(\SUMB[8][41] ), .CO(
        \CARRYB[9][40] ), .S(\SUMB[9][40] ) );
  FA1A S2_18_39 ( .A(\ab[39][18] ), .B(\CARRYB[17][39] ), .CI(\SUMB[17][40] ), 
        .CO(\CARRYB[18][39] ), .S(\SUMB[18][39] ) );
  FA1P S1_43_0 ( .A(n2200), .B(\CARRYB[42][0] ), .CI(\SUMB[42][1] ), .CO(
        \CARRYB[43][0] ), .S(\A1[41] ) );
  FA1P S2_39_9 ( .A(\CARRYB[38][9] ), .B(n570), .CI(\SUMB[38][10] ), .CO(
        \CARRYB[39][9] ), .S(\SUMB[39][9] ) );
  FA1P S2_3_12 ( .A(n351), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), .CO(
        \CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1 S2_37_25 ( .A(\ab[37][25] ), .B(\CARRYB[36][25] ), .CI(\SUMB[36][26] ), 
        .CO(\CARRYB[37][25] ), .S(\SUMB[37][25] ) );
  FA1P S2_45_8 ( .A(\CARRYB[44][8] ), .B(n521), .CI(\SUMB[44][9] ), .CO(
        \CARRYB[45][8] ), .S(\SUMB[45][8] ) );
  FA1 S2_46_8 ( .A(n503), .B(\CARRYB[45][8] ), .CI(\SUMB[45][9] ), .CO(
        \CARRYB[46][8] ), .S(\SUMB[46][8] ) );
  FA1P S2_34_5 ( .A(n403), .B(\CARRYB[33][5] ), .CI(\SUMB[33][6] ), .CO(
        \CARRYB[34][5] ), .S(\SUMB[34][5] ) );
  FA1P S2_2_10 ( .A(n345), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), .CO(
        \CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1 S2_3_10 ( .A(n355), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), .CO(
        \CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1P S2_22_6 ( .A(n441), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), .CO(
        \CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA1AP S2_16_40 ( .A(\ab[40][16] ), .B(\CARRYB[15][40] ), .CI(\SUMB[15][41] ), 
        .CO(\CARRYB[16][40] ), .S(\SUMB[16][40] ) );
  FA1P S2_40_32 ( .A(\ab[40][32] ), .B(\CARRYB[39][32] ), .CI(\SUMB[39][33] ), 
        .CO(\CARRYB[40][32] ), .S(\SUMB[40][32] ) );
  FA1P S2_26_40 ( .A(\ab[40][26] ), .B(\CARRYB[25][40] ), .CI(\SUMB[25][41] ), 
        .CO(\CARRYB[26][40] ), .S(\SUMB[26][40] ) );
  FA1A S2_18_33 ( .A(\CARRYB[17][33] ), .B(\ab[33][18] ), .CI(\SUMB[17][34] ), 
        .CO(\CARRYB[18][33] ), .S(\SUMB[18][33] ) );
  FA1P S2_11_39 ( .A(\ab[39][11] ), .B(\CARRYB[10][39] ), .CI(\SUMB[10][40] ), 
        .CO(\CARRYB[11][39] ), .S(\SUMB[11][39] ) );
  FA1 S2_26_36 ( .A(\CARRYB[25][36] ), .B(\ab[36][26] ), .CI(\SUMB[25][37] ), 
        .CO(\CARRYB[26][36] ), .S(\SUMB[26][36] ) );
  FA1AP S2_22_24 ( .A(\ab[24][22] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA1P S2_26_4 ( .A(n362), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), .CO(
        \CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA1P S2_27_4 ( .A(n2309), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), .CO(
        \CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA1A S1_30_0 ( .A(n2169), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), .CO(
        \CARRYB[30][0] ), .S(\A1[28] ) );
  FA1 S2_29_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA1P S2_41_31 ( .A(\ab[41][31] ), .B(\CARRYB[40][31] ), .CI(\SUMB[40][32] ), 
        .CO(\CARRYB[41][31] ), .S(\SUMB[41][31] ) );
  FA1P S2_44_19 ( .A(\CARRYB[43][19] ), .B(\ab[44][19] ), .CI(\SUMB[43][20] ), 
        .CO(\CARRYB[44][19] ), .S(\SUMB[44][19] ) );
  FA1 S2_29_20 ( .A(\CARRYB[28][20] ), .B(\ab[29][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA1AP S2_21_33 ( .A(\CARRYB[20][33] ), .B(\ab[33][21] ), .CI(\SUMB[20][34] ), 
        .CO(\CARRYB[21][33] ), .S(\SUMB[21][33] ) );
  FA1P S2_43_17 ( .A(\ab[43][17] ), .B(\CARRYB[42][17] ), .CI(\SUMB[42][18] ), 
        .CO(\CARRYB[43][17] ), .S(\SUMB[43][17] ) );
  FA1P S2_25_21 ( .A(\CARRYB[24][21] ), .B(\ab[25][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA1P S2_44_9 ( .A(\CARRYB[43][9] ), .B(\ab[9][44] ), .CI(\SUMB[43][10] ), 
        .CO(\CARRYB[44][9] ), .S(\SUMB[44][9] ) );
  FA1AP S2_34_11 ( .A(n632), .B(\CARRYB[33][11] ), .CI(\SUMB[33][12] ), .CO(
        \CARRYB[34][11] ), .S(\SUMB[34][11] ) );
  FA1P S2_38_23 ( .A(\ab[38][23] ), .B(\CARRYB[37][23] ), .CI(\SUMB[37][24] ), 
        .CO(\CARRYB[38][23] ), .S(\SUMB[38][23] ) );
  FA1P S2_21_22 ( .A(\ab[22][21] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA1AP S2_9_37 ( .A(n569), .B(\CARRYB[8][37] ), .CI(\SUMB[8][38] ), .CO(
        \CARRYB[9][37] ), .S(\SUMB[9][37] ) );
  FA1A S2_9_17 ( .A(n574), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), .CO(
        \CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1A S2_33_10 ( .A(n614), .B(\CARRYB[32][10] ), .CI(\SUMB[32][11] ), .CO(
        \CARRYB[33][10] ), .S(\SUMB[33][10] ) );
  FA1A S2_17_14 ( .A(n710), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), .CO(
        \CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA1 S2_12_35 ( .A(\SUMB[11][36] ), .B(\CARRYB[11][35] ), .CI(n672), .CO(
        \CARRYB[12][35] ), .S(\SUMB[12][35] ) );
  FA1P S3_6_46 ( .A(n457), .B(\CARRYB[5][46] ), .CI(n303), .CO(\CARRYB[6][46] ), .S(\SUMB[6][46] ) );
  FA1AP S4_29 ( .A(\ab[47][29] ), .B(\CARRYB[46][29] ), .CI(\SUMB[46][30] ), 
        .CO(\CARRYB[47][29] ), .S(\SUMB[47][29] ) );
  FA1AP S2_38_5 ( .A(\CARRYB[37][5] ), .B(n413), .CI(\SUMB[37][6] ), .CO(
        \CARRYB[38][5] ), .S(\SUMB[38][5] ) );
  FA1A S1_29_0 ( .A(n2171), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), .CO(
        \CARRYB[29][0] ), .S(\A1[27] ) );
  FA1 S2_38_4 ( .A(n370), .B(\CARRYB[37][4] ), .CI(\SUMB[37][5] ), .CO(
        \CARRYB[38][4] ), .S(\SUMB[38][4] ) );
  FA1P S2_35_34 ( .A(\ab[35][34] ), .B(\CARRYB[34][34] ), .CI(\SUMB[34][35] ), 
        .CO(\CARRYB[35][34] ), .S(\SUMB[35][34] ) );
  FA1P S4_7 ( .A(\ab[7][47] ), .B(\CARRYB[46][7] ), .CI(\SUMB[46][8] ), .CO(
        \CARRYB[47][7] ), .S(\SUMB[47][7] ) );
  FA1 S2_32_11 ( .A(\SUMB[31][12] ), .B(\CARRYB[31][11] ), .CI(n622), .CO(
        \CARRYB[32][11] ), .S(\SUMB[32][11] ) );
  FA1AP S4_17 ( .A(\ab[47][17] ), .B(\CARRYB[46][17] ), .CI(\SUMB[46][18] ), 
        .CO(\CARRYB[47][17] ), .S(\SUMB[47][17] ) );
  FA1AP S2_38_19 ( .A(\ab[38][19] ), .B(\CARRYB[37][19] ), .CI(\SUMB[37][20] ), 
        .CO(\CARRYB[38][19] ), .S(\SUMB[38][19] ) );
  FA1P S2_39_32 ( .A(\ab[39][32] ), .B(\CARRYB[38][32] ), .CI(\SUMB[38][33] ), 
        .CO(\CARRYB[39][32] ), .S(\SUMB[39][32] ) );
  FA1A S2_28_28 ( .A(\CARRYB[27][28] ), .B(n2375), .CI(\SUMB[27][29] ), .CO(
        \CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA1P S2_6_30 ( .A(\CARRYB[5][30] ), .B(n431), .CI(\SUMB[5][31] ), .CO(
        \CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA1AP S2_3_32 ( .A(n2283), .B(\CARRYB[2][32] ), .CI(\SUMB[2][33] ), .CO(
        \CARRYB[3][32] ), .S(\SUMB[3][32] ) );
  FA1AP S4_20 ( .A(\ab[47][20] ), .B(\CARRYB[46][20] ), .CI(\SUMB[46][21] ), 
        .CO(\CARRYB[47][20] ), .S(\SUMB[47][20] ) );
  FA1A S2_26_14 ( .A(n708), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), .CO(
        \CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA1 S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA1AP S2_9_27 ( .A(\CARRYB[8][27] ), .B(n573), .CI(\SUMB[8][28] ), .CO(
        \CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S2_27_14 ( .A(\CARRYB[26][14] ), .B(n712), .CI(\SUMB[26][15] ), .CO(
        \CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA1AP S2_35_27 ( .A(\ab[35][27] ), .B(\CARRYB[34][27] ), .CI(\SUMB[34][28] ), 
        .CO(\CARRYB[35][27] ), .S(\SUMB[35][27] ) );
  FA1P S2_40_22 ( .A(\ab[40][22] ), .B(\CARRYB[39][22] ), .CI(\SUMB[39][23] ), 
        .CO(\CARRYB[40][22] ), .S(\SUMB[40][22] ) );
  FA1P S2_41_20 ( .A(\ab[41][20] ), .B(\CARRYB[40][20] ), .CI(\SUMB[40][21] ), 
        .CO(\CARRYB[41][20] ), .S(\SUMB[41][20] ) );
  FA1A S2_34_7 ( .A(\CARRYB[33][7] ), .B(n481), .CI(\SUMB[33][8] ), .CO(
        \CARRYB[34][7] ), .S(\SUMB[34][7] ) );
  FA1P S2_4_1 ( .A(n2253), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1 S2_5_1 ( .A(n2219), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1 S4_0 ( .A(n1276), .B(\CARRYB[46][0] ), .CI(\SUMB[46][1] ), .CO(
        \CARRYB[47][0] ), .S(\SUMB[47][0] ) );
  FA1AP S2_41_26 ( .A(\ab[41][26] ), .B(\CARRYB[40][26] ), .CI(\SUMB[40][27] ), 
        .CO(\CARRYB[41][26] ), .S(\SUMB[41][26] ) );
  FA1A S2_44_7 ( .A(\CARRYB[43][7] ), .B(n486), .CI(\SUMB[43][8] ), .CO(
        \CARRYB[44][7] ), .S(\SUMB[44][7] ) );
  FA1A S2_7_12 ( .A(\CARRYB[6][12] ), .B(n508), .CI(\SUMB[6][13] ), .CO(
        \CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_35_15 ( .A(\ab[35][15] ), .B(\CARRYB[34][15] ), .CI(\SUMB[34][16] ), 
        .CO(\CARRYB[35][15] ), .S(\SUMB[35][15] ) );
  FA1A S2_29_1 ( .A(n2164), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), .CO(
        \CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA1AP S2_9_32 ( .A(\CARRYB[8][32] ), .B(n568), .CI(\SUMB[8][33] ), .CO(
        \CARRYB[9][32] ), .S(\SUMB[9][32] ) );
  FA1AP S2_40_20 ( .A(\CARRYB[39][20] ), .B(\ab[40][20] ), .CI(\SUMB[39][21] ), 
        .CO(\CARRYB[40][20] ), .S(\SUMB[40][20] ) );
  FA1AP S4_10 ( .A(\CARRYB[46][10] ), .B(\ab[47][10] ), .CI(\SUMB[46][11] ), 
        .CO(\CARRYB[47][10] ), .S(\SUMB[47][10] ) );
  FA1P S2_2_40 ( .A(\SUMB[1][41] ), .B(\CARRYB[1][40] ), .CI(n2250), .CO(
        \CARRYB[2][40] ), .S(\SUMB[2][40] ) );
  FA1P S2_3_40 ( .A(n2295), .B(\CARRYB[2][40] ), .CI(\SUMB[2][41] ), .CO(
        \CARRYB[3][40] ), .S(\SUMB[3][40] ) );
  FA1 S2_37_28 ( .A(\CARRYB[36][28] ), .B(\ab[37][28] ), .CI(\SUMB[36][29] ), 
        .CO(\CARRYB[37][28] ), .S(\SUMB[37][28] ) );
  FA1A S1_25_0 ( .A(n2235), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), .CO(
        \CARRYB[25][0] ), .S(\A1[23] ) );
  FA1P S2_4_8 ( .A(n391), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1P S2_32_5 ( .A(n407), .B(\CARRYB[31][5] ), .CI(\SUMB[31][6] ), .CO(
        \CARRYB[32][5] ), .S(\SUMB[32][5] ) );
  FA1P S2_33_5 ( .A(n401), .B(\CARRYB[32][5] ), .CI(\SUMB[32][6] ), .CO(
        \CARRYB[33][5] ), .S(\SUMB[33][5] ) );
  FA1 S2_9_7 ( .A(n509), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1P S2_12_8 ( .A(n532), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), .CO(
        \CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1P S2_13_7 ( .A(n480), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), .CO(
        \CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_18_6 ( .A(n464), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), .CO(
        \CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA1AP S2_41_10 ( .A(\CARRYB[40][10] ), .B(\ab[41][10] ), .CI(\SUMB[40][11] ), 
        .CO(\CARRYB[41][10] ), .S(\SUMB[41][10] ) );
  FA1 S2_40_19 ( .A(\CARRYB[39][19] ), .B(\ab[40][19] ), .CI(\SUMB[39][20] ), 
        .CO(\CARRYB[40][19] ), .S(\SUMB[40][19] ) );
  FA1A S2_35_25 ( .A(\CARRYB[34][25] ), .B(\ab[35][25] ), .CI(\SUMB[34][26] ), 
        .CO(\CARRYB[35][25] ), .S(\SUMB[35][25] ) );
  FA1AP S2_33_26 ( .A(\ab[33][26] ), .B(\CARRYB[32][26] ), .CI(\SUMB[32][27] ), 
        .CO(\CARRYB[33][26] ), .S(\SUMB[33][26] ) );
  FA1 S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA1A S2_15_13 ( .A(\CARRYB[14][13] ), .B(n691), .CI(\SUMB[14][14] ), .CO(
        \CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA1P S2_39_20 ( .A(\CARRYB[38][20] ), .B(\ab[39][20] ), .CI(\SUMB[38][21] ), 
        .CO(\CARRYB[39][20] ), .S(\SUMB[39][20] ) );
  FA1P S2_43_10 ( .A(\CARRYB[42][10] ), .B(\ab[43][10] ), .CI(\SUMB[42][11] ), 
        .CO(\CARRYB[43][10] ), .S(\SUMB[43][10] ) );
  FA1P S2_2_16 ( .A(n319), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), .CO(
        \CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1P S2_3_16 ( .A(\CARRYB[2][16] ), .B(n337), .CI(\SUMB[2][17] ), .CO(
        \CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1AP S2_42_8 ( .A(n550), .B(\CARRYB[41][8] ), .CI(\SUMB[41][9] ), .CO(
        \CARRYB[42][8] ), .S(\SUMB[42][8] ) );
  FA1AP S2_11_35 ( .A(n609), .B(\CARRYB[10][35] ), .CI(\SUMB[10][36] ), .CO(
        \CARRYB[11][35] ), .S(\SUMB[11][35] ) );
  FA1AP S2_13_16 ( .A(n686), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), .CO(
        \CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA1P S2_7_24 ( .A(n500), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), .CO(
        \CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA1AP S2_43_24 ( .A(\CARRYB[42][24] ), .B(\ab[43][24] ), .CI(\SUMB[42][25] ), 
        .CO(\CARRYB[43][24] ), .S(\SUMB[43][24] ) );
  FA1A S2_2_32 ( .A(n2211), .B(\CARRYB[1][32] ), .CI(\SUMB[1][33] ), .CO(
        \CARRYB[2][32] ), .S(\SUMB[2][32] ) );
  FA1A S2_46_3 ( .A(\CARRYB[45][3] ), .B(n2282), .CI(\SUMB[45][4] ), .CO(
        \CARRYB[46][3] ), .S(\SUMB[46][3] ) );
  FA1AP S2_36_20 ( .A(\ab[36][20] ), .B(\CARRYB[35][20] ), .CI(\SUMB[35][21] ), 
        .CO(\CARRYB[36][20] ), .S(\SUMB[36][20] ) );
  FA1P S2_6_7 ( .A(n482), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1P S2_3_8 ( .A(n350), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1P S2_23_2 ( .A(n2199), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), .CO(
        \CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA1 S2_2_26 ( .A(n2258), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), .CO(
        \CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1P S2_8_36 ( .A(n543), .B(\CARRYB[7][36] ), .CI(\SUMB[7][37] ), .CO(
        \CARRYB[8][36] ), .S(\SUMB[8][36] ) );
  FA1AP S2_30_29 ( .A(\ab[30][29] ), .B(\CARRYB[29][29] ), .CI(\SUMB[29][30] ), 
        .CO(\CARRYB[30][29] ), .S(\SUMB[30][29] ) );
  FA1AP S2_19_33 ( .A(\CARRYB[18][33] ), .B(\ab[33][19] ), .CI(\SUMB[18][34] ), 
        .CO(\CARRYB[19][33] ), .S(\SUMB[19][33] ) );
  FA1AP S2_12_32 ( .A(\CARRYB[11][32] ), .B(n669), .CI(\SUMB[11][33] ), .CO(
        \CARRYB[12][32] ), .S(\SUMB[12][32] ) );
  FA1P S2_42_5 ( .A(\CARRYB[41][5] ), .B(n454), .CI(\SUMB[41][6] ), .CO(
        \CARRYB[42][5] ), .S(\SUMB[42][5] ) );
  FA1AP S2_15_33 ( .A(\ab[33][15] ), .B(\CARRYB[14][33] ), .CI(\SUMB[14][34] ), 
        .CO(\CARRYB[15][33] ), .S(\SUMB[15][33] ) );
  FA1P S2_38_14 ( .A(\ab[38][14] ), .B(\CARRYB[37][14] ), .CI(\SUMB[37][15] ), 
        .CO(\CARRYB[38][14] ), .S(\SUMB[38][14] ) );
  FA1P S2_39_14 ( .A(\ab[39][14] ), .B(\CARRYB[38][14] ), .CI(\SUMB[38][15] ), 
        .CO(\CARRYB[39][14] ), .S(\SUMB[39][14] ) );
  FA1 S2_24_1 ( .A(n2240), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), .CO(
        \CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA1P S2_33_30 ( .A(\ab[33][30] ), .B(\CARRYB[32][30] ), .CI(\SUMB[32][31] ), 
        .CO(\CARRYB[33][30] ), .S(\SUMB[33][30] ) );
  FA1P S2_2_33 ( .A(n2212), .B(\CARRYB[1][33] ), .CI(\SUMB[1][34] ), .CO(
        \CARRYB[2][33] ), .S(\SUMB[2][33] ) );
  FA1AP S2_43_25 ( .A(\ab[43][25] ), .B(\CARRYB[42][25] ), .CI(\SUMB[42][26] ), 
        .CO(\CARRYB[43][25] ), .S(\SUMB[43][25] ) );
  FA1P S2_9_22 ( .A(n565), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), .CO(
        \CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA1AP S2_10_22 ( .A(n617), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), .CO(
        \CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA1P S2_28_14 ( .A(n706), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), .CO(
        \CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA1 S2_17_17 ( .A(\CARRYB[16][17] ), .B(n2355), .CI(\SUMB[16][18] ), .CO(
        \CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA1A S2_44_4 ( .A(\CARRYB[43][4] ), .B(n382), .CI(\SUMB[43][5] ), .CO(
        \CARRYB[44][4] ), .S(\SUMB[44][4] ) );
  FA1AP S2_34_12 ( .A(\CARRYB[33][12] ), .B(n674), .CI(\SUMB[33][13] ), .CO(
        \CARRYB[34][12] ), .S(\SUMB[34][12] ) );
  FA1P S2_20_22 ( .A(\SUMB[19][23] ), .B(\CARRYB[19][22] ), .CI(\ab[22][20] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA1A S2_43_28 ( .A(\ab[43][28] ), .B(\CARRYB[42][28] ), .CI(\SUMB[42][29] ), 
        .CO(\CARRYB[43][28] ), .S(\SUMB[43][28] ) );
  FA1 S2_17_38 ( .A(\ab[38][17] ), .B(\CARRYB[16][38] ), .CI(\SUMB[16][39] ), 
        .CO(\CARRYB[17][38] ), .S(\SUMB[17][38] ) );
  FA1P S1_40_0 ( .A(n2205), .B(\CARRYB[39][0] ), .CI(\SUMB[39][1] ), .CO(
        \CARRYB[40][0] ), .S(\A1[38] ) );
  FA1AP S2_36_12 ( .A(\CARRYB[35][12] ), .B(\ab[36][12] ), .CI(\SUMB[35][13] ), 
        .CO(\CARRYB[36][12] ), .S(\SUMB[36][12] ) );
  FA1A S2_2_29 ( .A(\CARRYB[1][29] ), .B(n2238), .CI(\SUMB[1][30] ), .CO(
        \CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1AP S2_6_36 ( .A(\CARRYB[5][36] ), .B(n443), .CI(\SUMB[5][37] ), .CO(
        \CARRYB[6][36] ), .S(\SUMB[6][36] ) );
  FA1P S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA1AP S2_29_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA1P S2_5_4 ( .A(n390), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1P S2_7_4 ( .A(n369), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1P S2_22_37 ( .A(\CARRYB[21][37] ), .B(\ab[37][22] ), .CI(\SUMB[21][38] ), 
        .CO(\CARRYB[22][37] ), .S(\SUMB[22][37] ) );
  FA1P S2_46_25 ( .A(\CARRYB[45][25] ), .B(\ab[46][25] ), .CI(\SUMB[45][26] ), 
        .CO(\CARRYB[46][25] ), .S(\SUMB[46][25] ) );
  FA1AP S2_38_26 ( .A(\CARRYB[37][26] ), .B(\ab[38][26] ), .CI(\SUMB[37][27] ), 
        .CO(\CARRYB[38][26] ), .S(\SUMB[38][26] ) );
  FA1 S2_20_1 ( .A(n270), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), .CO(
        \CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1P S1_39_0 ( .A(n334), .B(\CARRYB[38][0] ), .CI(\SUMB[38][1] ), .CO(
        \CARRYB[39][0] ), .S(\A1[37] ) );
  FA1AP S2_25_31 ( .A(\ab[31][25] ), .B(\CARRYB[24][31] ), .CI(\SUMB[24][32] ), 
        .CO(\CARRYB[25][31] ), .S(\SUMB[25][31] ) );
  FA1A S2_22_23 ( .A(\CARRYB[21][23] ), .B(\ab[23][22] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA1AP S2_7_14 ( .A(n513), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1 S2_16_12 ( .A(\CARRYB[15][12] ), .B(n312), .CI(\SUMB[15][13] ), .CO(
        \CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA1P S2_22_27 ( .A(\CARRYB[21][27] ), .B(\ab[27][22] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA1P S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA1P S2_36_23 ( .A(\ab[36][23] ), .B(\CARRYB[35][23] ), .CI(\SUMB[35][24] ), 
        .CO(\CARRYB[36][23] ), .S(\SUMB[36][23] ) );
  FA1P S2_37_23 ( .A(\ab[37][23] ), .B(\CARRYB[36][23] ), .CI(\SUMB[36][24] ), 
        .CO(\CARRYB[37][23] ), .S(\SUMB[37][23] ) );
  FA1A S2_23_30 ( .A(\CARRYB[22][30] ), .B(\ab[30][23] ), .CI(\SUMB[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FA1A S2_18_23 ( .A(\ab[23][18] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA1A S2_21_21 ( .A(n2362), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), .CO(
        \CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA1A S2_30_8 ( .A(\CARRYB[29][8] ), .B(n541), .CI(\SUMB[29][9] ), .CO(
        \CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA1 S2_5_22 ( .A(\CARRYB[4][22] ), .B(n380), .CI(\SUMB[4][23] ), .CO(
        \CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1AP S2_29_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA1AP S2_19_27 ( .A(\ab[27][19] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA1AP S2_26_26 ( .A(\CARRYB[25][26] ), .B(n2370), .CI(\SUMB[25][27] ), .CO(
        \CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA1 S2_23_29 ( .A(\ab[29][23] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA1A S2_18_29 ( .A(\CARRYB[17][29] ), .B(\ab[29][18] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA1A S2_37_21 ( .A(\ab[37][21] ), .B(\CARRYB[36][21] ), .CI(\SUMB[36][22] ), 
        .CO(\CARRYB[37][21] ), .S(\SUMB[37][21] ) );
  FA1AP S2_30_20 ( .A(\CARRYB[29][20] ), .B(\ab[30][20] ), .CI(\SUMB[29][21] ), 
        .CO(\CARRYB[30][20] ), .S(\SUMB[30][20] ) );
  FA1P S2_11_23 ( .A(n642), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), .CO(
        \CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1P S2_40_12 ( .A(\ab[40][12] ), .B(\CARRYB[39][12] ), .CI(\SUMB[39][13] ), 
        .CO(\CARRYB[40][12] ), .S(\SUMB[40][12] ) );
  FA1 S2_35_21 ( .A(\SUMB[34][22] ), .B(\CARRYB[34][21] ), .CI(\ab[35][21] ), 
        .CO(\CARRYB[35][21] ), .S(\SUMB[35][21] ) );
  FA1P S2_42_17 ( .A(\ab[42][17] ), .B(\CARRYB[41][17] ), .CI(\SUMB[41][18] ), 
        .CO(\CARRYB[42][17] ), .S(\SUMB[42][17] ) );
  FA1AP S2_19_8 ( .A(n540), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), .CO(
        \CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1P S2_25_40 ( .A(\ab[40][25] ), .B(\CARRYB[24][40] ), .CI(\SUMB[24][41] ), 
        .CO(\CARRYB[25][40] ), .S(\SUMB[25][40] ) );
  FA1P S2_40_34 ( .A(\ab[40][34] ), .B(\CARRYB[39][34] ), .CI(\SUMB[39][35] ), 
        .CO(\CARRYB[40][34] ), .S(\SUMB[40][34] ) );
  FA1A S2_30_24 ( .A(\ab[30][24] ), .B(\CARRYB[29][24] ), .CI(\SUMB[29][25] ), 
        .CO(\CARRYB[30][24] ), .S(\SUMB[30][24] ) );
  FA1A S2_33_29 ( .A(\CARRYB[32][29] ), .B(\ab[33][29] ), .CI(\SUMB[32][30] ), 
        .CO(\CARRYB[33][29] ), .S(\SUMB[33][29] ) );
  FA1 S2_29_25 ( .A(\CARRYB[28][25] ), .B(\ab[29][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA1AP S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA1AP S2_39_6 ( .A(\CARRYB[38][6] ), .B(n463), .CI(\SUMB[38][7] ), .CO(
        \CARRYB[39][6] ), .S(\SUMB[39][6] ) );
  FA1A S2_8_21 ( .A(\CARRYB[7][21] ), .B(n526), .CI(\SUMB[7][22] ), .CO(
        \CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA1 S2_18_30 ( .A(\ab[30][18] ), .B(\CARRYB[17][30] ), .CI(\SUMB[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA1P S2_2_43 ( .A(n2252), .B(\CARRYB[1][43] ), .CI(\SUMB[1][44] ), .CO(
        \CARRYB[2][43] ), .S(\SUMB[2][43] ) );
  FA1 S2_41_8 ( .A(n546), .B(\CARRYB[40][8] ), .CI(\SUMB[40][9] ), .CO(
        \CARRYB[41][8] ), .S(\SUMB[41][8] ) );
  FA1P S3_5_46 ( .A(n305), .B(\CARRYB[4][46] ), .CI(n406), .CO(\CARRYB[5][46] ), .S(\SUMB[5][46] ) );
  FA1AP S2_8_15 ( .A(n527), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), .CO(
        \CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1AP S2_2_24 ( .A(\CARRYB[1][24] ), .B(n2259), .CI(\SUMB[1][25] ), .CO(
        \CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA1P S2_20_28 ( .A(\CARRYB[19][28] ), .B(\ab[28][20] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA1AP S2_15_34 ( .A(\ab[34][15] ), .B(\CARRYB[14][34] ), .CI(\SUMB[14][35] ), 
        .CO(\CARRYB[15][34] ), .S(\SUMB[15][34] ) );
  FA1AP S2_19_35 ( .A(\CARRYB[18][35] ), .B(\ab[35][19] ), .CI(\SUMB[18][36] ), 
        .CO(\CARRYB[19][35] ), .S(\SUMB[19][35] ) );
  FA1AP S2_18_26 ( .A(\ab[26][18] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA1AP S2_16_30 ( .A(\CARRYB[15][30] ), .B(\ab[30][16] ), .CI(\SUMB[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA1P S2_34_15 ( .A(\CARRYB[33][15] ), .B(\ab[34][15] ), .CI(\SUMB[33][16] ), 
        .CO(\CARRYB[34][15] ), .S(\SUMB[34][15] ) );
  FA1A S2_38_13 ( .A(\ab[38][13] ), .B(\CARRYB[37][13] ), .CI(\SUMB[37][14] ), 
        .CO(\CARRYB[38][13] ), .S(\SUMB[38][13] ) );
  FA1P S2_8_33 ( .A(n537), .B(\CARRYB[7][33] ), .CI(\SUMB[7][34] ), .CO(
        \CARRYB[8][33] ), .S(\SUMB[8][33] ) );
  FA1 S2_28_36 ( .A(\ab[36][28] ), .B(\CARRYB[27][36] ), .CI(\SUMB[27][37] ), 
        .CO(\CARRYB[28][36] ), .S(\SUMB[28][36] ) );
  FA1AP S2_4_29 ( .A(\CARRYB[3][29] ), .B(n2299), .CI(\SUMB[3][30] ), .CO(
        \CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1 S2_15_24 ( .A(n726), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), .CO(
        \CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA1A S2_4_10 ( .A(n373), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), .CO(
        \CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1 S2_16_21 ( .A(\ab[21][16] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA1 S2_18_34 ( .A(\ab[34][18] ), .B(\CARRYB[17][34] ), .CI(\SUMB[17][35] ), 
        .CO(\CARRYB[18][34] ), .S(\SUMB[18][34] ) );
  FA1AP S2_19_34 ( .A(\ab[34][19] ), .B(\CARRYB[18][34] ), .CI(\SUMB[18][35] ), 
        .CO(\CARRYB[19][34] ), .S(\SUMB[19][34] ) );
  FA1A S2_36_14 ( .A(\ab[36][14] ), .B(\CARRYB[35][14] ), .CI(\SUMB[35][15] ), 
        .CO(\CARRYB[36][14] ), .S(\SUMB[36][14] ) );
  FA1P S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA1P S2_17_23 ( .A(\ab[23][17] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA1A S2_16_24 ( .A(\ab[24][16] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA1A S2_23_33 ( .A(\ab[33][23] ), .B(\CARRYB[22][33] ), .CI(\SUMB[22][34] ), 
        .CO(\CARRYB[23][33] ), .S(\SUMB[23][33] ) );
  FA1P S2_28_7 ( .A(n471), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), .CO(
        \CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA1P S2_29_7 ( .A(n502), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), .CO(
        \CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA1P S2_39_3 ( .A(n2305), .B(\CARRYB[38][3] ), .CI(\SUMB[38][4] ), .CO(
        \CARRYB[39][3] ), .S(\SUMB[39][3] ) );
  FA1A S2_11_12 ( .A(n644), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), .CO(
        \CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1P S2_35_31 ( .A(\ab[35][31] ), .B(\CARRYB[34][31] ), .CI(\SUMB[34][32] ), 
        .CO(\CARRYB[35][31] ), .S(\SUMB[35][31] ) );
  FA1 S2_6_17 ( .A(n436), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), .CO(
        \CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1P S2_24_12 ( .A(\CARRYB[23][12] ), .B(n660), .CI(\SUMB[23][13] ), .CO(
        \CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA1A S2_25_14 ( .A(n711), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), .CO(
        \CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA1P S2_39_16 ( .A(\CARRYB[38][16] ), .B(\ab[39][16] ), .CI(\SUMB[38][17] ), 
        .CO(\CARRYB[39][16] ), .S(\SUMB[39][16] ) );
  FA1P S2_42_15 ( .A(\ab[42][15] ), .B(\CARRYB[41][15] ), .CI(\SUMB[41][16] ), 
        .CO(\CARRYB[42][15] ), .S(\SUMB[42][15] ) );
  FA1AP S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA1P S2_32_10 ( .A(\CARRYB[31][10] ), .B(n598), .CI(\SUMB[31][11] ), .CO(
        \CARRYB[32][10] ), .S(\SUMB[32][10] ) );
  FA1 S2_46_28 ( .A(\ab[46][28] ), .B(\CARRYB[45][28] ), .CI(\SUMB[45][29] ), 
        .CO(\CARRYB[46][28] ), .S(\SUMB[46][28] ) );
  FA1A S2_23_16 ( .A(\CARRYB[22][16] ), .B(\ab[23][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA1A S2_9_16 ( .A(\CARRYB[8][16] ), .B(n548), .CI(\SUMB[8][17] ), .CO(
        \CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1A S2_31_11 ( .A(\CARRYB[30][11] ), .B(n631), .CI(\SUMB[30][12] ), .CO(
        \CARRYB[31][11] ), .S(\SUMB[31][11] ) );
  FA1P S2_24_29 ( .A(\CARRYB[23][29] ), .B(\ab[29][24] ), .CI(\SUMB[23][30] ), 
        .CO(\CARRYB[24][29] ), .S(\SUMB[24][29] ) );
  FA1A S2_17_33 ( .A(\ab[33][17] ), .B(\CARRYB[16][33] ), .CI(\SUMB[16][34] ), 
        .CO(\CARRYB[17][33] ), .S(\SUMB[17][33] ) );
  FA1 S2_10_15 ( .A(n588), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), .CO(
        \CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1P S2_2_18 ( .A(\CARRYB[1][18] ), .B(n2216), .CI(\SUMB[1][19] ), .CO(
        \CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1 S2_14_33 ( .A(\CARRYB[13][33] ), .B(\ab[33][14] ), .CI(\SUMB[13][34] ), 
        .CO(\CARRYB[14][33] ), .S(\SUMB[14][33] ) );
  FA1 S2_31_28 ( .A(\CARRYB[30][28] ), .B(\ab[31][28] ), .CI(\SUMB[30][29] ), 
        .CO(\CARRYB[31][28] ), .S(\SUMB[31][28] ) );
  FA1P S2_45_9 ( .A(\CARRYB[44][9] ), .B(\ab[9][45] ), .CI(\SUMB[44][10] ), 
        .CO(\CARRYB[45][9] ), .S(\SUMB[45][9] ) );
  FA1P S2_30_22 ( .A(\ab[30][22] ), .B(\CARRYB[29][22] ), .CI(\SUMB[29][23] ), 
        .CO(\CARRYB[30][22] ), .S(\SUMB[30][22] ) );
  FA1P S2_31_22 ( .A(\CARRYB[30][22] ), .B(\ab[31][22] ), .CI(\SUMB[30][23] ), 
        .CO(\CARRYB[31][22] ), .S(\SUMB[31][22] ) );
  FA1P S2_29_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA1P S2_6_31 ( .A(n465), .B(\CARRYB[5][31] ), .CI(\SUMB[5][32] ), .CO(
        \CARRYB[6][31] ), .S(\SUMB[6][31] ) );
  FA1 S2_18_12 ( .A(\SUMB[17][13] ), .B(\CARRYB[17][12] ), .CI(n664), .CO(
        \CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA1 S2_27_8 ( .A(n524), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), .CO(
        \CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA1P S2_34_18 ( .A(\ab[34][18] ), .B(\CARRYB[33][18] ), .CI(\SUMB[33][19] ), 
        .CO(\CARRYB[34][18] ), .S(\SUMB[34][18] ) );
  FA1P S2_24_38 ( .A(\ab[38][24] ), .B(\CARRYB[23][38] ), .CI(\SUMB[23][39] ), 
        .CO(\CARRYB[24][38] ), .S(\SUMB[24][38] ) );
  FA1AP S2_42_30 ( .A(\ab[42][30] ), .B(\CARRYB[41][30] ), .CI(\SUMB[41][31] ), 
        .CO(\CARRYB[42][30] ), .S(\SUMB[42][30] ) );
  FA1AP S2_41_29 ( .A(\ab[41][29] ), .B(\CARRYB[40][29] ), .CI(\SUMB[40][30] ), 
        .CO(\CARRYB[41][29] ), .S(\SUMB[41][29] ) );
  FA1A S2_17_12 ( .A(\CARRYB[16][12] ), .B(n677), .CI(\SUMB[16][13] ), .CO(
        \CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA1AP S2_13_19 ( .A(\CARRYB[12][19] ), .B(n679), .CI(\SUMB[12][20] ), .CO(
        \CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA1P S2_16_23 ( .A(\CARRYB[15][23] ), .B(\ab[23][16] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA1P S2_17_1 ( .A(n2231), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), .CO(
        \CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1 S1_24_0 ( .A(n2236), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), .CO(
        \CARRYB[24][0] ), .S(\A1[22] ) );
  FA1AP S2_13_33 ( .A(\ab[33][13] ), .B(\CARRYB[12][33] ), .CI(\SUMB[12][34] ), 
        .CO(\CARRYB[13][33] ), .S(\SUMB[13][33] ) );
  FA1P S2_40_6 ( .A(n458), .B(\SUMB[39][7] ), .CI(\CARRYB[39][6] ), .CO(
        \CARRYB[40][6] ), .S(\SUMB[40][6] ) );
  FA1P S2_34_16 ( .A(\ab[34][16] ), .B(\CARRYB[33][16] ), .CI(\SUMB[33][17] ), 
        .CO(\CARRYB[34][16] ), .S(\SUMB[34][16] ) );
  FA1P S2_36_15 ( .A(\ab[36][15] ), .B(\CARRYB[35][15] ), .CI(\SUMB[35][16] ), 
        .CO(\CARRYB[36][15] ), .S(\SUMB[36][15] ) );
  FA1AP S2_32_12 ( .A(\CARRYB[31][12] ), .B(n669), .CI(\SUMB[31][13] ), .CO(
        \CARRYB[32][12] ), .S(\SUMB[32][12] ) );
  FA1A S2_24_15 ( .A(\CARRYB[23][15] ), .B(n726), .CI(\SUMB[23][16] ), .CO(
        \CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA1 S2_36_13 ( .A(\SUMB[35][14] ), .B(\CARRYB[35][13] ), .CI(\ab[36][13] ), 
        .CO(\CARRYB[36][13] ), .S(\SUMB[36][13] ) );
  FA1P S2_23_10 ( .A(\CARRYB[22][10] ), .B(n603), .CI(\SUMB[22][11] ), .CO(
        \CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA1 S2_42_29 ( .A(\CARRYB[41][29] ), .B(\ab[42][29] ), .CI(\SUMB[41][30] ), 
        .CO(\CARRYB[42][29] ), .S(\SUMB[42][29] ) );
  FA1P S2_35_32 ( .A(\ab[35][32] ), .B(\CARRYB[34][32] ), .CI(\SUMB[34][33] ), 
        .CO(\CARRYB[35][32] ), .S(\SUMB[35][32] ) );
  FA1AP S2_36_33 ( .A(\CARRYB[35][33] ), .B(\ab[36][33] ), .CI(\SUMB[35][34] ), 
        .CO(\CARRYB[36][33] ), .S(\SUMB[36][33] ) );
  FA1A S2_2_30 ( .A(\CARRYB[1][30] ), .B(n2208), .CI(\SUMB[1][31] ), .CO(
        \CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  FA1P S2_41_25 ( .A(\CARRYB[40][25] ), .B(\ab[41][25] ), .CI(\SUMB[40][26] ), 
        .CO(\CARRYB[41][25] ), .S(\SUMB[41][25] ) );
  FA1P S2_34_14 ( .A(\CARRYB[33][14] ), .B(\ab[34][14] ), .CI(\SUMB[33][15] ), 
        .CO(\CARRYB[34][14] ), .S(\SUMB[34][14] ) );
  FA1 S2_32_15 ( .A(\CARRYB[31][15] ), .B(\ab[32][15] ), .CI(\SUMB[31][16] ), 
        .CO(\CARRYB[32][15] ), .S(\SUMB[32][15] ) );
  FA1A S2_36_10 ( .A(\CARRYB[35][10] ), .B(n601), .CI(\SUMB[35][11] ), .CO(
        \CARRYB[36][10] ), .S(\SUMB[36][10] ) );
  FA1 S2_38_7 ( .A(\CARRYB[37][7] ), .B(n490), .CI(\SUMB[37][8] ), .CO(
        \CARRYB[38][7] ), .S(\SUMB[38][7] ) );
  FA1P S2_41_6 ( .A(n493), .B(\CARRYB[40][6] ), .CI(\SUMB[40][7] ), .CO(
        \CARRYB[41][6] ), .S(\SUMB[41][6] ) );
  FA1AP S2_37_8 ( .A(n551), .B(\CARRYB[36][8] ), .CI(\SUMB[36][9] ), .CO(
        \CARRYB[37][8] ), .S(\SUMB[37][8] ) );
  FA1P S2_10_18 ( .A(n602), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), .CO(
        \CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1A S2_33_15 ( .A(\CARRYB[32][15] ), .B(\ab[33][15] ), .CI(\SUMB[32][16] ), 
        .CO(\CARRYB[33][15] ), .S(\SUMB[33][15] ) );
  FA1P S2_12_13 ( .A(\CARRYB[11][13] ), .B(n654), .CI(\SUMB[11][14] ), .CO(
        \CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1 S2_10_31 ( .A(n585), .B(\CARRYB[9][31] ), .CI(\SUMB[9][32] ), .CO(
        \CARRYB[10][31] ), .S(\SUMB[10][31] ) );
  FA1A S2_22_10 ( .A(\CARRYB[21][10] ), .B(n617), .CI(\SUMB[21][11] ), .CO(
        \CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA1P S2_25_25 ( .A(n2369), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), .CO(
        \CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA1AP S2_13_30 ( .A(n692), .B(\CARRYB[12][30] ), .CI(\SUMB[12][31] ), .CO(
        \CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA1P S2_16_20 ( .A(\CARRYB[15][20] ), .B(\ab[20][16] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA1A S2_45_7 ( .A(n494), .B(\CARRYB[44][7] ), .CI(\SUMB[44][8] ), .CO(
        \CARRYB[45][7] ), .S(\SUMB[45][7] ) );
  FA1A S2_2_19 ( .A(\CARRYB[1][19] ), .B(n2215), .CI(\SUMB[1][20] ), .CO(
        \CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA1AP S2_25_33 ( .A(\CARRYB[24][33] ), .B(\ab[33][25] ), .CI(\SUMB[24][34] ), 
        .CO(\CARRYB[25][33] ), .S(\SUMB[25][33] ) );
  FA1 S2_36_9 ( .A(\SUMB[35][10] ), .B(\CARRYB[35][9] ), .CI(n567), .CO(
        \CARRYB[36][9] ), .S(\SUMB[36][9] ) );
  FA1AP S2_32_13 ( .A(\CARRYB[31][13] ), .B(n694), .CI(\SUMB[31][14] ), .CO(
        \CARRYB[32][13] ), .S(\SUMB[32][13] ) );
  FA1 S2_45_26 ( .A(\CARRYB[44][26] ), .B(\ab[45][26] ), .CI(\SUMB[44][27] ), 
        .CO(\CARRYB[45][26] ), .S(\SUMB[45][26] ) );
  FA1 S2_22_26 ( .A(\ab[26][22] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA1A S2_40_13 ( .A(\CARRYB[39][13] ), .B(\ab[40][13] ), .CI(\SUMB[39][14] ), 
        .CO(\CARRYB[40][13] ), .S(\SUMB[40][13] ) );
  FA1A S2_17_31 ( .A(\ab[31][17] ), .B(\CARRYB[16][31] ), .CI(\SUMB[16][32] ), 
        .CO(\CARRYB[17][31] ), .S(\SUMB[17][31] ) );
  FA1 S2_22_30 ( .A(\CARRYB[21][30] ), .B(\ab[30][22] ), .CI(\SUMB[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA1AP S2_17_28 ( .A(\ab[28][17] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA1 S2_17_27 ( .A(\ab[27][17] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA1AP S2_45_15 ( .A(\ab[45][15] ), .B(\CARRYB[44][15] ), .CI(\SUMB[44][16] ), 
        .CO(\CARRYB[45][15] ), .S(\SUMB[45][15] ) );
  FA1AP S2_45_14 ( .A(\CARRYB[44][14] ), .B(\ab[45][14] ), .CI(\SUMB[44][15] ), 
        .CO(\CARRYB[45][14] ), .S(\SUMB[45][14] ) );
  FA1 S2_9_30 ( .A(n592), .B(\CARRYB[8][30] ), .CI(\SUMB[8][31] ), .CO(
        \CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA1 S2_20_27 ( .A(\ab[27][20] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA1A S2_11_25 ( .A(n633), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), .CO(
        \CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1P S2_41_21 ( .A(\ab[41][21] ), .B(\CARRYB[40][21] ), .CI(\SUMB[40][22] ), 
        .CO(\CARRYB[41][21] ), .S(\SUMB[41][21] ) );
  FA1P S2_17_30 ( .A(\CARRYB[16][30] ), .B(\ab[30][17] ), .CI(\SUMB[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA1 S2_2_25 ( .A(\CARRYB[1][25] ), .B(n2207), .CI(\SUMB[1][26] ), .CO(
        \CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1P S2_4_9 ( .A(n387), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1P S2_11_8 ( .A(n542), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(
        \CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1P S2_33_4 ( .A(n2306), .B(\CARRYB[32][4] ), .CI(\SUMB[32][5] ), .CO(
        \CARRYB[33][4] ), .S(\SUMB[33][4] ) );
  FA1 S2_40_3 ( .A(n2295), .B(\CARRYB[39][3] ), .CI(\SUMB[39][4] ), .CO(
        \CARRYB[40][3] ), .S(\SUMB[40][3] ) );
  FA1A S2_7_9 ( .A(n509), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_15_1 ( .A(n2218), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1P S2_16_1 ( .A(n2187), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), .CO(
        \CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1P S2_18_1 ( .A(n2168), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), .CO(
        \CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA1A S2_20_24 ( .A(\ab[24][20] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA1P S2_2_20 ( .A(n2176), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), .CO(
        \CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1A S2_8_26 ( .A(n523), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), .CO(
        \CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1AP S2_6_27 ( .A(n442), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), .CO(
        \CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA1A S2_29_36 ( .A(\ab[36][29] ), .B(\CARRYB[28][36] ), .CI(\SUMB[28][37] ), 
        .CO(\CARRYB[29][36] ), .S(\SUMB[29][36] ) );
  FA1 S1_28_0 ( .A(n2174), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), .CO(
        \CARRYB[28][0] ), .S(\A1[26] ) );
  FA1AP S2_27_35 ( .A(\CARRYB[26][35] ), .B(\ab[35][27] ), .CI(\SUMB[26][36] ), 
        .CO(\CARRYB[27][35] ), .S(\SUMB[27][35] ) );
  FA1P S4_33 ( .A(\ab[47][33] ), .B(\CARRYB[46][33] ), .CI(\SUMB[46][34] ), 
        .CO(\CARRYB[47][33] ), .S(\SUMB[47][33] ) );
  FA1A S2_40_31 ( .A(\ab[40][31] ), .B(\CARRYB[39][31] ), .CI(\SUMB[39][32] ), 
        .CO(\CARRYB[40][31] ), .S(\SUMB[40][31] ) );
  FA1A S2_25_36 ( .A(\CARRYB[24][36] ), .B(\ab[36][25] ), .CI(\SUMB[24][37] ), 
        .CO(\CARRYB[25][36] ), .S(\SUMB[25][36] ) );
  FA1 S2_24_26 ( .A(\CARRYB[23][26] ), .B(\ab[26][24] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA1P S2_31_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FA1A S2_40_29 ( .A(\CARRYB[39][29] ), .B(\ab[40][29] ), .CI(\SUMB[39][30] ), 
        .CO(\CARRYB[40][29] ), .S(\SUMB[40][29] ) );
  FA1P S2_46_7 ( .A(\CARRYB[45][7] ), .B(n306), .CI(\SUMB[45][8] ), .CO(
        \CARRYB[46][7] ), .S(\SUMB[46][7] ) );
  FA1A S2_9_29 ( .A(n575), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), .CO(
        \CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1 S2_37_24 ( .A(\CARRYB[36][24] ), .B(\ab[37][24] ), .CI(\SUMB[36][25] ), 
        .CO(\CARRYB[37][24] ), .S(\SUMB[37][24] ) );
  FA1P S1_6_0 ( .A(n285), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1 S2_40_30 ( .A(\ab[40][30] ), .B(\CARRYB[39][30] ), .CI(\SUMB[39][31] ), 
        .CO(\CARRYB[40][30] ), .S(\SUMB[40][30] ) );
  FA1P S2_36_32 ( .A(\ab[36][32] ), .B(\CARRYB[35][32] ), .CI(\SUMB[35][33] ), 
        .CO(\CARRYB[36][32] ), .S(\SUMB[36][32] ) );
  FA1P S2_33_33 ( .A(n2392), .B(\CARRYB[32][33] ), .CI(\SUMB[32][34] ), .CO(
        \CARRYB[33][33] ), .S(\SUMB[33][33] ) );
  FA1P S2_38_31 ( .A(\ab[38][31] ), .B(\CARRYB[37][31] ), .CI(\SUMB[37][32] ), 
        .CO(\CARRYB[38][31] ), .S(\SUMB[38][31] ) );
  FA1 S2_43_21 ( .A(\ab[43][21] ), .B(\CARRYB[42][21] ), .CI(\SUMB[42][22] ), 
        .CO(\CARRYB[43][21] ), .S(\SUMB[43][21] ) );
  FA1P S2_5_35 ( .A(n374), .B(\CARRYB[4][35] ), .CI(\SUMB[4][36] ), .CO(
        \CARRYB[5][35] ), .S(\SUMB[5][35] ) );
  FA1P S2_15_30 ( .A(\ab[30][15] ), .B(\CARRYB[14][30] ), .CI(\SUMB[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA1A S2_42_3 ( .A(n2296), .B(\CARRYB[41][3] ), .CI(\SUMB[41][4] ), .CO(
        \CARRYB[42][3] ), .S(\SUMB[42][3] ) );
  FA1P S2_43_3 ( .A(n2297), .B(\CARRYB[42][3] ), .CI(\SUMB[42][4] ), .CO(
        \CARRYB[43][3] ), .S(\SUMB[43][3] ) );
  FA1 S2_7_27 ( .A(\CARRYB[6][27] ), .B(n498), .CI(\SUMB[6][28] ), .CO(
        \CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1A S2_23_27 ( .A(\CARRYB[22][27] ), .B(\ab[27][23] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA1A S2_38_11 ( .A(\ab[38][11] ), .B(\CARRYB[37][11] ), .CI(\SUMB[37][12] ), 
        .CO(\CARRYB[38][11] ), .S(\SUMB[38][11] ) );
  FA1 S2_38_38 ( .A(n2404), .B(\CARRYB[37][38] ), .CI(\SUMB[37][39] ), .CO(
        \CARRYB[38][38] ), .S(\SUMB[38][38] ) );
  FA1P S2_17_34 ( .A(\ab[34][17] ), .B(\CARRYB[16][34] ), .CI(\SUMB[16][35] ), 
        .CO(\CARRYB[17][34] ), .S(\SUMB[17][34] ) );
  FA1A S2_32_28 ( .A(\ab[32][28] ), .B(\CARRYB[31][28] ), .CI(\SUMB[31][29] ), 
        .CO(\CARRYB[32][28] ), .S(\SUMB[32][28] ) );
  FA1 S2_19_31 ( .A(\ab[31][19] ), .B(\CARRYB[18][31] ), .CI(\SUMB[18][32] ), 
        .CO(\CARRYB[19][31] ), .S(\SUMB[19][31] ) );
  FA1P S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA1 S2_33_27 ( .A(\SUMB[32][28] ), .B(\CARRYB[32][27] ), .CI(\ab[33][27] ), 
        .CO(\CARRYB[33][27] ), .S(\SUMB[33][27] ) );
  FA1A S2_21_20 ( .A(\CARRYB[20][20] ), .B(\ab[21][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA1AP S2_19_21 ( .A(\CARRYB[18][21] ), .B(\ab[21][19] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA1P S2_40_21 ( .A(\ab[40][21] ), .B(\CARRYB[39][21] ), .CI(\SUMB[39][22] ), 
        .CO(\CARRYB[40][21] ), .S(\SUMB[40][21] ) );
  FA1P S2_8_40 ( .A(n545), .B(\CARRYB[7][40] ), .CI(\SUMB[7][41] ), .CO(
        \CARRYB[8][40] ), .S(\SUMB[8][40] ) );
  FA1AP S2_31_24 ( .A(\CARRYB[30][24] ), .B(\ab[31][24] ), .CI(\SUMB[30][25] ), 
        .CO(\CARRYB[31][24] ), .S(\SUMB[31][24] ) );
  FA1 S2_37_22 ( .A(\SUMB[36][23] ), .B(\CARRYB[36][22] ), .CI(\ab[37][22] ), 
        .CO(\CARRYB[37][22] ), .S(\SUMB[37][22] ) );
  FA1P S2_3_20 ( .A(n2280), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), .CO(
        \CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1P S2_7_36 ( .A(n501), .B(\CARRYB[6][36] ), .CI(\SUMB[6][37] ), .CO(
        \CARRYB[7][36] ), .S(\SUMB[7][36] ) );
  FA1P S2_37_6 ( .A(\SUMB[36][7] ), .B(\CARRYB[36][6] ), .CI(n440), .CO(
        \CARRYB[37][6] ), .S(\SUMB[37][6] ) );
  FA1P S2_12_36 ( .A(\ab[36][12] ), .B(\CARRYB[11][36] ), .CI(\SUMB[11][37] ), 
        .CO(\CARRYB[12][36] ), .S(\SUMB[12][36] ) );
  FA1AP S2_11_36 ( .A(n643), .B(\CARRYB[10][36] ), .CI(\SUMB[10][37] ), .CO(
        \CARRYB[11][36] ), .S(\SUMB[11][36] ) );
  FA1P S2_14_35 ( .A(\ab[35][14] ), .B(\CARRYB[13][35] ), .CI(\SUMB[13][36] ), 
        .CO(\CARRYB[14][35] ), .S(\SUMB[14][35] ) );
  FA1P S2_15_17 ( .A(\CARRYB[14][17] ), .B(n717), .CI(\SUMB[14][18] ), .CO(
        \CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA1 S2_34_22 ( .A(\CARRYB[33][22] ), .B(\ab[34][22] ), .CI(\SUMB[33][23] ), 
        .CO(\CARRYB[34][22] ), .S(\SUMB[34][22] ) );
  FA1P S2_16_15 ( .A(n722), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), .CO(
        \CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA1 S2_10_39 ( .A(n640), .B(\CARRYB[9][39] ), .CI(\SUMB[9][40] ), .CO(
        \CARRYB[10][39] ), .S(\SUMB[10][39] ) );
  FA1A S2_10_14 ( .A(\CARRYB[9][14] ), .B(n595), .CI(\SUMB[9][15] ), .CO(
        \CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1AP S2_20_16 ( .A(\CARRYB[19][16] ), .B(\ab[20][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA1P S2_27_15 ( .A(\CARRYB[26][15] ), .B(n718), .CI(\SUMB[26][16] ), .CO(
        \CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA1A S2_42_11 ( .A(\ab[42][11] ), .B(\CARRYB[41][11] ), .CI(\SUMB[41][12] ), 
        .CO(\CARRYB[42][11] ), .S(\SUMB[42][11] ) );
  FA1A S2_23_15 ( .A(\CARRYB[22][15] ), .B(n716), .CI(\SUMB[22][16] ), .CO(
        \CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA1A S2_21_16 ( .A(\CARRYB[20][16] ), .B(\ab[21][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA1A S2_22_16 ( .A(\CARRYB[21][16] ), .B(\ab[22][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA1 S2_17_26 ( .A(\ab[26][17] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA1A S2_18_25 ( .A(\ab[25][18] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA1 S2_37_30 ( .A(\ab[37][30] ), .B(\CARRYB[36][30] ), .CI(\SUMB[36][31] ), 
        .CO(\CARRYB[37][30] ), .S(\SUMB[37][30] ) );
  FA1 S2_14_29 ( .A(n702), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), .CO(
        \CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA1AP S2_11_26 ( .A(\CARRYB[10][26] ), .B(n630), .CI(\SUMB[10][27] ), .CO(
        \CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1 S2_18_11 ( .A(\CARRYB[17][11] ), .B(n638), .CI(\SUMB[17][12] ), .CO(
        \CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA1AP S2_19_11 ( .A(\CARRYB[18][11] ), .B(n618), .CI(\SUMB[18][12] ), .CO(
        \CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA1AP S2_36_11 ( .A(\CARRYB[35][11] ), .B(n643), .CI(\SUMB[35][12] ), .CO(
        \CARRYB[36][11] ), .S(\SUMB[36][11] ) );
  FA1P S2_39_21 ( .A(\ab[39][21] ), .B(\CARRYB[38][21] ), .CI(\SUMB[38][22] ), 
        .CO(\CARRYB[39][21] ), .S(\SUMB[39][21] ) );
  FA1P S2_7_13 ( .A(n480), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), .CO(
        \CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1P S2_6_13 ( .A(n461), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), .CO(
        \CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1AP S2_11_17 ( .A(n629), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), .CO(
        \CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1A S2_11_28 ( .A(\CARRYB[10][28] ), .B(n628), .CI(\SUMB[10][29] ), .CO(
        \CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1 S2_20_21 ( .A(\CARRYB[19][21] ), .B(\ab[21][20] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA1AP S2_38_25 ( .A(\CARRYB[37][25] ), .B(\ab[38][25] ), .CI(\SUMB[37][26] ), 
        .CO(\CARRYB[38][25] ), .S(\SUMB[38][25] ) );
  FA1P S2_13_31 ( .A(n685), .B(\CARRYB[12][31] ), .CI(\SUMB[12][32] ), .CO(
        \CARRYB[13][31] ), .S(\SUMB[13][31] ) );
  FA1A S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA1 S2_7_34 ( .A(\CARRYB[6][34] ), .B(n481), .CI(\SUMB[6][35] ), .CO(
        \CARRYB[7][34] ), .S(\SUMB[7][34] ) );
  FA1 S2_21_30 ( .A(\ab[30][21] ), .B(\CARRYB[20][30] ), .CI(\SUMB[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA1P S2_23_26 ( .A(\CARRYB[22][26] ), .B(\ab[26][23] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA1P S2_31_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FA1P S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA1P S2_15_39 ( .A(\CARRYB[14][39] ), .B(\ab[39][15] ), .CI(\SUMB[14][40] ), 
        .CO(\CARRYB[15][39] ), .S(\SUMB[15][39] ) );
  FA1P S2_33_31 ( .A(\CARRYB[32][31] ), .B(\ab[33][31] ), .CI(\SUMB[32][32] ), 
        .CO(\CARRYB[33][31] ), .S(\SUMB[33][31] ) );
  FA1P S2_46_33 ( .A(\ab[46][33] ), .B(\CARRYB[45][33] ), .CI(\SUMB[45][34] ), 
        .CO(\CARRYB[46][33] ), .S(\SUMB[46][33] ) );
  FA1 S2_30_28 ( .A(\CARRYB[29][28] ), .B(\ab[30][28] ), .CI(\SUMB[29][29] ), 
        .CO(\CARRYB[30][28] ), .S(\SUMB[30][28] ) );
  FA1A S2_25_10 ( .A(n591), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), .CO(
        \CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA1A S2_38_21 ( .A(\CARRYB[37][21] ), .B(\ab[38][21] ), .CI(\SUMB[37][22] ), 
        .CO(\CARRYB[38][21] ), .S(\SUMB[38][21] ) );
  FA1P S2_30_12 ( .A(\SUMB[29][13] ), .B(\CARRYB[29][12] ), .CI(n662), .CO(
        \CARRYB[30][12] ), .S(\SUMB[30][12] ) );
  FA1 S2_24_13 ( .A(n690), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), .CO(
        \CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA1AP S2_30_14 ( .A(\CARRYB[29][14] ), .B(n705), .CI(\SUMB[29][15] ), .CO(
        \CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FA1P S2_18_19 ( .A(\CARRYB[17][19] ), .B(\ab[19][18] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA1A S1_7_0 ( .A(n2255), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_12_0 ( .A(n2183), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), .CO(
        \CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S2_26_1 ( .A(n2220), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), .CO(
        \CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA1A S2_7_1 ( .A(n2244), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_3_1 ( .A(n2429), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_12_1 ( .A(n2192), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), .CO(
        \CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S2_11_1 ( .A(n2180), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(
        \CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_27_2 ( .A(n2209), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), .CO(
        \CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA1A S2_4_3 ( .A(n344), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_8_3 ( .A(n350), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_7_2 ( .A(n338), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_2_3 ( .A(n301), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S4_39 ( .A(\ab[47][39] ), .B(\CARRYB[46][39] ), .CI(\SUMB[46][40] ), 
        .CO(\CARRYB[47][39] ), .S(\SUMB[47][39] ) );
  FA1A S4_15 ( .A(\ab[47][15] ), .B(\CARRYB[46][15] ), .CI(\SUMB[46][16] ), 
        .CO(\CARRYB[47][15] ), .S(\SUMB[47][15] ) );
  FA1A S3_46_46 ( .A(n256), .B(\CARRYB[45][46] ), .CI(\ab[47][45] ), .CO(
        \CARRYB[46][46] ), .S(\SUMB[46][46] ) );
  FA1A S4_45 ( .A(\ab[47][45] ), .B(\CARRYB[46][45] ), .CI(\SUMB[46][46] ), 
        .CO(\CARRYB[47][45] ), .S(\SUMB[47][45] ) );
  FA1A S4_44 ( .A(\ab[47][44] ), .B(\CARRYB[46][44] ), .CI(\SUMB[46][45] ), 
        .CO(\CARRYB[47][44] ), .S(\SUMB[47][44] ) );
  FA1A S4_13 ( .A(\ab[47][13] ), .B(\CARRYB[46][13] ), .CI(\SUMB[46][14] ), 
        .CO(\CARRYB[47][13] ), .S(\SUMB[47][13] ) );
  FA1A S4_14 ( .A(\ab[47][14] ), .B(\CARRYB[46][14] ), .CI(\SUMB[46][15] ), 
        .CO(\CARRYB[47][14] ), .S(\SUMB[47][14] ) );
  FA1A S2_5_3 ( .A(n2310), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S3_45_46 ( .A(\ab[46][45] ), .B(\CARRYB[44][46] ), .CI(\ab[47][44] ), 
        .CO(\CARRYB[45][46] ), .S(\SUMB[45][46] ) );
  FA1A S2_23_4 ( .A(n353), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), .CO(
        \CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA1A S2_12_4 ( .A(n386), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), .CO(
        \CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_10_4 ( .A(n373), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_4 ( .A(n387), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_45_37 ( .A(\ab[45][37] ), .B(\CARRYB[44][37] ), .CI(\SUMB[44][38] ), 
        .CO(\CARRYB[45][37] ), .S(\SUMB[45][37] ) );
  FA1A S2_45_45 ( .A(n263), .B(\CARRYB[44][45] ), .CI(\SUMB[44][46] ), .CO(
        \CARRYB[45][45] ), .S(\SUMB[45][45] ) );
  FA1A S2_44_10 ( .A(\ab[44][10] ), .B(\CARRYB[43][10] ), .CI(\SUMB[43][11] ), 
        .CO(\CARRYB[44][10] ), .S(\SUMB[44][10] ) );
  FA1A S2_3_5 ( .A(n2310), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_11_5 ( .A(n418), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(
        \CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_9_6 ( .A(n484), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_5 ( .A(n419), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_44_38 ( .A(\ab[44][38] ), .B(\CARRYB[43][38] ), .CI(\SUMB[43][39] ), 
        .CO(\CARRYB[44][38] ), .S(\SUMB[44][38] ) );
  FA1A S3_43_46 ( .A(\ab[46][43] ), .B(\CARRYB[42][46] ), .CI(\ab[47][42] ), 
        .CO(\CARRYB[43][46] ), .S(\SUMB[43][46] ) );
  FA1A S2_33_7 ( .A(n510), .B(\CARRYB[32][7] ), .CI(\SUMB[32][8] ), .CO(
        \CARRYB[33][7] ), .S(\SUMB[33][7] ) );
  FA1A S2_8_6 ( .A(n483), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_8_7 ( .A(n518), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_7_6 ( .A(n482), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_2_8 ( .A(n336), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_42_23 ( .A(\ab[42][23] ), .B(\CARRYB[41][23] ), .CI(\SUMB[41][24] ), 
        .CO(\CARRYB[42][23] ), .S(\SUMB[42][23] ) );
  FA1A S2_39_27 ( .A(\CARRYB[38][27] ), .B(\ab[39][27] ), .CI(\SUMB[38][28] ), 
        .CO(\CARRYB[39][27] ), .S(\SUMB[39][27] ) );
  FA1A S2_42_36 ( .A(\ab[42][36] ), .B(\CARRYB[41][36] ), .CI(\SUMB[41][37] ), 
        .CO(\CARRYB[42][36] ), .S(\SUMB[42][36] ) );
  FA1A S2_43_39 ( .A(\ab[43][39] ), .B(\CARRYB[42][39] ), .CI(\SUMB[42][40] ), 
        .CO(\CARRYB[43][39] ), .S(\SUMB[43][39] ) );
  FA1A S2_43_38 ( .A(\ab[43][38] ), .B(\CARRYB[42][38] ), .CI(\SUMB[42][39] ), 
        .CO(\CARRYB[43][38] ), .S(\SUMB[43][38] ) );
  FA1A S2_14_7 ( .A(n513), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), .CO(
        \CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_42_45 ( .A(\ab[45][42] ), .B(\CARRYB[41][45] ), .CI(\SUMB[41][46] ), 
        .CO(\CARRYB[42][45] ), .S(\SUMB[42][45] ) );
  FA1A S3_41_46 ( .A(\ab[46][41] ), .B(\CARRYB[40][46] ), .CI(\ab[47][40] ), 
        .CO(\CARRYB[41][46] ), .S(\SUMB[41][46] ) );
  FA1A S2_9_8 ( .A(n552), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_8_8 ( .A(n2336), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_5_10 ( .A(n424), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), .CO(
        \CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_40_35 ( .A(\ab[40][35] ), .B(\CARRYB[39][35] ), .CI(\SUMB[39][36] ), 
        .CO(\CARRYB[40][35] ), .S(\SUMB[40][35] ) );
  FA1A S2_41_39 ( .A(\ab[41][39] ), .B(\CARRYB[40][39] ), .CI(\SUMB[40][40] ), 
        .CO(\CARRYB[41][39] ), .S(\SUMB[41][39] ) );
  FA1A S2_41_42 ( .A(\ab[42][41] ), .B(\CARRYB[40][42] ), .CI(\SUMB[40][43] ), 
        .CO(\CARRYB[41][42] ), .S(\SUMB[41][42] ) );
  FA1A S2_41_45 ( .A(\ab[45][41] ), .B(\CARRYB[40][45] ), .CI(\SUMB[40][46] ), 
        .CO(\CARRYB[41][45] ), .S(\SUMB[41][45] ) );
  FA1A S2_41_40 ( .A(\ab[41][40] ), .B(\CARRYB[40][40] ), .CI(\SUMB[40][41] ), 
        .CO(\CARRYB[41][40] ), .S(\SUMB[41][40] ) );
  FA1A S2_12_10 ( .A(n615), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), .CO(
        \CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_38_32 ( .A(\ab[38][32] ), .B(\CARRYB[37][32] ), .CI(\SUMB[37][33] ), 
        .CO(\CARRYB[38][32] ), .S(\SUMB[38][32] ) );
  FA1A S2_40_40 ( .A(n2411), .B(\CARRYB[39][40] ), .CI(\SUMB[39][41] ), .CO(
        \CARRYB[40][40] ), .S(\SUMB[40][40] ) );
  FA1A S2_11_11 ( .A(n2341), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), .CO(
        \CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_39_41 ( .A(\ab[41][39] ), .B(\CARRYB[38][41] ), .CI(\SUMB[38][42] ), 
        .CO(\CARRYB[39][41] ), .S(\SUMB[39][41] ) );
  FA1A S2_39_42 ( .A(\ab[42][39] ), .B(\CARRYB[38][42] ), .CI(\SUMB[38][43] ), 
        .CO(\CARRYB[39][42] ), .S(\SUMB[39][42] ) );
  FA1A S2_2_12 ( .A(n287), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_38_41 ( .A(\ab[41][38] ), .B(\CARRYB[37][41] ), .CI(\SUMB[37][42] ), 
        .CO(\CARRYB[38][41] ), .S(\SUMB[38][41] ) );
  FA1A S2_36_41 ( .A(\ab[41][36] ), .B(\CARRYB[35][41] ), .CI(\SUMB[35][42] ), 
        .CO(\CARRYB[36][41] ), .S(\SUMB[36][41] ) );
  FA1A S3_37_46 ( .A(\ab[46][37] ), .B(\CARRYB[36][46] ), .CI(\ab[47][36] ), 
        .CO(\CARRYB[37][46] ), .S(\SUMB[37][46] ) );
  FA1A S2_28_13 ( .A(\CARRYB[27][13] ), .B(n697), .CI(\SUMB[27][14] ), .CO(
        \CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA1A S2_9_13 ( .A(n572), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), .CO(
        \CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_35_42 ( .A(\ab[42][35] ), .B(\CARRYB[34][42] ), .CI(\SUMB[34][43] ), 
        .CO(\CARRYB[35][42] ), .S(\SUMB[35][42] ) );
  FA1A S2_36_42 ( .A(\ab[42][36] ), .B(\CARRYB[35][42] ), .CI(\SUMB[35][43] ), 
        .CO(\CARRYB[36][42] ), .S(\SUMB[36][42] ) );
  FA1A S2_37_43 ( .A(\ab[43][37] ), .B(\CARRYB[36][43] ), .CI(\SUMB[36][44] ), 
        .CO(\CARRYB[37][43] ), .S(\SUMB[37][43] ) );
  FA1A S2_37_45 ( .A(\ab[45][37] ), .B(\CARRYB[36][45] ), .CI(\SUMB[36][46] ), 
        .CO(\CARRYB[37][45] ), .S(\SUMB[37][45] ) );
  FA1A S2_37_44 ( .A(\ab[44][37] ), .B(\CARRYB[36][44] ), .CI(\SUMB[36][45] ), 
        .CO(\CARRYB[37][44] ), .S(\SUMB[37][44] ) );
  FA1A S2_32_19 ( .A(\CARRYB[31][19] ), .B(\ab[32][19] ), .CI(\SUMB[31][20] ), 
        .CO(\CARRYB[32][19] ), .S(\SUMB[32][19] ) );
  FA1A S3_36_46 ( .A(\ab[46][36] ), .B(\CARRYB[35][46] ), .CI(\ab[47][35] ), 
        .CO(\CARRYB[36][46] ), .S(\SUMB[36][46] ) );
  FA1A S2_31_16 ( .A(\CARRYB[30][16] ), .B(\ab[31][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FA1A S2_34_42 ( .A(\ab[42][34] ), .B(\CARRYB[33][42] ), .CI(\SUMB[33][43] ), 
        .CO(\CARRYB[34][42] ), .S(\SUMB[34][42] ) );
  FA1A S2_34_43 ( .A(\ab[43][34] ), .B(\CARRYB[33][43] ), .CI(\SUMB[33][44] ), 
        .CO(\CARRYB[34][43] ), .S(\SUMB[34][43] ) );
  FA1A S2_35_43 ( .A(\ab[43][35] ), .B(\CARRYB[34][43] ), .CI(\SUMB[34][44] ), 
        .CO(\CARRYB[35][43] ), .S(\SUMB[35][43] ) );
  FA1A S2_30_21 ( .A(\ab[30][21] ), .B(\CARRYB[29][21] ), .CI(\SUMB[29][22] ), 
        .CO(\CARRYB[30][21] ), .S(\SUMB[30][21] ) );
  FA1A S3_35_46 ( .A(\ab[46][35] ), .B(\CARRYB[34][46] ), .CI(\ab[47][34] ), 
        .CO(\CARRYB[35][46] ), .S(\SUMB[35][46] ) );
  FA1A S2_7_17 ( .A(\CARRYB[6][17] ), .B(n488), .CI(\SUMB[6][18] ), .CO(
        \CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1A S2_5_15 ( .A(n423), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), .CO(
        \CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_33_40 ( .A(\ab[40][33] ), .B(\CARRYB[32][40] ), .CI(\SUMB[32][41] ), 
        .CO(\CARRYB[33][40] ), .S(\SUMB[33][40] ) );
  FA1A S2_35_44 ( .A(\ab[44][35] ), .B(\CARRYB[34][44] ), .CI(\SUMB[34][45] ), 
        .CO(\CARRYB[35][44] ), .S(\SUMB[35][44] ) );
  FA1A S2_33_43 ( .A(\ab[43][33] ), .B(\CARRYB[32][43] ), .CI(\SUMB[32][44] ), 
        .CO(\CARRYB[33][43] ), .S(\SUMB[33][43] ) );
  FA1A S2_33_44 ( .A(\ab[44][33] ), .B(\CARRYB[32][44] ), .CI(\SUMB[32][45] ), 
        .CO(\CARRYB[33][44] ), .S(\SUMB[33][44] ) );
  FA1A S2_34_45 ( .A(\ab[45][34] ), .B(\CARRYB[33][45] ), .CI(\SUMB[33][46] ), 
        .CO(\CARRYB[34][45] ), .S(\SUMB[34][45] ) );
  FA1A S2_32_43 ( .A(\ab[43][32] ), .B(\CARRYB[31][43] ), .CI(\SUMB[31][44] ), 
        .CO(\CARRYB[32][43] ), .S(\SUMB[32][43] ) );
  FA1A S2_32_44 ( .A(\ab[44][32] ), .B(\CARRYB[31][44] ), .CI(\SUMB[31][45] ), 
        .CO(\CARRYB[32][44] ), .S(\SUMB[32][44] ) );
  FA1A S2_32_45 ( .A(\ab[45][32] ), .B(\CARRYB[31][45] ), .CI(\SUMB[31][46] ), 
        .CO(\CARRYB[32][45] ), .S(\SUMB[32][45] ) );
  FA1A S2_12_21 ( .A(n667), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), .CO(
        \CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA1A S2_29_42 ( .A(\ab[42][29] ), .B(\CARRYB[28][42] ), .CI(\SUMB[28][43] ), 
        .CO(\CARRYB[29][42] ), .S(\SUMB[29][42] ) );
  FA1A S2_31_45 ( .A(\ab[45][31] ), .B(\CARRYB[30][45] ), .CI(\SUMB[30][46] ), 
        .CO(\CARRYB[31][45] ), .S(\SUMB[31][45] ) );
  FA1A S3_31_46 ( .A(\ab[46][31] ), .B(\CARRYB[30][46] ), .CI(\ab[47][30] ), 
        .CO(\CARRYB[31][46] ), .S(\SUMB[31][46] ) );
  FA1A S3_32_46 ( .A(\ab[46][32] ), .B(\CARRYB[31][46] ), .CI(\ab[47][31] ), 
        .CO(\CARRYB[32][46] ), .S(\SUMB[32][46] ) );
  FA1A S2_23_31 ( .A(\CARRYB[22][31] ), .B(\ab[31][23] ), .CI(\SUMB[22][32] ), 
        .CO(\CARRYB[23][31] ), .S(\SUMB[23][31] ) );
  FA1A S3_30_46 ( .A(\ab[46][30] ), .B(\CARRYB[29][46] ), .CI(\ab[47][29] ), 
        .CO(\CARRYB[30][46] ), .S(\SUMB[30][46] ) );
  FA1A S3_29_46 ( .A(\ab[46][29] ), .B(\CARRYB[28][46] ), .CI(\ab[47][28] ), 
        .CO(\CARRYB[29][46] ), .S(\SUMB[29][46] ) );
  FA1A S2_15_23 ( .A(\CARRYB[14][23] ), .B(n716), .CI(\SUMB[14][24] ), .CO(
        \CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA1A S2_25_43 ( .A(\ab[43][25] ), .B(\CARRYB[24][43] ), .CI(\SUMB[24][44] ), 
        .CO(\CARRYB[25][43] ), .S(\SUMB[25][43] ) );
  FA1A S2_23_44 ( .A(\ab[44][23] ), .B(\CARRYB[22][44] ), .CI(\SUMB[22][45] ), 
        .CO(\CARRYB[23][44] ), .S(\SUMB[23][44] ) );
  FA1A S2_25_44 ( .A(\ab[44][25] ), .B(\CARRYB[24][44] ), .CI(\SUMB[24][45] ), 
        .CO(\CARRYB[25][44] ), .S(\SUMB[25][44] ) );
  FA1A S2_17_32 ( .A(\ab[32][17] ), .B(\CARRYB[16][32] ), .CI(\SUMB[16][33] ), 
        .CO(\CARRYB[17][32] ), .S(\SUMB[17][32] ) );
  FA1A S2_14_26 ( .A(n708), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), .CO(
        \CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA1A S2_16_34 ( .A(\ab[34][16] ), .B(\CARRYB[15][34] ), .CI(\SUMB[15][35] ), 
        .CO(\CARRYB[16][34] ), .S(\SUMB[16][34] ) );
  FA1A S3_20_46 ( .A(\ab[46][20] ), .B(\CARRYB[19][46] ), .CI(\ab[47][19] ), 
        .CO(\CARRYB[20][46] ), .S(\SUMB[20][46] ) );
  FA1A S2_11_31 ( .A(\CARRYB[10][31] ), .B(n631), .CI(\SUMB[10][32] ), .CO(
        \CARRYB[11][31] ), .S(\SUMB[11][31] ) );
  FA1A S2_10_29 ( .A(\CARRYB[9][29] ), .B(n605), .CI(\SUMB[9][30] ), .CO(
        \CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1A S3_19_46 ( .A(\ab[46][19] ), .B(\CARRYB[18][46] ), .CI(\ab[47][18] ), 
        .CO(\CARRYB[19][46] ), .S(\SUMB[19][46] ) );
  FA1A S2_5_31 ( .A(n416), .B(\CARRYB[4][31] ), .CI(\SUMB[4][32] ), .CO(
        \CARRYB[5][31] ), .S(\SUMB[5][31] ) );
  FA1A S3_18_46 ( .A(\ab[46][18] ), .B(\CARRYB[17][46] ), .CI(\ab[47][17] ), 
        .CO(\CARRYB[18][46] ), .S(\SUMB[18][46] ) );
  FA1A S2_7_33 ( .A(n510), .B(\CARRYB[6][33] ), .CI(\SUMB[6][34] ), .CO(
        \CARRYB[7][33] ), .S(\SUMB[7][33] ) );
  FA1A S2_8_39 ( .A(n547), .B(\CARRYB[7][39] ), .CI(\SUMB[7][40] ), .CO(
        \CARRYB[8][39] ), .S(\SUMB[8][39] ) );
  FA1A S2_7_37 ( .A(\CARRYB[6][37] ), .B(n472), .CI(\SUMB[6][38] ), .CO(
        \CARRYB[7][37] ), .S(\SUMB[7][37] ) );
  FA1A S2_6_37 ( .A(n440), .B(\CARRYB[5][37] ), .CI(\SUMB[5][38] ), .CO(
        \CARRYB[6][37] ), .S(\SUMB[6][37] ) );
  FA1A S2_5_2 ( .A(n2267), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_9_2 ( .A(n2254), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_29_2 ( .A(n2238), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), .CO(
        \CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA1A S2_45_18 ( .A(\ab[45][18] ), .B(\CARRYB[44][18] ), .CI(\SUMB[44][19] ), 
        .CO(\CARRYB[45][18] ), .S(\SUMB[45][18] ) );
  FA1A S2_45_5 ( .A(\CARRYB[44][5] ), .B(n394), .CI(\SUMB[44][6] ), .CO(
        \CARRYB[45][5] ), .S(\SUMB[45][5] ) );
  FA1A S2_20_5 ( .A(n402), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), .CO(
        \CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA1A S2_41_14 ( .A(\CARRYB[40][14] ), .B(\ab[41][14] ), .CI(\SUMB[40][15] ), 
        .CO(\CARRYB[41][14] ), .S(\SUMB[41][14] ) );
  FA1A S2_24_9 ( .A(\CARRYB[23][9] ), .B(n571), .CI(\SUMB[23][10] ), .CO(
        \CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA1A S2_35_33 ( .A(\ab[35][33] ), .B(\CARRYB[34][33] ), .CI(\SUMB[34][34] ), 
        .CO(\CARRYB[35][33] ), .S(\SUMB[35][33] ) );
  FA1A S2_31_17 ( .A(\CARRYB[30][17] ), .B(\ab[31][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FA1A S2_28_30 ( .A(\CARRYB[27][30] ), .B(\ab[30][28] ), .CI(\SUMB[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA1A S2_29_35 ( .A(\ab[35][29] ), .B(\CARRYB[28][35] ), .CI(\SUMB[28][36] ), 
        .CO(\CARRYB[29][35] ), .S(\SUMB[29][35] ) );
  FA1AP S2_28_39 ( .A(\ab[39][28] ), .B(\CARRYB[27][39] ), .CI(\SUMB[27][40] ), 
        .CO(\CARRYB[28][39] ), .S(\SUMB[28][39] ) );
  FA1AP S2_27_38 ( .A(\ab[38][27] ), .B(\CARRYB[26][38] ), .CI(\SUMB[26][39] ), 
        .CO(\CARRYB[27][38] ), .S(\SUMB[27][38] ) );
  FA1A S2_27_39 ( .A(\ab[39][27] ), .B(\CARRYB[26][39] ), .CI(\SUMB[26][40] ), 
        .CO(\CARRYB[27][39] ), .S(\SUMB[27][39] ) );
  FA1AP S2_26_38 ( .A(\ab[38][26] ), .B(\CARRYB[25][38] ), .CI(\SUMB[25][39] ), 
        .CO(\CARRYB[26][38] ), .S(\SUMB[26][38] ) );
  FA1A S2_20_31 ( .A(\CARRYB[19][31] ), .B(\ab[31][20] ), .CI(\SUMB[19][32] ), 
        .CO(\CARRYB[20][31] ), .S(\SUMB[20][31] ) );
  FA1A S2_13_24 ( .A(n690), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), .CO(
        \CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA1A S2_9_26 ( .A(\CARRYB[8][26] ), .B(n564), .CI(\SUMB[8][27] ), .CO(
        \CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1A S2_15_36 ( .A(\ab[36][15] ), .B(\CARRYB[14][36] ), .CI(\SUMB[14][37] ), 
        .CO(\CARRYB[15][36] ), .S(\SUMB[15][36] ) );
  FA1AP S2_13_27 ( .A(\CARRYB[12][27] ), .B(n682), .CI(\SUMB[12][28] ), .CO(
        \CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA1P S2_30_44 ( .A(\ab[44][30] ), .B(\CARRYB[29][44] ), .CI(\SUMB[29][45] ), 
        .CO(\CARRYB[30][44] ), .S(\SUMB[30][44] ) );
  FA1P S2_6_42 ( .A(n478), .B(\CARRYB[5][42] ), .CI(\SUMB[5][43] ), .CO(
        \CARRYB[6][42] ), .S(\SUMB[6][42] ) );
  FA1P S2_7_42 ( .A(n505), .B(\CARRYB[6][42] ), .CI(\SUMB[6][43] ), .CO(
        \CARRYB[7][42] ), .S(\SUMB[7][42] ) );
  FA1P S2_26_45 ( .A(\ab[45][26] ), .B(\CARRYB[25][45] ), .CI(\SUMB[25][46] ), 
        .CO(\CARRYB[26][45] ), .S(\SUMB[26][45] ) );
  FA1P S2_46_43 ( .A(\ab[46][43] ), .B(\CARRYB[45][43] ), .CI(\SUMB[45][44] ), 
        .CO(\CARRYB[46][43] ), .S(\SUMB[46][43] ) );
  FA1AP S4_43 ( .A(\ab[47][43] ), .B(\CARRYB[46][43] ), .CI(\SUMB[46][44] ), 
        .CO(\CARRYB[47][43] ), .S(\SUMB[47][43] ) );
  FA1P S2_8_45 ( .A(n521), .B(\CARRYB[7][45] ), .CI(\SUMB[7][46] ), .CO(
        \CARRYB[8][45] ), .S(\SUMB[8][45] ) );
  FA1P S2_9_45 ( .A(\ab[9][45] ), .B(\CARRYB[8][45] ), .CI(\SUMB[8][46] ), 
        .CO(\CARRYB[9][45] ), .S(\SUMB[9][45] ) );
  FA1AP S2_11_42 ( .A(\ab[42][11] ), .B(\CARRYB[10][42] ), .CI(\SUMB[10][43] ), 
        .CO(\CARRYB[11][42] ), .S(\SUMB[11][42] ) );
  FA1P S2_5_44 ( .A(\SUMB[4][45] ), .B(\CARRYB[4][44] ), .CI(n439), .CO(
        \CARRYB[5][44] ), .S(\SUMB[5][44] ) );
  FA1P S2_4_42 ( .A(n384), .B(\CARRYB[3][42] ), .CI(\SUMB[3][43] ), .CO(
        \CARRYB[4][42] ), .S(\SUMB[4][42] ) );
  FA1P S2_5_42 ( .A(n454), .B(\CARRYB[4][42] ), .CI(\SUMB[4][43] ), .CO(
        \CARRYB[5][42] ), .S(\SUMB[5][42] ) );
  FA1P S2_6_45 ( .A(n485), .B(\CARRYB[5][45] ), .CI(\SUMB[5][46] ), .CO(
        \CARRYB[6][45] ), .S(\SUMB[6][45] ) );
  FA1P S2_7_45 ( .A(n494), .B(\CARRYB[6][45] ), .CI(\SUMB[6][46] ), .CO(
        \CARRYB[7][45] ), .S(\SUMB[7][45] ) );
  FA1P S2_5_41 ( .A(n444), .B(\CARRYB[4][41] ), .CI(\SUMB[4][42] ), .CO(
        \CARRYB[5][41] ), .S(\SUMB[5][41] ) );
  FA1P S2_6_41 ( .A(n493), .B(\CARRYB[5][41] ), .CI(\SUMB[5][42] ), .CO(
        \CARRYB[6][41] ), .S(\SUMB[6][41] ) );
  FA1P S2_6_44 ( .A(n453), .B(\CARRYB[5][44] ), .CI(\SUMB[5][45] ), .CO(
        \CARRYB[6][44] ), .S(\SUMB[6][44] ) );
  FA1P S2_10_42 ( .A(\CARRYB[9][42] ), .B(\ab[42][10] ), .CI(\SUMB[9][43] ), 
        .CO(\CARRYB[10][42] ), .S(\SUMB[10][42] ) );
  FA1P S2_20_41 ( .A(\ab[41][20] ), .B(\CARRYB[19][41] ), .CI(\SUMB[19][42] ), 
        .CO(\CARRYB[20][41] ), .S(\SUMB[20][41] ) );
  FA1 S2_44_44 ( .A(n280), .B(\CARRYB[43][44] ), .CI(\SUMB[43][45] ), .CO(
        \CARRYB[44][44] ), .S(\SUMB[44][44] ) );
  FA1P S2_18_41 ( .A(\ab[41][18] ), .B(\CARRYB[17][41] ), .CI(\SUMB[17][42] ), 
        .CO(\CARRYB[18][41] ), .S(\SUMB[18][41] ) );
  FA1P S2_19_41 ( .A(\ab[41][19] ), .B(\CARRYB[18][41] ), .CI(\SUMB[18][42] ), 
        .CO(\CARRYB[19][41] ), .S(\SUMB[19][41] ) );
  FA1P S2_19_42 ( .A(\ab[42][19] ), .B(\CARRYB[18][42] ), .CI(\SUMB[18][43] ), 
        .CO(\CARRYB[19][42] ), .S(\SUMB[19][42] ) );
  FA1P S2_10_45 ( .A(\ab[45][10] ), .B(\CARRYB[9][45] ), .CI(\SUMB[9][46] ), 
        .CO(\CARRYB[10][45] ), .S(\SUMB[10][45] ) );
  FA1P S2_11_45 ( .A(\ab[45][11] ), .B(\CARRYB[10][45] ), .CI(\SUMB[10][46] ), 
        .CO(\CARRYB[11][45] ), .S(\SUMB[11][45] ) );
  FA1 S2_37_36 ( .A(\ab[37][36] ), .B(\CARRYB[36][36] ), .CI(\SUMB[36][37] ), 
        .CO(\CARRYB[37][36] ), .S(\SUMB[37][36] ) );
  FA1P S2_44_43 ( .A(\ab[44][43] ), .B(\CARRYB[43][43] ), .CI(\SUMB[43][44] ), 
        .CO(\CARRYB[44][43] ), .S(\SUMB[44][43] ) );
  FA1P S2_45_43 ( .A(\ab[45][43] ), .B(\CARRYB[44][43] ), .CI(\SUMB[44][44] ), 
        .CO(\CARRYB[45][43] ), .S(\SUMB[45][43] ) );
  FA1P S2_36_36 ( .A(n2399), .B(\CARRYB[35][36] ), .CI(\SUMB[35][37] ), .CO(
        \CARRYB[36][36] ), .S(\SUMB[36][36] ) );
  FA1P S2_16_41 ( .A(\ab[41][16] ), .B(\CARRYB[15][41] ), .CI(\SUMB[15][42] ), 
        .CO(\CARRYB[16][41] ), .S(\SUMB[16][41] ) );
  FA1P S2_16_43 ( .A(\ab[43][16] ), .B(\CARRYB[15][43] ), .CI(\SUMB[15][44] ), 
        .CO(\CARRYB[16][43] ), .S(\SUMB[16][43] ) );
  FA1P S2_38_35 ( .A(\ab[38][35] ), .B(\CARRYB[37][35] ), .CI(\SUMB[37][36] ), 
        .CO(\CARRYB[38][35] ), .S(\SUMB[38][35] ) );
  FA1 S2_39_35 ( .A(\ab[39][35] ), .B(\CARRYB[38][35] ), .CI(\SUMB[38][36] ), 
        .CO(\CARRYB[39][35] ), .S(\SUMB[39][35] ) );
  FA1P S2_14_43 ( .A(\ab[43][14] ), .B(\CARRYB[13][43] ), .CI(\SUMB[13][44] ), 
        .CO(\CARRYB[14][43] ), .S(\SUMB[14][43] ) );
  FA1P S2_34_36 ( .A(\ab[36][34] ), .B(\CARRYB[33][36] ), .CI(\SUMB[33][37] ), 
        .CO(\CARRYB[34][36] ), .S(\SUMB[34][36] ) );
  FA1P S2_35_36 ( .A(\ab[36][35] ), .B(\CARRYB[34][36] ), .CI(\SUMB[34][37] ), 
        .CO(\CARRYB[35][36] ), .S(\SUMB[35][36] ) );
  FA1P S2_14_44 ( .A(\ab[44][14] ), .B(\CARRYB[13][44] ), .CI(\SUMB[13][45] ), 
        .CO(\CARRYB[14][44] ), .S(\SUMB[14][44] ) );
  FA1AP S2_23_41 ( .A(\ab[41][23] ), .B(\CARRYB[22][41] ), .CI(\SUMB[22][42] ), 
        .CO(\CARRYB[23][41] ), .S(\SUMB[23][41] ) );
  FA1P S2_42_44 ( .A(\ab[44][42] ), .B(\CARRYB[41][44] ), .CI(\SUMB[41][45] ), 
        .CO(\CARRYB[42][44] ), .S(\SUMB[42][44] ) );
  FA1P S2_43_44 ( .A(\ab[44][43] ), .B(\CARRYB[42][44] ), .CI(\SUMB[42][45] ), 
        .CO(\CARRYB[43][44] ), .S(\SUMB[43][44] ) );
  FA1P S2_42_43 ( .A(\ab[43][42] ), .B(\CARRYB[41][43] ), .CI(\SUMB[41][44] ), 
        .CO(\CARRYB[42][43] ), .S(\SUMB[42][43] ) );
  FA1P S3_3_46 ( .A(n2282), .B(\CARRYB[2][46] ), .CI(n339), .CO(
        \CARRYB[3][46] ), .S(\SUMB[3][46] ) );
  FA1A S2_46_1 ( .A(n2196), .B(\CARRYB[45][1] ), .CI(\SUMB[45][2] ), .CO(
        \CARRYB[46][1] ), .S(\SUMB[46][1] ) );
  FA1P S2_37_35 ( .A(\ab[37][35] ), .B(\CARRYB[36][35] ), .CI(\SUMB[36][36] ), 
        .CO(\CARRYB[37][35] ), .S(\SUMB[37][35] ) );
  FA1P S2_13_45 ( .A(\ab[45][13] ), .B(\CARRYB[12][45] ), .CI(\SUMB[12][46] ), 
        .CO(\CARRYB[13][45] ), .S(\SUMB[13][45] ) );
  FA1P S2_20_42 ( .A(\ab[42][20] ), .B(\CARRYB[19][42] ), .CI(\SUMB[19][43] ), 
        .CO(\CARRYB[20][42] ), .S(\SUMB[20][42] ) );
  FA1P S2_18_44 ( .A(\ab[44][18] ), .B(\CARRYB[17][44] ), .CI(\SUMB[17][45] ), 
        .CO(\CARRYB[18][44] ), .S(\SUMB[18][44] ) );
  FA1P S2_19_44 ( .A(\ab[44][19] ), .B(\CARRYB[18][44] ), .CI(\SUMB[18][45] ), 
        .CO(\CARRYB[19][44] ), .S(\SUMB[19][44] ) );
  FA1P S2_21_41 ( .A(\ab[41][21] ), .B(\CARRYB[20][41] ), .CI(\SUMB[20][42] ), 
        .CO(\CARRYB[21][41] ), .S(\SUMB[21][41] ) );
  FA1 S2_22_41 ( .A(\ab[41][22] ), .B(\CARRYB[21][41] ), .CI(\SUMB[21][42] ), 
        .CO(\CARRYB[22][41] ), .S(\SUMB[22][41] ) );
  FA1P S2_33_36 ( .A(\CARRYB[32][36] ), .B(\ab[36][33] ), .CI(\SUMB[32][37] ), 
        .CO(\CARRYB[33][36] ), .S(\SUMB[33][36] ) );
  FA1P S2_18_43 ( .A(\ab[43][18] ), .B(\CARRYB[17][43] ), .CI(\SUMB[17][44] ), 
        .CO(\CARRYB[18][43] ), .S(\SUMB[18][43] ) );
  FA1P S2_46_41 ( .A(\ab[46][41] ), .B(\CARRYB[45][41] ), .CI(\SUMB[45][42] ), 
        .CO(\CARRYB[46][41] ), .S(\SUMB[46][41] ) );
  FA1P S4_35 ( .A(\ab[47][35] ), .B(\CARRYB[46][35] ), .CI(\SUMB[46][36] ), 
        .CO(\CARRYB[47][35] ), .S(\SUMB[47][35] ) );
  FA1P S2_43_43 ( .A(n737), .B(\CARRYB[42][43] ), .CI(\SUMB[42][44] ), .CO(
        \CARRYB[43][43] ), .S(\SUMB[43][43] ) );
  FA1P S2_44_35 ( .A(\ab[44][35] ), .B(\CARRYB[43][35] ), .CI(\SUMB[43][36] ), 
        .CO(\CARRYB[44][35] ), .S(\SUMB[44][35] ) );
  FA1P S2_45_35 ( .A(\ab[45][35] ), .B(\CARRYB[44][35] ), .CI(\SUMB[44][36] ), 
        .CO(\CARRYB[45][35] ), .S(\SUMB[45][35] ) );
  FA1 S2_44_41 ( .A(\ab[44][41] ), .B(\CARRYB[43][41] ), .CI(\SUMB[43][42] ), 
        .CO(\CARRYB[44][41] ), .S(\SUMB[44][41] ) );
  FA1AP S2_45_41 ( .A(\ab[45][41] ), .B(\CARRYB[44][41] ), .CI(\SUMB[44][42] ), 
        .CO(\CARRYB[45][41] ), .S(\SUMB[45][41] ) );
  FA1 S2_40_43 ( .A(\ab[43][40] ), .B(\CARRYB[39][43] ), .CI(\SUMB[39][44] ), 
        .CO(\CARRYB[40][43] ), .S(\SUMB[40][43] ) );
  FA1P S2_39_1 ( .A(n2221), .B(\CARRYB[38][1] ), .CI(\SUMB[38][2] ), .CO(
        \CARRYB[39][1] ), .S(\SUMB[39][1] ) );
  FA1P S2_43_33 ( .A(\ab[43][33] ), .B(\CARRYB[42][33] ), .CI(\SUMB[42][34] ), 
        .CO(\CARRYB[43][33] ), .S(\SUMB[43][33] ) );
  FA1P S2_44_33 ( .A(\ab[44][33] ), .B(\CARRYB[43][33] ), .CI(\SUMB[43][34] ), 
        .CO(\CARRYB[44][33] ), .S(\SUMB[44][33] ) );
  FA1P S2_28_45 ( .A(\ab[45][28] ), .B(\CARRYB[27][45] ), .CI(\SUMB[27][46] ), 
        .CO(\CARRYB[28][45] ), .S(\SUMB[28][45] ) );
  FA1P S2_38_2 ( .A(n2249), .B(\CARRYB[37][2] ), .CI(\SUMB[37][3] ), .CO(
        \CARRYB[38][2] ), .S(\SUMB[38][2] ) );
  FA1P S2_39_2 ( .A(n2261), .B(\CARRYB[38][2] ), .CI(\SUMB[38][3] ), .CO(
        \CARRYB[39][2] ), .S(\SUMB[39][2] ) );
  FA1P S2_27_45 ( .A(\ab[45][27] ), .B(\CARRYB[26][45] ), .CI(\SUMB[26][46] ), 
        .CO(\CARRYB[27][45] ), .S(\SUMB[27][45] ) );
  FA1P S2_24_45 ( .A(\ab[45][24] ), .B(\CARRYB[23][45] ), .CI(\SUMB[23][46] ), 
        .CO(\CARRYB[24][45] ), .S(\SUMB[24][45] ) );
  FA1P S2_25_45 ( .A(\ab[45][25] ), .B(\CARRYB[24][45] ), .CI(\SUMB[24][46] ), 
        .CO(\CARRYB[25][45] ), .S(\SUMB[25][45] ) );
  FA1P S2_40_44 ( .A(\ab[44][40] ), .B(\CARRYB[39][44] ), .CI(\SUMB[39][45] ), 
        .CO(\CARRYB[40][44] ), .S(\SUMB[40][44] ) );
  FA1P S2_41_44 ( .A(\ab[44][41] ), .B(\CARRYB[40][44] ), .CI(\SUMB[40][45] ), 
        .CO(\CARRYB[41][44] ), .S(\SUMB[41][44] ) );
  FA1P S2_39_37 ( .A(\ab[39][37] ), .B(\CARRYB[38][37] ), .CI(\SUMB[38][38] ), 
        .CO(\CARRYB[39][37] ), .S(\SUMB[39][37] ) );
  FA1A S2_40_37 ( .A(\ab[40][37] ), .B(\CARRYB[39][37] ), .CI(\SUMB[39][38] ), 
        .CO(\CARRYB[40][37] ), .S(\SUMB[40][37] ) );
  FA1P S2_31_33 ( .A(\CARRYB[30][33] ), .B(\ab[33][31] ), .CI(\SUMB[30][34] ), 
        .CO(\CARRYB[31][33] ), .S(\SUMB[31][33] ) );
  FA1P S2_32_33 ( .A(\ab[33][32] ), .B(\CARRYB[31][33] ), .CI(\SUMB[31][34] ), 
        .CO(\CARRYB[32][33] ), .S(\SUMB[32][33] ) );
  FA1 S2_9_39 ( .A(n570), .B(\CARRYB[8][39] ), .CI(\SUMB[8][40] ), .CO(
        \CARRYB[9][39] ), .S(\SUMB[9][39] ) );
  FA1P S2_33_32 ( .A(\CARRYB[32][32] ), .B(\ab[33][32] ), .CI(\SUMB[32][33] ), 
        .CO(\CARRYB[33][32] ), .S(\SUMB[33][32] ) );
  FA1P S2_34_32 ( .A(\ab[34][32] ), .B(\CARRYB[33][32] ), .CI(\SUMB[33][33] ), 
        .CO(\CARRYB[34][32] ), .S(\SUMB[34][32] ) );
  FA1 S2_12_38 ( .A(\ab[38][12] ), .B(\CARRYB[11][38] ), .CI(\SUMB[11][39] ), 
        .CO(\CARRYB[12][38] ), .S(\SUMB[12][38] ) );
  FA1 S2_13_38 ( .A(\ab[38][13] ), .B(\CARRYB[12][38] ), .CI(\SUMB[12][39] ), 
        .CO(\CARRYB[13][38] ), .S(\SUMB[13][38] ) );
  FA1P S2_42_41 ( .A(\ab[42][41] ), .B(\CARRYB[41][41] ), .CI(\SUMB[41][42] ), 
        .CO(\CARRYB[42][41] ), .S(\SUMB[42][41] ) );
  FA1AP S2_43_41 ( .A(\ab[43][41] ), .B(\CARRYB[42][41] ), .CI(\SUMB[42][42] ), 
        .CO(\CARRYB[43][41] ), .S(\SUMB[43][41] ) );
  FA1P S2_32_3 ( .A(n2283), .B(\CARRYB[31][3] ), .CI(\SUMB[31][4] ), .CO(
        \CARRYB[32][3] ), .S(\SUMB[32][3] ) );
  FA1P S2_41_43 ( .A(\ab[43][41] ), .B(\CARRYB[40][43] ), .CI(\SUMB[40][44] ), 
        .CO(\CARRYB[41][43] ), .S(\SUMB[41][43] ) );
  FA1 S2_45_40 ( .A(\ab[45][40] ), .B(\CARRYB[44][40] ), .CI(\SUMB[44][41] ), 
        .CO(\CARRYB[45][40] ), .S(\SUMB[45][40] ) );
  FA1 S2_46_40 ( .A(\ab[46][40] ), .B(\CARRYB[45][40] ), .CI(\SUMB[45][41] ), 
        .CO(\CARRYB[46][40] ), .S(\SUMB[46][40] ) );
  FA1P S2_7_40 ( .A(n492), .B(\CARRYB[6][40] ), .CI(\SUMB[6][41] ), .CO(
        \CARRYB[7][40] ), .S(\SUMB[7][40] ) );
  FA1P S2_38_44 ( .A(\ab[44][38] ), .B(\CARRYB[37][44] ), .CI(\SUMB[37][45] ), 
        .CO(\CARRYB[38][44] ), .S(\SUMB[38][44] ) );
  FA1P S2_39_44 ( .A(\ab[44][39] ), .B(\CARRYB[38][44] ), .CI(\SUMB[38][45] ), 
        .CO(\CARRYB[39][44] ), .S(\SUMB[39][44] ) );
  FA1P S2_34_37 ( .A(\ab[37][34] ), .B(\CARRYB[33][37] ), .CI(\SUMB[33][38] ), 
        .CO(\CARRYB[34][37] ), .S(\SUMB[34][37] ) );
  FA1P S2_38_17 ( .A(\ab[38][17] ), .B(\CARRYB[37][17] ), .CI(\SUMB[37][18] ), 
        .CO(\CARRYB[38][17] ), .S(\SUMB[38][17] ) );
  FA1P S2_39_43 ( .A(\ab[43][39] ), .B(\CARRYB[38][43] ), .CI(\SUMB[38][44] ), 
        .CO(\CARRYB[39][43] ), .S(\SUMB[39][43] ) );
  FA1A S2_12_37 ( .A(\ab[37][12] ), .B(\CARRYB[11][37] ), .CI(\SUMB[11][38] ), 
        .CO(\CARRYB[12][37] ), .S(\SUMB[12][37] ) );
  FA1AP S2_13_37 ( .A(\CARRYB[12][37] ), .B(\ab[37][13] ), .CI(\SUMB[12][38] ), 
        .CO(\CARRYB[13][37] ), .S(\SUMB[13][37] ) );
  FA1P S2_37_2 ( .A(n318), .B(\CARRYB[36][2] ), .CI(\SUMB[36][3] ), .CO(
        \CARRYB[37][2] ), .S(\SUMB[37][2] ) );
  FA1P S2_30_3 ( .A(n2273), .B(\CARRYB[29][3] ), .CI(\SUMB[29][4] ), .CO(
        \CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA1AP S2_10_38 ( .A(\CARRYB[9][38] ), .B(n613), .CI(\SUMB[9][39] ), .CO(
        \CARRYB[10][38] ), .S(\SUMB[10][38] ) );
  FA1P S2_11_38 ( .A(\ab[38][11] ), .B(\CARRYB[10][38] ), .CI(\SUMB[10][39] ), 
        .CO(\CARRYB[11][38] ), .S(\SUMB[11][38] ) );
  FA1P S2_30_43 ( .A(\ab[43][30] ), .B(\CARRYB[29][43] ), .CI(\SUMB[29][44] ), 
        .CO(\CARRYB[30][43] ), .S(\SUMB[30][43] ) );
  FA1AP S2_31_43 ( .A(\ab[43][31] ), .B(\CARRYB[30][43] ), .CI(\SUMB[30][44] ), 
        .CO(\CARRYB[31][43] ), .S(\SUMB[31][43] ) );
  FA1AP S2_40_39 ( .A(\ab[40][39] ), .B(\CARRYB[39][39] ), .CI(\SUMB[39][40] ), 
        .CO(\CARRYB[40][39] ), .S(\SUMB[40][39] ) );
  FA1AP S2_38_40 ( .A(\ab[40][38] ), .B(\CARRYB[37][40] ), .CI(\SUMB[37][41] ), 
        .CO(\CARRYB[38][40] ), .S(\SUMB[38][40] ) );
  FA1 S2_39_39 ( .A(n2408), .B(\CARRYB[38][39] ), .CI(\SUMB[38][40] ), .CO(
        \CARRYB[39][39] ), .S(\SUMB[39][39] ) );
  FA1P S2_36_17 ( .A(\ab[36][17] ), .B(\CARRYB[35][17] ), .CI(\SUMB[35][18] ), 
        .CO(\CARRYB[36][17] ), .S(\SUMB[36][17] ) );
  FA1P S2_37_17 ( .A(\CARRYB[36][17] ), .B(\ab[37][17] ), .CI(\SUMB[36][18] ), 
        .CO(\CARRYB[37][17] ), .S(\SUMB[37][17] ) );
  FA1 S2_40_41 ( .A(\ab[41][40] ), .B(\CARRYB[39][41] ), .CI(\SUMB[39][42] ), 
        .CO(\CARRYB[40][41] ), .S(\SUMB[40][41] ) );
  FA1AP S2_41_41 ( .A(n316), .B(\CARRYB[40][41] ), .CI(\SUMB[40][42] ), .CO(
        \CARRYB[41][41] ), .S(\SUMB[41][41] ) );
  FA1P S2_35_41 ( .A(\ab[41][35] ), .B(\CARRYB[34][41] ), .CI(\SUMB[34][42] ), 
        .CO(\CARRYB[35][41] ), .S(\SUMB[35][41] ) );
  FA1P S2_23_45 ( .A(\ab[45][23] ), .B(\CARRYB[22][45] ), .CI(\SUMB[22][46] ), 
        .CO(\CARRYB[23][45] ), .S(\SUMB[23][45] ) );
  FA1P S2_5_38 ( .A(n413), .B(\CARRYB[4][38] ), .CI(\SUMB[4][39] ), .CO(
        \CARRYB[5][38] ), .S(\SUMB[5][38] ) );
  FA1 S2_28_44 ( .A(\ab[44][28] ), .B(\CARRYB[27][44] ), .CI(\SUMB[27][45] ), 
        .CO(\CARRYB[28][44] ), .S(\SUMB[28][44] ) );
  FA1AP S2_29_44 ( .A(\ab[44][29] ), .B(\CARRYB[28][44] ), .CI(\SUMB[28][45] ), 
        .CO(\CARRYB[29][44] ), .S(\SUMB[29][44] ) );
  FA1P S2_26_3 ( .A(n2288), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), .CO(
        \CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA1P S2_27_3 ( .A(n2274), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), .CO(
        \CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA1AP S2_40_38 ( .A(\ab[40][38] ), .B(\CARRYB[39][38] ), .CI(\SUMB[39][39] ), 
        .CO(\CARRYB[40][38] ), .S(\SUMB[40][38] ) );
  FA1A S2_36_39 ( .A(\ab[39][36] ), .B(\CARRYB[35][39] ), .CI(\SUMB[35][40] ), 
        .CO(\CARRYB[36][39] ), .S(\SUMB[36][39] ) );
  FA1AP S2_34_40 ( .A(\ab[40][34] ), .B(\CARRYB[33][40] ), .CI(\SUMB[33][41] ), 
        .CO(\CARRYB[34][40] ), .S(\SUMB[34][40] ) );
  FA1 S2_35_39 ( .A(\ab[39][35] ), .B(\CARRYB[34][39] ), .CI(\SUMB[34][40] ), 
        .CO(\CARRYB[35][39] ), .S(\SUMB[35][39] ) );
  FA1P S3_27_46 ( .A(\ab[46][27] ), .B(\CARRYB[26][46] ), .CI(\ab[47][26] ), 
        .CO(\CARRYB[27][46] ), .S(\SUMB[27][46] ) );
  FA1P S2_24_2 ( .A(n2259), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), .CO(
        \CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA1 S2_25_2 ( .A(n2207), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), .CO(
        \CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA1P S2_19_3 ( .A(n2272), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), .CO(
        \CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1P S2_20_3 ( .A(n2280), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), .CO(
        \CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1P S2_21_2 ( .A(n2264), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), .CO(
        \CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1P S2_22_2 ( .A(n2263), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), .CO(
        \CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA1 S2_30_42 ( .A(\ab[42][30] ), .B(\CARRYB[29][42] ), .CI(\SUMB[29][43] ), 
        .CO(\CARRYB[30][42] ), .S(\SUMB[30][42] ) );
  FA1 S2_28_43 ( .A(\ab[43][28] ), .B(\CARRYB[27][43] ), .CI(\SUMB[27][44] ), 
        .CO(\CARRYB[28][43] ), .S(\SUMB[28][43] ) );
  FA1AP S2_29_43 ( .A(\ab[43][29] ), .B(\CARRYB[28][43] ), .CI(\SUMB[28][44] ), 
        .CO(\CARRYB[29][43] ), .S(\SUMB[29][43] ) );
  FA1P S2_35_17 ( .A(\CARRYB[34][17] ), .B(\ab[35][17] ), .CI(\SUMB[34][18] ), 
        .CO(\CARRYB[35][17] ), .S(\SUMB[35][17] ) );
  FA1P S2_4_39 ( .A(n383), .B(\CARRYB[3][39] ), .CI(\SUMB[3][40] ), .CO(
        \CARRYB[4][39] ), .S(\SUMB[4][39] ) );
  FA1 S2_29_41 ( .A(\ab[41][29] ), .B(\CARRYB[28][41] ), .CI(\SUMB[28][42] ), 
        .CO(\CARRYB[29][41] ), .S(\SUMB[29][41] ) );
  FA1A S2_30_41 ( .A(\ab[41][30] ), .B(\CARRYB[29][41] ), .CI(\SUMB[29][42] ), 
        .CO(\CARRYB[30][41] ), .S(\SUMB[30][41] ) );
  FA1P S2_17_45 ( .A(\ab[45][17] ), .B(\CARRYB[16][45] ), .CI(\SUMB[16][46] ), 
        .CO(\CARRYB[17][45] ), .S(\SUMB[17][45] ) );
  FA1P S2_18_45 ( .A(\ab[45][18] ), .B(\CARRYB[17][45] ), .CI(\SUMB[17][46] ), 
        .CO(\CARRYB[18][45] ), .S(\SUMB[18][45] ) );
  FA1P S2_13_36 ( .A(\ab[36][13] ), .B(\CARRYB[12][36] ), .CI(\SUMB[12][37] ), 
        .CO(\CARRYB[13][36] ), .S(\SUMB[13][36] ) );
  FA1A S2_6_39 ( .A(\CARRYB[5][39] ), .B(n463), .CI(\SUMB[5][40] ), .CO(
        \CARRYB[6][39] ), .S(\SUMB[6][39] ) );
  FA1P S2_31_39 ( .A(\ab[39][31] ), .B(\CARRYB[30][39] ), .CI(\SUMB[30][40] ), 
        .CO(\CARRYB[31][39] ), .S(\SUMB[31][39] ) );
  FA1P S2_32_38 ( .A(\ab[38][32] ), .B(\CARRYB[31][38] ), .CI(\SUMB[31][39] ), 
        .CO(\CARRYB[32][38] ), .S(\SUMB[32][38] ) );
  FA1AP S2_31_41 ( .A(\ab[41][31] ), .B(\CARRYB[30][41] ), .CI(\SUMB[30][42] ), 
        .CO(\CARRYB[31][41] ), .S(\SUMB[31][41] ) );
  FA1 S2_32_40 ( .A(\ab[40][32] ), .B(\CARRYB[31][40] ), .CI(\SUMB[31][41] ), 
        .CO(\CARRYB[32][40] ), .S(\SUMB[32][40] ) );
  FA1P S2_30_38 ( .A(\ab[38][30] ), .B(\CARRYB[29][38] ), .CI(\SUMB[29][39] ), 
        .CO(\CARRYB[30][38] ), .S(\SUMB[30][38] ) );
  FA1P S2_31_38 ( .A(\ab[38][31] ), .B(\CARRYB[30][38] ), .CI(\SUMB[30][39] ), 
        .CO(\CARRYB[31][38] ), .S(\SUMB[31][38] ) );
  FA1AP S2_28_42 ( .A(\ab[42][28] ), .B(\CARRYB[27][42] ), .CI(\SUMB[27][43] ), 
        .CO(\CARRYB[28][42] ), .S(\SUMB[28][42] ) );
  FA1P S2_16_44 ( .A(\ab[44][16] ), .B(\CARRYB[15][44] ), .CI(\SUMB[15][45] ), 
        .CO(\CARRYB[16][44] ), .S(\SUMB[16][44] ) );
  FA1P S3_25_46 ( .A(\ab[46][25] ), .B(\CARRYB[24][46] ), .CI(\ab[47][24] ), 
        .CO(\CARRYB[25][46] ), .S(\SUMB[25][46] ) );
  FA1P S3_26_46 ( .A(\ab[46][26] ), .B(\CARRYB[25][46] ), .CI(\ab[47][25] ), 
        .CO(\CARRYB[26][46] ), .S(\SUMB[26][46] ) );
  FA1P S2_28_34 ( .A(\CARRYB[27][34] ), .B(\ab[34][28] ), .CI(\SUMB[27][35] ), 
        .CO(\CARRYB[28][34] ), .S(\SUMB[28][34] ) );
  FA1P S2_28_41 ( .A(\ab[41][28] ), .B(\CARRYB[27][41] ), .CI(\SUMB[27][42] ), 
        .CO(\CARRYB[28][41] ), .S(\SUMB[28][41] ) );
  FA1P S2_45_13 ( .A(\CARRYB[44][13] ), .B(\ab[45][13] ), .CI(\SUMB[44][14] ), 
        .CO(\CARRYB[45][13] ), .S(\SUMB[45][13] ) );
  FA1P S2_33_37 ( .A(\ab[37][33] ), .B(\CARRYB[32][37] ), .CI(\SUMB[32][38] ), 
        .CO(\CARRYB[33][37] ), .S(\SUMB[33][37] ) );
  FA1AP S2_27_18 ( .A(\CARRYB[26][18] ), .B(\ab[27][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA1P S2_31_36 ( .A(\ab[36][31] ), .B(\CARRYB[30][36] ), .CI(\SUMB[30][37] ), 
        .CO(\CARRYB[31][36] ), .S(\SUMB[31][36] ) );
  FA1 S2_18_22 ( .A(\ab[22][18] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA1P S2_19_22 ( .A(\CARRYB[18][22] ), .B(\ab[22][19] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA1P S2_14_5 ( .A(n417), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(
        \CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1P S2_16_45 ( .A(\ab[45][16] ), .B(\CARRYB[15][45] ), .CI(\SUMB[15][46] ), 
        .CO(\CARRYB[16][45] ), .S(\SUMB[16][45] ) );
  FA1 S2_26_44 ( .A(\ab[44][26] ), .B(\CARRYB[25][44] ), .CI(\SUMB[25][45] ), 
        .CO(\CARRYB[26][44] ), .S(\SUMB[26][44] ) );
  FA1AP S2_27_44 ( .A(\ab[44][27] ), .B(\CARRYB[26][44] ), .CI(\SUMB[26][45] ), 
        .CO(\CARRYB[27][44] ), .S(\SUMB[27][44] ) );
  FA1P S2_17_4 ( .A(n371), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), .CO(
        \CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1P S2_36_1 ( .A(n2197), .B(\CARRYB[35][1] ), .CI(\SUMB[35][2] ), .CO(
        \CARRYB[36][1] ), .S(\SUMB[36][1] ) );
  FA1 S2_37_1 ( .A(n15), .B(\CARRYB[36][1] ), .CI(\SUMB[36][2] ), .CO(
        \CARRYB[37][1] ), .S(\SUMB[37][1] ) );
  FA1P S2_29_32 ( .A(\ab[32][29] ), .B(\CARRYB[28][32] ), .CI(\SUMB[28][33] ), 
        .CO(\CARRYB[29][32] ), .S(\SUMB[29][32] ) );
  FA1AP S2_36_31 ( .A(\ab[36][31] ), .B(\CARRYB[35][31] ), .CI(\SUMB[35][32] ), 
        .CO(\CARRYB[36][31] ), .S(\SUMB[36][31] ) );
  FA1AP S2_4_40 ( .A(n414), .B(\CARRYB[3][40] ), .CI(\SUMB[3][41] ), .CO(
        \CARRYB[4][40] ), .S(\SUMB[4][40] ) );
  FA1A S2_2_41 ( .A(n2251), .B(\CARRYB[1][41] ), .CI(\SUMB[1][42] ), .CO(
        \CARRYB[2][41] ), .S(\SUMB[2][41] ) );
  FA1P S2_30_39 ( .A(\ab[39][30] ), .B(\CARRYB[29][39] ), .CI(\SUMB[29][40] ), 
        .CO(\CARRYB[30][39] ), .S(\SUMB[30][39] ) );
  FA1P S2_18_3 ( .A(n2278), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), .CO(
        \CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1P S2_19_2 ( .A(n2215), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), .CO(
        \CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1P S2_20_2 ( .A(n2176), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), .CO(
        \CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA1P S1_37_0 ( .A(n320), .B(\CARRYB[36][0] ), .CI(\SUMB[36][1] ), .CO(
        \CARRYB[37][0] ), .S(\A1[35] ) );
  FA1P S1_38_0 ( .A(n2226), .B(\CARRYB[37][0] ), .CI(\SUMB[37][1] ), .CO(
        \CARRYB[38][0] ), .S(\A1[36] ) );
  FA1 S2_25_42 ( .A(\ab[42][25] ), .B(\CARRYB[24][42] ), .CI(\SUMB[24][43] ), 
        .CO(\CARRYB[25][42] ), .S(\SUMB[25][42] ) );
  FA1 S2_20_44 ( .A(\ab[44][20] ), .B(\CARRYB[19][44] ), .CI(\SUMB[19][45] ), 
        .CO(\CARRYB[20][44] ), .S(\SUMB[20][44] ) );
  FA1AP S2_21_44 ( .A(\ab[44][21] ), .B(\CARRYB[20][44] ), .CI(\SUMB[20][45] ), 
        .CO(\CARRYB[21][44] ), .S(\SUMB[21][44] ) );
  FA1P S2_25_34 ( .A(\CARRYB[24][34] ), .B(\ab[34][25] ), .CI(\SUMB[24][35] ), 
        .CO(\CARRYB[25][34] ), .S(\SUMB[25][34] ) );
  FA1P S2_26_34 ( .A(\ab[34][26] ), .B(\CARRYB[25][34] ), .CI(\SUMB[25][35] ), 
        .CO(\CARRYB[26][34] ), .S(\SUMB[26][34] ) );
  FA1P S2_21_43 ( .A(\ab[43][21] ), .B(\CARRYB[20][43] ), .CI(\SUMB[20][44] ), 
        .CO(\CARRYB[21][43] ), .S(\SUMB[21][43] ) );
  FA1P S2_15_6 ( .A(n449), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(
        \CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA1P S2_16_6 ( .A(n445), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), .CO(
        \CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1P S2_10_41 ( .A(\ab[41][10] ), .B(\CARRYB[9][41] ), .CI(\SUMB[9][42] ), 
        .CO(\CARRYB[10][41] ), .S(\SUMB[10][41] ) );
  FA1P S2_46_36 ( .A(\ab[46][36] ), .B(\CARRYB[45][36] ), .CI(\SUMB[45][37] ), 
        .CO(\CARRYB[46][36] ), .S(\SUMB[46][36] ) );
  FA1AP S4_36 ( .A(\ab[47][36] ), .B(\CARRYB[46][36] ), .CI(\SUMB[46][37] ), 
        .CO(\CARRYB[47][36] ), .S(\SUMB[47][36] ) );
  FA1AP S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA1P S2_4_25 ( .A(n364), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), .CO(
        \CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1 S2_5_25 ( .A(n404), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), .CO(
        \CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1P S2_30_1 ( .A(n2167), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), .CO(
        \CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA1P S3_23_46 ( .A(\ab[46][23] ), .B(\CARRYB[22][46] ), .CI(\ab[47][22] ), 
        .CO(\CARRYB[23][46] ), .S(\SUMB[23][46] ) );
  FA1P S3_24_46 ( .A(\ab[46][24] ), .B(\CARRYB[23][46] ), .CI(\ab[47][23] ), 
        .CO(\CARRYB[24][46] ), .S(\SUMB[24][46] ) );
  FA1P S2_26_41 ( .A(\ab[41][26] ), .B(\CARRYB[25][41] ), .CI(\SUMB[25][42] ), 
        .CO(\CARRYB[26][41] ), .S(\SUMB[26][41] ) );
  FA1P S2_42_35 ( .A(\ab[42][35] ), .B(\CARRYB[41][35] ), .CI(\SUMB[41][36] ), 
        .CO(\CARRYB[42][35] ), .S(\SUMB[42][35] ) );
  FA1P S2_43_35 ( .A(\ab[43][35] ), .B(\CARRYB[42][35] ), .CI(\SUMB[42][36] ), 
        .CO(\CARRYB[43][35] ), .S(\SUMB[43][35] ) );
  FA1P S2_14_45 ( .A(\ab[45][14] ), .B(\CARRYB[13][45] ), .CI(\SUMB[13][46] ), 
        .CO(\CARRYB[14][45] ), .S(\SUMB[14][45] ) );
  FA1P S2_15_45 ( .A(\ab[45][15] ), .B(\CARRYB[14][45] ), .CI(\SUMB[14][46] ), 
        .CO(\CARRYB[15][45] ), .S(\SUMB[15][45] ) );
  FA1P S2_17_3 ( .A(n2279), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), .CO(
        \CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1P S2_21_42 ( .A(\ab[42][21] ), .B(\CARRYB[20][42] ), .CI(\SUMB[20][43] ), 
        .CO(\CARRYB[21][42] ), .S(\SUMB[21][42] ) );
  FA1P S2_17_44 ( .A(\ab[44][17] ), .B(\CARRYB[16][44] ), .CI(\SUMB[16][45] ), 
        .CO(\CARRYB[17][44] ), .S(\SUMB[17][44] ) );
  FA1AP S4_31 ( .A(\ab[47][31] ), .B(\CARRYB[46][31] ), .CI(\SUMB[46][32] ), 
        .CO(\CARRYB[47][31] ), .S(\SUMB[47][31] ) );
  FA1P S2_15_5 ( .A(n423), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1P S2_16_4 ( .A(n359), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), .CO(
        \CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1AP S4_37 ( .A(\ab[47][37] ), .B(\CARRYB[46][37] ), .CI(\SUMB[46][38] ), 
        .CO(\CARRYB[47][37] ), .S(\SUMB[47][37] ) );
  FA1AP S2_27_43 ( .A(\ab[43][27] ), .B(\CARRYB[26][43] ), .CI(\SUMB[26][44] ), 
        .CO(\CARRYB[27][43] ), .S(\SUMB[27][43] ) );
  FA1P S2_12_5 ( .A(n405), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), .CO(
        \CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1P S2_12_6 ( .A(n466), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), .CO(
        \CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1P S2_13_5 ( .A(n422), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), .CO(
        \CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1P S2_30_16 ( .A(\CARRYB[29][16] ), .B(\ab[30][16] ), .CI(\SUMB[29][17] ), 
        .CO(\CARRYB[30][16] ), .S(\SUMB[30][16] ) );
  FA1P S2_44_36 ( .A(\ab[44][36] ), .B(\CARRYB[43][36] ), .CI(\SUMB[43][37] ), 
        .CO(\CARRYB[44][36] ), .S(\SUMB[44][36] ) );
  FA1P S2_45_36 ( .A(\ab[45][36] ), .B(\CARRYB[44][36] ), .CI(\SUMB[44][37] ), 
        .CO(\CARRYB[45][36] ), .S(\SUMB[45][36] ) );
  FA1 S2_4_24 ( .A(n365), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), .CO(
        \CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1P S2_15_4 ( .A(n367), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1 S2_35_29 ( .A(\ab[35][29] ), .B(\CARRYB[34][29] ), .CI(\SUMB[34][30] ), 
        .CO(\CARRYB[35][29] ), .S(\SUMB[35][29] ) );
  FA1P S2_44_37 ( .A(\ab[44][37] ), .B(\CARRYB[43][37] ), .CI(\SUMB[43][38] ), 
        .CO(\CARRYB[44][37] ), .S(\SUMB[44][37] ) );
  FA1P S2_22_38 ( .A(\SUMB[21][39] ), .B(\CARRYB[21][38] ), .CI(\ab[38][22] ), 
        .CO(\CARRYB[22][38] ), .S(\SUMB[22][38] ) );
  FA1P S2_23_38 ( .A(\ab[38][23] ), .B(\CARRYB[22][38] ), .CI(\SUMB[22][39] ), 
        .CO(\CARRYB[23][38] ), .S(\SUMB[23][38] ) );
  FA1 S2_28_1 ( .A(n2186), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), .CO(
        \CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA1P S2_46_38 ( .A(\ab[46][38] ), .B(\CARRYB[45][38] ), .CI(\SUMB[45][39] ), 
        .CO(\CARRYB[46][38] ), .S(\SUMB[46][38] ) );
  FA1AP S4_38 ( .A(\ab[47][38] ), .B(\CARRYB[46][38] ), .CI(\SUMB[46][39] ), 
        .CO(\CARRYB[47][38] ), .S(\SUMB[47][38] ) );
  FA1P S2_19_1 ( .A(n2165), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), .CO(
        \CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1P S2_45_12 ( .A(\CARRYB[44][12] ), .B(\ab[45][12] ), .CI(\SUMB[44][13] ), 
        .CO(\CARRYB[45][12] ), .S(\SUMB[45][12] ) );
  FA1P S2_45_16 ( .A(\ab[45][16] ), .B(\CARRYB[44][16] ), .CI(\SUMB[44][17] ), 
        .CO(\CARRYB[45][16] ), .S(\SUMB[45][16] ) );
  FA1 S2_43_23 ( .A(\ab[43][23] ), .B(\CARRYB[42][23] ), .CI(\SUMB[42][24] ), 
        .CO(\CARRYB[43][23] ), .S(\SUMB[43][23] ) );
  FA1P S2_34_41 ( .A(\ab[41][34] ), .B(\CARRYB[33][41] ), .CI(\SUMB[33][42] ), 
        .CO(\CARRYB[34][41] ), .S(\SUMB[34][41] ) );
  FA1P S2_35_40 ( .A(\ab[40][35] ), .B(\CARRYB[34][40] ), .CI(\SUMB[34][41] ), 
        .CO(\CARRYB[35][40] ), .S(\SUMB[35][40] ) );
  FA1 S2_30_17 ( .A(\ab[30][17] ), .B(\CARRYB[29][17] ), .CI(\SUMB[29][18] ), 
        .CO(\CARRYB[30][17] ), .S(\SUMB[30][17] ) );
  FA1AP S2_16_36 ( .A(\ab[36][16] ), .B(\CARRYB[15][36] ), .CI(\SUMB[15][37] ), 
        .CO(\CARRYB[16][36] ), .S(\SUMB[16][36] ) );
  FA1 S2_17_36 ( .A(\ab[36][17] ), .B(\CARRYB[16][36] ), .CI(\SUMB[16][37] ), 
        .CO(\CARRYB[17][36] ), .S(\SUMB[17][36] ) );
  FA1A S2_18_24 ( .A(\CARRYB[17][24] ), .B(\ab[24][18] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA1AP S2_16_26 ( .A(\ab[26][16] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA1AP S2_16_25 ( .A(\CARRYB[15][25] ), .B(\ab[25][16] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA1P S2_23_5 ( .A(n408), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), .CO(
        \CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA1A S2_33_42 ( .A(\ab[42][33] ), .B(\CARRYB[32][42] ), .CI(\SUMB[32][43] ), 
        .CO(\CARRYB[33][42] ), .S(\SUMB[33][42] ) );
  FA1 S2_31_42 ( .A(\ab[42][31] ), .B(\CARRYB[30][42] ), .CI(\SUMB[30][43] ), 
        .CO(\CARRYB[31][42] ), .S(\SUMB[31][42] ) );
  FA1AP S2_13_3 ( .A(n2287), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), .CO(
        \CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S1_16_0 ( .A(n269), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), .CO(
        \CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S2_14_1 ( .A(n2241), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(
        \CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1 S1_14_0 ( .A(n286), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(
        \CARRYB[14][0] ), .S(\A1[12] ) );
  FA1AP S2_39_17 ( .A(\ab[39][17] ), .B(\CARRYB[38][17] ), .CI(\SUMB[38][18] ), 
        .CO(\CARRYB[39][17] ), .S(\SUMB[39][17] ) );
  FA1A S2_37_18 ( .A(\CARRYB[36][18] ), .B(\ab[37][18] ), .CI(\SUMB[36][19] ), 
        .CO(\CARRYB[37][18] ), .S(\SUMB[37][18] ) );
  FA1P S2_10_28 ( .A(\CARRYB[9][28] ), .B(n610), .CI(\SUMB[9][29] ), .CO(
        \CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1P S2_20_40 ( .A(\ab[40][20] ), .B(\CARRYB[19][40] ), .CI(\SUMB[19][41] ), 
        .CO(\CARRYB[20][40] ), .S(\SUMB[20][40] ) );
  FA1AP S2_34_17 ( .A(\CARRYB[33][17] ), .B(\ab[34][17] ), .CI(\SUMB[33][18] ), 
        .CO(\CARRYB[34][17] ), .S(\SUMB[34][17] ) );
  FA1AP S2_13_34 ( .A(\CARRYB[12][34] ), .B(\ab[34][13] ), .CI(\SUMB[12][35] ), 
        .CO(\CARRYB[13][34] ), .S(\SUMB[13][34] ) );
  FA1A S2_46_37 ( .A(\ab[46][37] ), .B(\CARRYB[45][37] ), .CI(\SUMB[45][38] ), 
        .CO(\CARRYB[46][37] ), .S(\SUMB[46][37] ) );
  FA1AP S2_44_39 ( .A(\ab[44][39] ), .B(\CARRYB[43][39] ), .CI(\SUMB[43][40] ), 
        .CO(\CARRYB[44][39] ), .S(\SUMB[44][39] ) );
  FA1P S2_24_43 ( .A(\ab[43][24] ), .B(\CARRYB[23][43] ), .CI(\SUMB[23][44] ), 
        .CO(\CARRYB[24][43] ), .S(\SUMB[24][43] ) );
  FA1P S2_22_44 ( .A(\ab[44][22] ), .B(\CARRYB[21][44] ), .CI(\SUMB[21][45] ), 
        .CO(\CARRYB[22][44] ), .S(\SUMB[22][44] ) );
  FA1P S2_22_43 ( .A(\ab[43][22] ), .B(\CARRYB[21][43] ), .CI(\SUMB[21][44] ), 
        .CO(\CARRYB[22][43] ), .S(\SUMB[22][43] ) );
  FA1A S2_10_33 ( .A(\CARRYB[9][33] ), .B(n614), .CI(\SUMB[9][34] ), .CO(
        \CARRYB[10][33] ), .S(\SUMB[10][33] ) );
  FA1 S2_33_20 ( .A(\ab[33][20] ), .B(\CARRYB[32][20] ), .CI(\SUMB[32][21] ), 
        .CO(\CARRYB[33][20] ), .S(\SUMB[33][20] ) );
  FA1 S2_26_31 ( .A(\ab[31][26] ), .B(\CARRYB[25][31] ), .CI(\SUMB[25][32] ), 
        .CO(\CARRYB[26][31] ), .S(\SUMB[26][31] ) );
  FA1A S2_41_16 ( .A(\CARRYB[40][16] ), .B(\ab[41][16] ), .CI(\SUMB[40][17] ), 
        .CO(\CARRYB[41][16] ), .S(\SUMB[41][16] ) );
  FA1AP S2_45_24 ( .A(\ab[45][24] ), .B(\CARRYB[44][24] ), .CI(\SUMB[44][25] ), 
        .CO(\CARRYB[45][24] ), .S(\SUMB[45][24] ) );
  FA1AP S2_14_27 ( .A(n712), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), .CO(
        \CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA1A S2_32_34 ( .A(\ab[34][32] ), .B(\CARRYB[31][34] ), .CI(\SUMB[31][35] ), 
        .CO(\CARRYB[32][34] ), .S(\SUMB[32][34] ) );
  FA1AP S2_30_35 ( .A(\ab[35][30] ), .B(\CARRYB[29][35] ), .CI(\SUMB[29][36] ), 
        .CO(\CARRYB[30][35] ), .S(\SUMB[30][35] ) );
  FA1 S2_26_35 ( .A(\ab[35][26] ), .B(\CARRYB[25][35] ), .CI(\SUMB[25][36] ), 
        .CO(\CARRYB[26][35] ), .S(\SUMB[26][35] ) );
  FA1P S3_21_46 ( .A(\ab[46][21] ), .B(\CARRYB[20][46] ), .CI(\ab[47][20] ), 
        .CO(\CARRYB[21][46] ), .S(\SUMB[21][46] ) );
  FA1P S2_14_22 ( .A(\CARRYB[13][22] ), .B(n700), .CI(\SUMB[13][23] ), .CO(
        \CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA1P S2_28_40 ( .A(\ab[40][28] ), .B(\CARRYB[27][40] ), .CI(\SUMB[27][41] ), 
        .CO(\CARRYB[28][40] ), .S(\SUMB[28][40] ) );
  FA1AP S2_24_22 ( .A(\CARRYB[23][22] ), .B(\ab[24][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA1AP S2_6_40 ( .A(n458), .B(\CARRYB[5][40] ), .CI(\SUMB[5][41] ), .CO(
        \CARRYB[6][40] ), .S(\SUMB[6][40] ) );
  FA1AP S2_4_41 ( .A(\CARRYB[3][41] ), .B(n379), .CI(\SUMB[3][42] ), .CO(
        \CARRYB[4][41] ), .S(\SUMB[4][41] ) );
  FA1AP S2_6_28 ( .A(n447), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), .CO(
        \CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1 S2_2_31 ( .A(n2198), .B(\CARRYB[1][31] ), .CI(\SUMB[1][32] ), .CO(
        \CARRYB[2][31] ), .S(\SUMB[2][31] ) );
  FA1P S2_45_32 ( .A(\ab[45][32] ), .B(\CARRYB[44][32] ), .CI(\SUMB[44][33] ), 
        .CO(\CARRYB[45][32] ), .S(\SUMB[45][32] ) );
  FA1P S2_32_32 ( .A(\CARRYB[31][32] ), .B(n2389), .CI(\SUMB[31][33] ), .CO(
        \CARRYB[32][32] ), .S(\SUMB[32][32] ) );
  FA1P S2_7_44 ( .A(n486), .B(\CARRYB[6][44] ), .CI(\SUMB[6][45] ), .CO(
        \CARRYB[7][44] ), .S(\SUMB[7][44] ) );
  FA1P S2_15_44 ( .A(\ab[44][15] ), .B(\CARRYB[14][44] ), .CI(\SUMB[14][45] ), 
        .CO(\CARRYB[15][44] ), .S(\SUMB[15][44] ) );
  FA1P S2_42_38 ( .A(\ab[42][38] ), .B(\CARRYB[41][38] ), .CI(\SUMB[41][39] ), 
        .CO(\CARRYB[42][38] ), .S(\SUMB[42][38] ) );
  FA1P S2_26_42 ( .A(\ab[42][26] ), .B(\CARRYB[25][42] ), .CI(\SUMB[25][43] ), 
        .CO(\CARRYB[26][42] ), .S(\SUMB[26][42] ) );
  FA1P S2_27_42 ( .A(\ab[42][27] ), .B(\CARRYB[26][42] ), .CI(\SUMB[26][43] ), 
        .CO(\CARRYB[27][42] ), .S(\SUMB[27][42] ) );
  FA1P S2_2_9 ( .A(n2254), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1P S2_3_9 ( .A(n2298), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1P S2_15_7 ( .A(n475), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1P S2_16_7 ( .A(n479), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), .CO(
        \CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1 S2_10_7 ( .A(n528), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1P S2_11_7 ( .A(n504), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(
        \CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1AP S2_24_3 ( .A(n2289), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), .CO(
        \CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA1P S2_3_44 ( .A(n2285), .B(\CARRYB[2][44] ), .CI(\SUMB[2][45] ), .CO(
        \CARRYB[3][44] ), .S(\SUMB[3][44] ) );
  FA1P S2_43_32 ( .A(\ab[43][32] ), .B(\CARRYB[42][32] ), .CI(\SUMB[42][33] ), 
        .CO(\CARRYB[43][32] ), .S(\SUMB[43][32] ) );
  FA1P S2_27_37 ( .A(\ab[37][27] ), .B(\CARRYB[26][37] ), .CI(\SUMB[26][38] ), 
        .CO(\CARRYB[27][37] ), .S(\SUMB[27][37] ) );
  FA1AP S2_5_30 ( .A(n392), .B(\CARRYB[4][30] ), .CI(\SUMB[4][31] ), .CO(
        \CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA1P S2_19_24 ( .A(\CARRYB[18][24] ), .B(\ab[24][19] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA1P S2_31_20 ( .A(\CARRYB[30][20] ), .B(\ab[31][20] ), .CI(\SUMB[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FA1AP S2_32_20 ( .A(\ab[32][20] ), .B(\CARRYB[31][20] ), .CI(\SUMB[31][21] ), 
        .CO(\CARRYB[32][20] ), .S(\SUMB[32][20] ) );
  FA1AP S2_7_29 ( .A(n502), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), .CO(
        \CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1P S2_21_23 ( .A(\ab[23][21] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA1P S2_27_41 ( .A(\ab[41][27] ), .B(\CARRYB[26][41] ), .CI(\SUMB[26][42] ), 
        .CO(\CARRYB[27][41] ), .S(\SUMB[27][41] ) );
  FA1P S2_24_41 ( .A(\ab[41][24] ), .B(\CARRYB[23][41] ), .CI(\SUMB[23][42] ), 
        .CO(\CARRYB[24][41] ), .S(\SUMB[24][41] ) );
  FA1P S2_25_41 ( .A(\ab[41][25] ), .B(\CARRYB[24][41] ), .CI(\SUMB[24][42] ), 
        .CO(\CARRYB[25][41] ), .S(\SUMB[25][41] ) );
  FA1AP S2_42_37 ( .A(\ab[42][37] ), .B(\CARRYB[41][37] ), .CI(\SUMB[41][38] ), 
        .CO(\CARRYB[42][37] ), .S(\SUMB[42][37] ) );
  FA1P S2_43_37 ( .A(\ab[43][37] ), .B(\CARRYB[42][37] ), .CI(\SUMB[42][38] ), 
        .CO(\CARRYB[43][37] ), .S(\SUMB[43][37] ) );
  FA1P S2_30_33 ( .A(\ab[33][30] ), .B(\CARRYB[29][33] ), .CI(\SUMB[29][34] ), 
        .CO(\CARRYB[30][33] ), .S(\SUMB[30][33] ) );
  FA1 S2_45_28 ( .A(\SUMB[44][29] ), .B(\CARRYB[44][28] ), .CI(\ab[45][28] ), 
        .CO(\CARRYB[45][28] ), .S(\SUMB[45][28] ) );
  FA1P S2_39_30 ( .A(\CARRYB[38][30] ), .B(\ab[39][30] ), .CI(\SUMB[38][31] ), 
        .CO(\CARRYB[39][30] ), .S(\SUMB[39][30] ) );
  FA1 S2_9_3 ( .A(n2298), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1 S2_10_3 ( .A(n355), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S1_18_0 ( .A(n2228), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), .CO(
        \CARRYB[18][0] ), .S(\A1[16] ) );
  FA1P S1_19_0 ( .A(n2190), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), .CO(
        \CARRYB[19][0] ), .S(\A1[17] ) );
  FA1P S1_26_0 ( .A(n2182), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), .CO(
        \CARRYB[26][0] ), .S(\A1[24] ) );
  FA1 S1_22_0 ( .A(n2316), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), .CO(
        \CARRYB[22][0] ), .S(\A1[20] ) );
  FA1 S2_22_1 ( .A(n2223), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), .CO(
        \CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA1 S4_1 ( .A(n2245), .B(\CARRYB[46][1] ), .CI(\SUMB[46][2] ), .CO(
        \CARRYB[47][1] ), .S(\SUMB[47][1] ) );
  FA1AP S2_4_23 ( .A(\CARRYB[3][23] ), .B(n353), .CI(\SUMB[3][24] ), .CO(
        \CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA1AP S2_40_9 ( .A(n593), .B(\CARRYB[39][9] ), .CI(\SUMB[39][10] ), .CO(
        \CARRYB[40][9] ), .S(\SUMB[40][9] ) );
  FA1AP S2_6_22 ( .A(\CARRYB[5][22] ), .B(n441), .CI(\SUMB[5][23] ), .CO(
        \CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA1 S2_7_22 ( .A(n506), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), .CO(
        \CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA1AP S2_31_30 ( .A(\ab[31][30] ), .B(\CARRYB[30][30] ), .CI(\SUMB[30][31] ), 
        .CO(\CARRYB[31][30] ), .S(\SUMB[31][30] ) );
  FA1P S2_32_29 ( .A(\CARRYB[31][29] ), .B(\ab[32][29] ), .CI(\SUMB[31][30] ), 
        .CO(\CARRYB[32][29] ), .S(\SUMB[32][29] ) );
  FA1P S2_39_28 ( .A(\ab[39][28] ), .B(\CARRYB[38][28] ), .CI(\SUMB[38][29] ), 
        .CO(\CARRYB[39][28] ), .S(\SUMB[39][28] ) );
  FA1 S2_14_37 ( .A(\CARRYB[13][37] ), .B(\ab[37][14] ), .CI(\SUMB[13][38] ), 
        .CO(\CARRYB[14][37] ), .S(\SUMB[14][37] ) );
  FA1P S2_30_30 ( .A(\CARRYB[29][30] ), .B(n2382), .CI(\SUMB[29][31] ), .CO(
        \CARRYB[30][30] ), .S(\SUMB[30][30] ) );
  FA1 S2_28_31 ( .A(\ab[31][28] ), .B(\CARRYB[27][31] ), .CI(\SUMB[27][32] ), 
        .CO(\CARRYB[28][31] ), .S(\SUMB[28][31] ) );
  FA1P S2_29_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA1P S2_17_21 ( .A(\CARRYB[16][21] ), .B(\ab[21][17] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA1P S2_14_23 ( .A(\CARRYB[13][23] ), .B(n693), .CI(\SUMB[13][24] ), .CO(
        \CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA1P S2_37_34 ( .A(\ab[37][34] ), .B(\CARRYB[36][34] ), .CI(\SUMB[36][35] ), 
        .CO(\CARRYB[37][34] ), .S(\SUMB[37][34] ) );
  FA1P S2_12_42 ( .A(\ab[42][12] ), .B(\CARRYB[11][42] ), .CI(\SUMB[11][43] ), 
        .CO(\CARRYB[12][42] ), .S(\SUMB[12][42] ) );
  FA1P S2_39_34 ( .A(\ab[39][34] ), .B(\CARRYB[38][34] ), .CI(\SUMB[38][35] ), 
        .CO(\CARRYB[39][34] ), .S(\SUMB[39][34] ) );
  FA1P S2_41_27 ( .A(\CARRYB[40][27] ), .B(\ab[41][27] ), .CI(\SUMB[40][28] ), 
        .CO(\CARRYB[41][27] ), .S(\SUMB[41][27] ) );
  FA1 S2_26_32 ( .A(\ab[32][26] ), .B(\CARRYB[25][32] ), .CI(\SUMB[25][33] ), 
        .CO(\CARRYB[26][32] ), .S(\SUMB[26][32] ) );
  FA1P S2_5_45 ( .A(n394), .B(\CARRYB[4][45] ), .CI(\SUMB[4][46] ), .CO(
        \CARRYB[5][45] ), .S(\SUMB[5][45] ) );
  FA1P S2_20_45 ( .A(\ab[45][20] ), .B(\CARRYB[19][45] ), .CI(\SUMB[19][46] ), 
        .CO(\CARRYB[20][45] ), .S(\SUMB[20][45] ) );
  FA1P S2_21_45 ( .A(\ab[45][21] ), .B(\CARRYB[20][45] ), .CI(\SUMB[20][46] ), 
        .CO(\CARRYB[21][45] ), .S(\SUMB[21][45] ) );
  FA1P S2_46_45 ( .A(\ab[46][45] ), .B(\CARRYB[45][45] ), .CI(\SUMB[45][46] ), 
        .CO(\CARRYB[46][45] ), .S(\SUMB[46][45] ) );
  FA1 S2_30_45 ( .A(\ab[45][30] ), .B(\CARRYB[29][45] ), .CI(\SUMB[29][46] ), 
        .CO(\CARRYB[30][45] ), .S(\SUMB[30][45] ) );
  FA1P S3_28_46 ( .A(\ab[46][28] ), .B(\CARRYB[27][46] ), .CI(\ab[47][27] ), 
        .CO(\CARRYB[28][46] ), .S(\SUMB[28][46] ) );
  FA1P S2_29_45 ( .A(\ab[45][29] ), .B(\CARRYB[28][45] ), .CI(\SUMB[28][46] ), 
        .CO(\CARRYB[29][45] ), .S(\SUMB[29][45] ) );
  FA1 S2_38_45 ( .A(\ab[45][38] ), .B(\CARRYB[37][45] ), .CI(\SUMB[37][46] ), 
        .CO(\CARRYB[38][45] ), .S(\SUMB[38][45] ) );
  FA1P S3_38_46 ( .A(\ab[46][38] ), .B(\CARRYB[37][46] ), .CI(\ab[47][37] ), 
        .CO(\CARRYB[38][46] ), .S(\SUMB[38][46] ) );
  FA1P S2_29_33 ( .A(\ab[33][29] ), .B(\CARRYB[28][33] ), .CI(\SUMB[28][34] ), 
        .CO(\CARRYB[29][33] ), .S(\SUMB[29][33] ) );
  FA1A S2_30_32 ( .A(\ab[32][30] ), .B(\CARRYB[29][32] ), .CI(\SUMB[29][33] ), 
        .CO(\CARRYB[30][32] ), .S(\SUMB[30][32] ) );
  FA1 S2_43_5 ( .A(\CARRYB[42][5] ), .B(n446), .CI(\SUMB[42][6] ), .CO(
        \CARRYB[43][5] ), .S(\SUMB[43][5] ) );
  FA1A S2_5_43 ( .A(n446), .B(\CARRYB[4][43] ), .CI(\SUMB[4][44] ), .CO(
        \CARRYB[5][43] ), .S(\SUMB[5][43] ) );
  FA1P S2_43_30 ( .A(\CARRYB[42][30] ), .B(\ab[43][30] ), .CI(\SUMB[42][31] ), 
        .CO(\CARRYB[43][30] ), .S(\SUMB[43][30] ) );
  FA1 S2_44_30 ( .A(\ab[44][30] ), .B(\CARRYB[43][30] ), .CI(\SUMB[43][31] ), 
        .CO(\CARRYB[44][30] ), .S(\SUMB[44][30] ) );
  FA1P S2_45_31 ( .A(\ab[45][31] ), .B(\CARRYB[44][31] ), .CI(\SUMB[44][32] ), 
        .CO(\CARRYB[45][31] ), .S(\SUMB[45][31] ) );
  FA1 S2_34_33 ( .A(\ab[34][33] ), .B(\CARRYB[33][33] ), .CI(\SUMB[33][34] ), 
        .CO(\CARRYB[34][33] ), .S(\SUMB[34][33] ) );
  FA1 S2_15_19 ( .A(\CARRYB[14][19] ), .B(n725), .CI(\SUMB[14][20] ), .CO(
        \CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA1AP S2_36_25 ( .A(\ab[36][25] ), .B(\CARRYB[35][25] ), .CI(\SUMB[35][26] ), 
        .CO(\CARRYB[36][25] ), .S(\SUMB[36][25] ) );
  FA1P S2_19_32 ( .A(\ab[32][19] ), .B(\CARRYB[18][32] ), .CI(\SUMB[18][33] ), 
        .CO(\CARRYB[19][32] ), .S(\SUMB[19][32] ) );
  FA1P S2_3_37 ( .A(\CARRYB[2][37] ), .B(n342), .CI(\SUMB[2][38] ), .CO(
        \CARRYB[3][37] ), .S(\SUMB[3][37] ) );
  FA1 S2_23_34 ( .A(\CARRYB[22][34] ), .B(\ab[34][23] ), .CI(\SUMB[22][35] ), 
        .CO(\CARRYB[23][34] ), .S(\SUMB[23][34] ) );
  FA1A S2_32_31 ( .A(\ab[32][31] ), .B(\CARRYB[31][31] ), .CI(\SUMB[31][32] ), 
        .CO(\CARRYB[32][31] ), .S(\SUMB[32][31] ) );
  FA1 S2_41_35 ( .A(\ab[41][35] ), .B(\CARRYB[40][35] ), .CI(\SUMB[40][36] ), 
        .CO(\CARRYB[41][35] ), .S(\SUMB[41][35] ) );
  FA1AP S2_14_25 ( .A(\CARRYB[13][25] ), .B(n711), .CI(\SUMB[13][26] ), .CO(
        \CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA1 S2_15_25 ( .A(\SUMB[14][26] ), .B(\CARRYB[14][25] ), .CI(n723), .CO(
        \CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA1P S2_30_34 ( .A(\CARRYB[29][34] ), .B(\ab[34][30] ), .CI(\SUMB[29][35] ), 
        .CO(\CARRYB[30][34] ), .S(\SUMB[30][34] ) );
  FA1P S2_44_31 ( .A(\ab[44][31] ), .B(\CARRYB[43][31] ), .CI(\SUMB[43][32] ), 
        .CO(\CARRYB[44][31] ), .S(\SUMB[44][31] ) );
  FA1P S2_42_32 ( .A(\ab[42][32] ), .B(\CARRYB[41][32] ), .CI(\SUMB[41][33] ), 
        .CO(\CARRYB[42][32] ), .S(\SUMB[42][32] ) );
  FA1P S2_29_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA1 S2_27_27 ( .A(n2372), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), .CO(
        \CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA1P S2_7_23 ( .A(n495), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), .CO(
        \CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA1P S2_37_10 ( .A(\CARRYB[36][10] ), .B(n599), .CI(\SUMB[36][11] ), .CO(
        \CARRYB[37][10] ), .S(\SUMB[37][10] ) );
  FA1AP S2_18_32 ( .A(\CARRYB[17][32] ), .B(\ab[32][18] ), .CI(\SUMB[17][33] ), 
        .CO(\CARRYB[18][32] ), .S(\SUMB[18][32] ) );
  FA1P S2_36_26 ( .A(\CARRYB[35][26] ), .B(\ab[36][26] ), .CI(\SUMB[35][27] ), 
        .CO(\CARRYB[36][26] ), .S(\SUMB[36][26] ) );
  FA1 S2_44_23 ( .A(\ab[44][23] ), .B(\CARRYB[43][23] ), .CI(\SUMB[43][24] ), 
        .CO(\CARRYB[44][23] ), .S(\SUMB[44][23] ) );
  FA1 S2_5_36 ( .A(\CARRYB[4][36] ), .B(n399), .CI(\SUMB[4][37] ), .CO(
        \CARRYB[5][36] ), .S(\SUMB[5][36] ) );
  FA1 S2_9_42 ( .A(\CARRYB[8][42] ), .B(n583), .CI(\SUMB[8][43] ), .CO(
        \CARRYB[9][42] ), .S(\SUMB[9][42] ) );
  FA1AP S2_20_36 ( .A(\ab[36][20] ), .B(\CARRYB[19][36] ), .CI(\SUMB[19][37] ), 
        .CO(\CARRYB[20][36] ), .S(\SUMB[20][36] ) );
  FA1AP S2_32_35 ( .A(\ab[35][32] ), .B(\CARRYB[31][35] ), .CI(\SUMB[31][36] ), 
        .CO(\CARRYB[32][35] ), .S(\SUMB[32][35] ) );
  FA1P S2_44_32 ( .A(\ab[44][32] ), .B(\CARRYB[43][32] ), .CI(\SUMB[43][33] ), 
        .CO(\CARRYB[44][32] ), .S(\SUMB[44][32] ) );
  FA1P S2_33_19 ( .A(\CARRYB[32][19] ), .B(\ab[33][19] ), .CI(\SUMB[32][20] ), 
        .CO(\CARRYB[33][19] ), .S(\SUMB[33][19] ) );
  FA1A S2_34_19 ( .A(\CARRYB[33][19] ), .B(\ab[34][19] ), .CI(\SUMB[33][20] ), 
        .CO(\CARRYB[34][19] ), .S(\SUMB[34][19] ) );
  FA1AP S2_16_18 ( .A(\CARRYB[15][18] ), .B(\ab[18][16] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA1AP S2_38_10 ( .A(\CARRYB[37][10] ), .B(n613), .CI(\SUMB[37][11] ), .CO(
        \CARRYB[38][10] ), .S(\SUMB[38][10] ) );
  FA1A S2_28_33 ( .A(\ab[33][28] ), .B(\CARRYB[27][33] ), .CI(\SUMB[27][34] ), 
        .CO(\CARRYB[28][33] ), .S(\SUMB[28][33] ) );
  FA1 S2_31_32 ( .A(\ab[32][31] ), .B(\CARRYB[30][32] ), .CI(\SUMB[30][33] ), 
        .CO(\CARRYB[31][32] ), .S(\SUMB[31][32] ) );
  FA1AP S2_20_13 ( .A(n688), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), .CO(
        \CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA1AP S2_28_10 ( .A(\CARRYB[27][10] ), .B(n610), .CI(\SUMB[27][11] ), .CO(
        \CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA1AP S2_15_20 ( .A(n724), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), .CO(
        \CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA1P S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA1AP S2_5_24 ( .A(\CARRYB[4][24] ), .B(n421), .CI(\SUMB[4][25] ), .CO(
        \CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1P S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), 
        .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FA1 S2_24_21 ( .A(\CARRYB[23][21] ), .B(\ab[24][21] ), .CI(\SUMB[23][22] ), 
        .CO(\CARRYB[24][21] ), .S(\SUMB[24][21] ) );
  FA1AP S2_28_20 ( .A(\CARRYB[27][20] ), .B(\ab[28][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA1P S2_41_33 ( .A(\ab[41][33] ), .B(\CARRYB[40][33] ), .CI(\SUMB[40][34] ), 
        .CO(\CARRYB[41][33] ), .S(\SUMB[41][33] ) );
  FA1P S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), 
        .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FA1P S2_35_18 ( .A(\CARRYB[34][18] ), .B(\ab[35][18] ), .CI(\SUMB[34][19] ), 
        .CO(\CARRYB[35][18] ), .S(\SUMB[35][18] ) );
  FA1P S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA1AP S2_29_31 ( .A(\ab[31][29] ), .B(\CARRYB[28][31] ), .CI(\SUMB[28][32] ), 
        .CO(\CARRYB[29][31] ), .S(\SUMB[29][31] ) );
  FA1P S2_9_21 ( .A(\CARRYB[8][21] ), .B(n561), .CI(\SUMB[8][22] ), .CO(
        \CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA1P S2_38_36 ( .A(\ab[38][36] ), .B(\CARRYB[37][36] ), .CI(\SUMB[37][37] ), 
        .CO(\CARRYB[38][36] ), .S(\SUMB[38][36] ) );
  FA1P S2_43_36 ( .A(\ab[43][36] ), .B(\CARRYB[42][36] ), .CI(\SUMB[42][37] ), 
        .CO(\CARRYB[43][36] ), .S(\SUMB[43][36] ) );
  FA1AP S2_29_37 ( .A(\ab[37][29] ), .B(\CARRYB[28][37] ), .CI(\SUMB[28][38] ), 
        .CO(\CARRYB[29][37] ), .S(\SUMB[29][37] ) );
  FA1P S2_35_35 ( .A(n300), .B(\CARRYB[34][35] ), .CI(\SUMB[34][36] ), .CO(
        \CARRYB[35][35] ), .S(\SUMB[35][35] ) );
  FA1 S2_32_36 ( .A(\ab[36][32] ), .B(\CARRYB[31][36] ), .CI(\SUMB[31][37] ), 
        .CO(\CARRYB[32][36] ), .S(\SUMB[32][36] ) );
  FA1 S2_8_42 ( .A(n550), .B(\CARRYB[7][42] ), .CI(\SUMB[7][43] ), .CO(
        \CARRYB[8][42] ), .S(\SUMB[8][42] ) );
  FA1 S2_14_39 ( .A(\ab[39][14] ), .B(\CARRYB[13][39] ), .CI(\SUMB[13][40] ), 
        .CO(\CARRYB[14][39] ), .S(\SUMB[14][39] ) );
  FA1AP S4_26 ( .A(\ab[47][26] ), .B(\CARRYB[46][26] ), .CI(\SUMB[46][27] ), 
        .CO(\CARRYB[47][26] ), .S(\SUMB[47][26] ) );
  FA1P S2_37_40 ( .A(\ab[40][37] ), .B(\CARRYB[36][40] ), .CI(\SUMB[36][41] ), 
        .CO(\CARRYB[37][40] ), .S(\SUMB[37][40] ) );
  FA1P S2_42_40 ( .A(\ab[42][40] ), .B(\CARRYB[41][40] ), .CI(\SUMB[41][41] ), 
        .CO(\CARRYB[42][40] ), .S(\SUMB[42][40] ) );
  FA1P S2_11_22 ( .A(\CARRYB[10][22] ), .B(n641), .CI(\SUMB[10][23] ), .CO(
        \CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1AP S2_44_11 ( .A(\ab[44][11] ), .B(\CARRYB[43][11] ), .CI(\SUMB[43][12] ), 
        .CO(\CARRYB[44][11] ), .S(\SUMB[44][11] ) );
  FA1P S2_45_10 ( .A(\SUMB[44][11] ), .B(\CARRYB[44][10] ), .CI(\ab[45][10] ), 
        .CO(\CARRYB[45][10] ), .S(\SUMB[45][10] ) );
  FA1P S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA1AP S2_18_37 ( .A(\ab[37][18] ), .B(\CARRYB[17][37] ), .CI(\SUMB[17][38] ), 
        .CO(\CARRYB[18][37] ), .S(\SUMB[18][37] ) );
  FA1P S2_16_22 ( .A(\CARRYB[15][22] ), .B(\ab[22][16] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA1A S2_17_22 ( .A(\CARRYB[16][22] ), .B(\ab[22][17] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA1 S2_12_23 ( .A(\CARRYB[11][23] ), .B(n666), .CI(\SUMB[11][24] ), .CO(
        \CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA1P S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA1AP S2_39_7 ( .A(n511), .B(\CARRYB[38][7] ), .CI(\SUMB[38][8] ), .CO(
        \CARRYB[39][7] ), .S(\SUMB[39][7] ) );
  FA1A S2_35_9 ( .A(n307), .B(\CARRYB[34][9] ), .CI(\SUMB[34][10] ), .CO(
        \CARRYB[35][9] ), .S(\SUMB[35][9] ) );
  FA1 S2_38_9 ( .A(n589), .B(\CARRYB[37][9] ), .CI(\SUMB[37][10] ), .CO(
        \CARRYB[38][9] ), .S(\SUMB[38][9] ) );
  FA1P S2_28_29 ( .A(\ab[29][28] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA1 S4_22 ( .A(\ab[47][22] ), .B(\CARRYB[46][22] ), .CI(\SUMB[46][23] ), 
        .CO(\CARRYB[47][22] ), .S(\SUMB[47][22] ) );
  FA1AP S2_30_9 ( .A(n592), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), .CO(
        \CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA1P S2_34_8 ( .A(n522), .B(\CARRYB[33][8] ), .CI(\SUMB[33][9] ), .CO(
        \CARRYB[34][8] ), .S(\SUMB[34][8] ) );
  FA1 S2_31_8 ( .A(\CARRYB[30][8] ), .B(n514), .CI(\SUMB[30][9] ), .CO(
        \CARRYB[31][8] ), .S(\SUMB[31][8] ) );
  FA1AP S2_40_4 ( .A(\CARRYB[39][4] ), .B(n414), .CI(\SUMB[39][5] ), .CO(
        \CARRYB[40][4] ), .S(\SUMB[40][4] ) );
  FA1P S2_32_9 ( .A(n568), .B(\CARRYB[31][9] ), .CI(\SUMB[31][10] ), .CO(
        \CARRYB[32][9] ), .S(\SUMB[32][9] ) );
  FA1A S2_14_19 ( .A(\CARRYB[13][19] ), .B(n699), .CI(\SUMB[13][20] ), .CO(
        \CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA1P S2_14_16 ( .A(\CARRYB[13][16] ), .B(n701), .CI(\SUMB[13][17] ), .CO(
        \CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA1P S2_17_15 ( .A(\CARRYB[16][15] ), .B(n717), .CI(\SUMB[16][16] ), .CO(
        \CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA1P S2_17_41 ( .A(\ab[41][17] ), .B(\CARRYB[16][41] ), .CI(\SUMB[16][42] ), 
        .CO(\CARRYB[17][41] ), .S(\SUMB[17][41] ) );
  FA1AP S2_25_37 ( .A(\ab[37][25] ), .B(\CARRYB[24][37] ), .CI(\SUMB[24][38] ), 
        .CO(\CARRYB[25][37] ), .S(\SUMB[25][37] ) );
  FA1AP S2_27_36 ( .A(\ab[36][27] ), .B(\CARRYB[26][36] ), .CI(\SUMB[26][37] ), 
        .CO(\CARRYB[27][36] ), .S(\SUMB[27][36] ) );
  FA1P S2_39_23 ( .A(\ab[39][23] ), .B(\CARRYB[38][23] ), .CI(\SUMB[38][24] ), 
        .CO(\CARRYB[39][23] ), .S(\SUMB[39][23] ) );
  FA1P S2_27_29 ( .A(\ab[29][27] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA1P S2_5_5 ( .A(n2331), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1P S2_11_4 ( .A(n388), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(
        \CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1 S2_33_2 ( .A(n2212), .B(\CARRYB[32][2] ), .CI(\SUMB[32][3] ), .CO(
        \CARRYB[33][2] ), .S(\SUMB[33][2] ) );
  FA1P S2_25_3 ( .A(n2269), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), .CO(
        \CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA1P S2_34_2 ( .A(n2213), .B(\CARRYB[33][2] ), .CI(\SUMB[33][3] ), .CO(
        \CARRYB[34][2] ), .S(\SUMB[34][2] ) );
  FA1 S2_24_44 ( .A(\ab[44][24] ), .B(\CARRYB[23][44] ), .CI(\SUMB[23][45] ), 
        .CO(\CARRYB[24][44] ), .S(\SUMB[24][44] ) );
  FA1 S2_40_42 ( .A(\ab[42][40] ), .B(\CARRYB[39][42] ), .CI(\SUMB[39][43] ), 
        .CO(\CARRYB[40][42] ), .S(\SUMB[40][42] ) );
  FA1P S2_38_43 ( .A(\ab[43][38] ), .B(\CARRYB[37][43] ), .CI(\SUMB[37][44] ), 
        .CO(\CARRYB[38][43] ), .S(\SUMB[38][43] ) );
  FA1P S4_41 ( .A(\ab[47][41] ), .B(\CARRYB[46][41] ), .CI(\SUMB[46][42] ), 
        .CO(\CARRYB[47][41] ), .S(\SUMB[47][41] ) );
  FA1A S2_19_45 ( .A(\ab[45][19] ), .B(\CARRYB[18][45] ), .CI(\SUMB[18][46] ), 
        .CO(\CARRYB[19][45] ), .S(\SUMB[19][45] ) );
  FA1A S2_22_45 ( .A(\ab[45][22] ), .B(\CARRYB[21][45] ), .CI(\SUMB[21][46] ), 
        .CO(\CARRYB[22][45] ), .S(\SUMB[22][45] ) );
  FA1 S2_25_30 ( .A(\ab[30][25] ), .B(\CARRYB[24][30] ), .CI(\SUMB[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA1 S2_36_28 ( .A(\ab[36][28] ), .B(\CARRYB[35][28] ), .CI(\SUMB[35][29] ), 
        .CO(\CARRYB[36][28] ), .S(\SUMB[36][28] ) );
  FA1 S2_22_22 ( .A(n2364), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), .CO(
        \CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA1P S2_23_22 ( .A(\CARRYB[22][22] ), .B(\ab[23][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA1P S2_36_24 ( .A(\ab[36][24] ), .B(\CARRYB[35][24] ), .CI(\SUMB[35][25] ), 
        .CO(\CARRYB[36][24] ), .S(\SUMB[36][24] ) );
  FA1A S2_2_37 ( .A(\CARRYB[1][37] ), .B(n318), .CI(\SUMB[1][38] ), .CO(
        \CARRYB[2][37] ), .S(\SUMB[2][37] ) );
  FA1 S2_25_13 ( .A(\CARRYB[24][13] ), .B(n683), .CI(\SUMB[24][14] ), .CO(
        \CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA1 S2_10_21 ( .A(n616), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), .CO(
        \CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1P S2_26_13 ( .A(\CARRYB[25][13] ), .B(n680), .CI(\SUMB[25][14] ), .CO(
        \CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA1AP S2_22_35 ( .A(\ab[35][22] ), .B(\CARRYB[21][35] ), .CI(\SUMB[21][36] ), 
        .CO(\CARRYB[22][35] ), .S(\SUMB[22][35] ) );
  FA1P S2_6_24 ( .A(n462), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), .CO(
        \CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1P S2_37_14 ( .A(\CARRYB[36][14] ), .B(\ab[37][14] ), .CI(\SUMB[36][15] ), 
        .CO(\CARRYB[37][14] ), .S(\SUMB[37][14] ) );
  FA1 S2_8_11 ( .A(n542), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), .CO(
        \CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1AP S2_9_11 ( .A(n594), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), .CO(
        \CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1 S2_30_6 ( .A(n431), .B(\CARRYB[29][6] ), .CI(\SUMB[29][7] ), .CO(
        \CARRYB[30][6] ), .S(\SUMB[30][6] ) );
  FA1P S2_31_6 ( .A(n465), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), .CO(
        \CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FA1 S2_35_6 ( .A(\CARRYB[34][6] ), .B(n409), .CI(\SUMB[34][7] ), .CO(
        \CARRYB[35][6] ), .S(\SUMB[35][6] ) );
  FA1AP S2_36_6 ( .A(\CARRYB[35][6] ), .B(n443), .CI(\SUMB[35][7] ), .CO(
        \CARRYB[36][6] ), .S(\SUMB[36][6] ) );
  FA1P S2_6_12 ( .A(n466), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), .CO(
        \CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1P S2_12_11 ( .A(n644), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), .CO(
        \CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1 S2_22_9 ( .A(n565), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), .CO(
        \CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA1P S2_18_16 ( .A(\CARRYB[17][16] ), .B(\ab[18][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA1P S2_9_38 ( .A(n589), .B(\CARRYB[8][38] ), .CI(\SUMB[8][39] ), .CO(
        \CARRYB[9][38] ), .S(\SUMB[9][38] ) );
  FA1P S2_7_39 ( .A(n511), .B(\CARRYB[6][39] ), .CI(\SUMB[6][40] ), .CO(
        \CARRYB[7][39] ), .S(\SUMB[7][39] ) );
  FA1AP S2_7_38 ( .A(n490), .B(\CARRYB[6][38] ), .CI(\SUMB[6][39] ), .CO(
        \CARRYB[7][38] ), .S(\SUMB[7][38] ) );
  FA1P S2_37_31 ( .A(\ab[37][31] ), .B(\CARRYB[36][31] ), .CI(\SUMB[36][32] ), 
        .CO(\CARRYB[37][31] ), .S(\SUMB[37][31] ) );
  FA1A S2_38_30 ( .A(\CARRYB[37][30] ), .B(\ab[38][30] ), .CI(\SUMB[37][31] ), 
        .CO(\CARRYB[38][30] ), .S(\SUMB[38][30] ) );
  FA1AP S2_34_13 ( .A(\ab[34][13] ), .B(\CARRYB[33][13] ), .CI(\SUMB[33][14] ), 
        .CO(\CARRYB[34][13] ), .S(\SUMB[34][13] ) );
  FA1AP S2_38_24 ( .A(\CARRYB[37][24] ), .B(\ab[38][24] ), .CI(\SUMB[37][25] ), 
        .CO(\CARRYB[38][24] ), .S(\SUMB[38][24] ) );
  FA1P S2_3_38 ( .A(\CARRYB[2][38] ), .B(n2294), .CI(\SUMB[2][39] ), .CO(
        \CARRYB[3][38] ), .S(\SUMB[3][38] ) );
  FA1P S2_9_35 ( .A(\CARRYB[8][35] ), .B(n307), .CI(\SUMB[8][36] ), .CO(
        \CARRYB[9][35] ), .S(\SUMB[9][35] ) );
  FA1A S2_31_26 ( .A(\ab[31][26] ), .B(\CARRYB[30][26] ), .CI(\SUMB[30][27] ), 
        .CO(\CARRYB[31][26] ), .S(\SUMB[31][26] ) );
  FA1AP S2_9_43 ( .A(n586), .B(\CARRYB[8][43] ), .CI(\SUMB[8][44] ), .CO(
        \CARRYB[9][43] ), .S(\SUMB[9][43] ) );
  FA1P S2_42_33 ( .A(\ab[42][33] ), .B(\CARRYB[41][33] ), .CI(\SUMB[41][34] ), 
        .CO(\CARRYB[42][33] ), .S(\SUMB[42][33] ) );
  FA1 S2_17_40 ( .A(\ab[40][17] ), .B(\CARRYB[16][40] ), .CI(\SUMB[16][41] ), 
        .CO(\CARRYB[17][40] ), .S(\SUMB[17][40] ) );
  FA1P S2_18_40 ( .A(\ab[40][18] ), .B(\CARRYB[17][40] ), .CI(\SUMB[17][41] ), 
        .CO(\CARRYB[18][40] ), .S(\SUMB[18][40] ) );
  FA1 S2_28_38 ( .A(\ab[38][28] ), .B(\CARRYB[27][38] ), .CI(\SUMB[27][39] ), 
        .CO(\CARRYB[28][38] ), .S(\SUMB[28][38] ) );
  FA1AP S2_3_25 ( .A(n2269), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), .CO(
        \CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA1 S2_30_11 ( .A(\CARRYB[29][11] ), .B(n623), .CI(\SUMB[29][12] ), .CO(
        \CARRYB[30][11] ), .S(\SUMB[30][11] ) );
  FA1P S2_34_9 ( .A(\CARRYB[33][9] ), .B(n555), .CI(\SUMB[33][10] ), .CO(
        \CARRYB[34][9] ), .S(\SUMB[34][9] ) );
  FA1 S2_17_18 ( .A(\ab[18][17] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA1AP S2_18_18 ( .A(\CARRYB[17][18] ), .B(n2356), .CI(\SUMB[17][19] ), .CO(
        \CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA1AP S2_44_28 ( .A(\ab[44][28] ), .B(\CARRYB[43][28] ), .CI(\SUMB[43][29] ), 
        .CO(\CARRYB[44][28] ), .S(\SUMB[44][28] ) );
  FA1A S2_25_32 ( .A(\ab[32][25] ), .B(\CARRYB[24][32] ), .CI(\SUMB[24][33] ), 
        .CO(\CARRYB[25][32] ), .S(\SUMB[25][32] ) );
  FA1AP S4_27 ( .A(\CARRYB[46][27] ), .B(\ab[47][27] ), .CI(\SUMB[46][28] ), 
        .CO(\CARRYB[47][27] ), .S(\SUMB[47][27] ) );
  FA1P S2_15_42 ( .A(\ab[42][15] ), .B(\CARRYB[14][42] ), .CI(\SUMB[14][43] ), 
        .CO(\CARRYB[15][42] ), .S(\SUMB[15][42] ) );
  FA1P S2_38_39 ( .A(\ab[39][38] ), .B(\CARRYB[37][39] ), .CI(\SUMB[37][40] ), 
        .CO(\CARRYB[38][39] ), .S(\SUMB[38][39] ) );
  FA1A S2_32_41 ( .A(\ab[41][32] ), .B(\CARRYB[31][41] ), .CI(\SUMB[31][42] ), 
        .CO(\CARRYB[32][41] ), .S(\SUMB[32][41] ) );
  FA1P S2_42_39 ( .A(\ab[42][39] ), .B(\CARRYB[41][39] ), .CI(\SUMB[41][40] ), 
        .CO(\CARRYB[42][39] ), .S(\SUMB[42][39] ) );
  FA1P S2_13_43 ( .A(\ab[43][13] ), .B(\CARRYB[12][43] ), .CI(\SUMB[12][44] ), 
        .CO(\CARRYB[13][43] ), .S(\SUMB[13][43] ) );
  FA1 S2_6_34 ( .A(n459), .B(\CARRYB[5][34] ), .CI(\SUMB[5][35] ), .CO(
        \CARRYB[6][34] ), .S(\SUMB[6][34] ) );
  FA1P S2_16_28 ( .A(\ab[28][16] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA1 S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA1P S2_38_15 ( .A(\CARRYB[37][15] ), .B(\ab[38][15] ), .CI(\SUMB[37][16] ), 
        .CO(\CARRYB[38][15] ), .S(\SUMB[38][15] ) );
  FA1AP S2_33_16 ( .A(\ab[33][16] ), .B(\CARRYB[32][16] ), .CI(\SUMB[32][17] ), 
        .CO(\CARRYB[33][16] ), .S(\SUMB[33][16] ) );
  FA1P S2_11_32 ( .A(n622), .B(\CARRYB[10][32] ), .CI(\SUMB[10][33] ), .CO(
        \CARRYB[11][32] ), .S(\SUMB[11][32] ) );
  FA1 S2_12_20 ( .A(\CARRYB[11][20] ), .B(n665), .CI(\SUMB[11][21] ), .CO(
        \CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA1P S2_29_11 ( .A(\CARRYB[28][11] ), .B(n639), .CI(\SUMB[28][12] ), .CO(
        \CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA1 S2_41_22 ( .A(\ab[41][22] ), .B(\CARRYB[40][22] ), .CI(\SUMB[40][23] ), 
        .CO(\CARRYB[41][22] ), .S(\SUMB[41][22] ) );
  FA1AP S2_42_22 ( .A(\ab[42][22] ), .B(\CARRYB[41][22] ), .CI(\SUMB[41][23] ), 
        .CO(\CARRYB[42][22] ), .S(\SUMB[42][22] ) );
  FA1P S2_24_30 ( .A(\ab[30][24] ), .B(\CARRYB[23][30] ), .CI(\SUMB[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA1AP S2_19_29 ( .A(\CARRYB[18][29] ), .B(\ab[29][19] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA1AP S2_21_28 ( .A(\CARRYB[20][28] ), .B(\ab[28][21] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA1A S2_37_16 ( .A(\CARRYB[36][16] ), .B(\ab[37][16] ), .CI(\SUMB[36][17] ), 
        .CO(\CARRYB[37][16] ), .S(\SUMB[37][16] ) );
  FA1A S2_9_28 ( .A(n563), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), .CO(
        \CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1AP S2_25_26 ( .A(\CARRYB[24][26] ), .B(\ab[26][25] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA1AP S2_2_39 ( .A(\CARRYB[1][39] ), .B(n2261), .CI(\SUMB[1][40] ), .CO(
        \CARRYB[2][39] ), .S(\SUMB[2][39] ) );
  FA1P S2_45_25 ( .A(\CARRYB[44][25] ), .B(\ab[45][25] ), .CI(\SUMB[44][26] ), 
        .CO(\CARRYB[45][25] ), .S(\SUMB[45][25] ) );
  FA1A S2_14_20 ( .A(n709), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), .CO(
        \CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA1A S2_16_19 ( .A(\ab[19][16] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA1AP S2_14_31 ( .A(\CARRYB[13][31] ), .B(\ab[31][14] ), .CI(\SUMB[13][32] ), 
        .CO(\CARRYB[14][31] ), .S(\SUMB[14][31] ) );
  FA1 S2_24_34 ( .A(\ab[34][24] ), .B(\CARRYB[23][34] ), .CI(\SUMB[23][35] ), 
        .CO(\CARRYB[24][34] ), .S(\SUMB[24][34] ) );
  FA1 S2_13_23 ( .A(\CARRYB[12][23] ), .B(n684), .CI(\SUMB[12][24] ), .CO(
        \CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA1AP S2_21_32 ( .A(\CARRYB[20][32] ), .B(\ab[32][21] ), .CI(\SUMB[20][33] ), 
        .CO(\CARRYB[21][32] ), .S(\SUMB[21][32] ) );
  FA1P S2_17_35 ( .A(\ab[35][17] ), .B(\CARRYB[16][35] ), .CI(\SUMB[16][36] ), 
        .CO(\CARRYB[17][35] ), .S(\SUMB[17][35] ) );
  FA1P S2_29_29 ( .A(n2378), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), .CO(
        \CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA1A S2_45_23 ( .A(\ab[45][23] ), .B(\CARRYB[44][23] ), .CI(\SUMB[44][24] ), 
        .CO(\CARRYB[45][23] ), .S(\SUMB[45][23] ) );
  FA1 S2_32_14 ( .A(\CARRYB[31][14] ), .B(\ab[32][14] ), .CI(\SUMB[31][15] ), 
        .CO(\CARRYB[32][14] ), .S(\SUMB[32][14] ) );
  FA1A S2_46_6 ( .A(n457), .B(\CARRYB[45][6] ), .CI(\SUMB[45][7] ), .CO(
        \CARRYB[46][6] ), .S(\SUMB[46][6] ) );
  FA1AP S2_40_23 ( .A(\ab[40][23] ), .B(\CARRYB[39][23] ), .CI(\SUMB[39][24] ), 
        .CO(\CARRYB[40][23] ), .S(\SUMB[40][23] ) );
  FA1AP S2_45_21 ( .A(\CARRYB[44][21] ), .B(\ab[45][21] ), .CI(\SUMB[44][22] ), 
        .CO(\CARRYB[45][21] ), .S(\SUMB[45][21] ) );
  FA1AP S2_34_26 ( .A(\CARRYB[33][26] ), .B(\ab[34][26] ), .CI(\SUMB[33][27] ), 
        .CO(\CARRYB[34][26] ), .S(\SUMB[34][26] ) );
  FA1AP S2_7_30 ( .A(\CARRYB[6][30] ), .B(n489), .CI(\SUMB[6][31] ), .CO(
        \CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA1P S2_8_30 ( .A(\CARRYB[7][30] ), .B(n541), .CI(\SUMB[7][31] ), .CO(
        \CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA1 S2_39_19 ( .A(\ab[39][19] ), .B(\CARRYB[38][19] ), .CI(\SUMB[38][20] ), 
        .CO(\CARRYB[39][19] ), .S(\SUMB[39][19] ) );
  FA1A S2_40_18 ( .A(\ab[40][18] ), .B(\CARRYB[39][18] ), .CI(\SUMB[39][19] ), 
        .CO(\CARRYB[40][18] ), .S(\SUMB[40][18] ) );
  FA1A S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA1A S2_24_24 ( .A(n2368), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), .CO(
        \CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA1 S2_41_18 ( .A(\CARRYB[40][18] ), .B(\ab[41][18] ), .CI(\SUMB[40][19] ), 
        .CO(\CARRYB[41][18] ), .S(\SUMB[41][18] ) );
  FA1A S2_44_27 ( .A(\ab[44][27] ), .B(\CARRYB[43][27] ), .CI(\SUMB[43][28] ), 
        .CO(\CARRYB[44][27] ), .S(\SUMB[44][27] ) );
  FA1AP S2_37_39 ( .A(\ab[39][37] ), .B(\CARRYB[36][39] ), .CI(\SUMB[36][40] ), 
        .CO(\CARRYB[37][39] ), .S(\SUMB[37][39] ) );
  FA1P S2_26_43 ( .A(\ab[43][26] ), .B(\CARRYB[25][43] ), .CI(\SUMB[25][44] ), 
        .CO(\CARRYB[26][43] ), .S(\SUMB[26][43] ) );
  FA1A S2_46_35 ( .A(\ab[46][35] ), .B(\CARRYB[45][35] ), .CI(\SUMB[45][36] ), 
        .CO(\CARRYB[46][35] ), .S(\SUMB[46][35] ) );
  FA1P S2_36_29 ( .A(\ab[36][29] ), .B(\CARRYB[35][29] ), .CI(\SUMB[35][30] ), 
        .CO(\CARRYB[36][29] ), .S(\SUMB[36][29] ) );
  FA1A S2_27_32 ( .A(\ab[32][27] ), .B(\CARRYB[26][32] ), .CI(\SUMB[26][33] ), 
        .CO(\CARRYB[27][32] ), .S(\SUMB[27][32] ) );
  FA1A S2_38_28 ( .A(\ab[38][28] ), .B(\CARRYB[37][28] ), .CI(\SUMB[37][29] ), 
        .CO(\CARRYB[38][28] ), .S(\SUMB[38][28] ) );
  FA1AP S2_13_14 ( .A(n675), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), .CO(
        \CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1 S2_25_9 ( .A(\CARRYB[24][9] ), .B(n557), .CI(\SUMB[24][10] ), .CO(
        \CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA1P S2_38_6 ( .A(n456), .B(\CARRYB[37][6] ), .CI(\SUMB[37][7] ), .CO(
        \CARRYB[38][6] ), .S(\SUMB[38][6] ) );
  FA1A S2_25_19 ( .A(\CARRYB[24][19] ), .B(\ab[25][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA1P S2_6_35 ( .A(\CARRYB[5][35] ), .B(n409), .CI(\SUMB[5][36] ), .CO(
        \CARRYB[6][35] ), .S(\SUMB[6][35] ) );
  FA1P S2_42_13 ( .A(\CARRYB[41][13] ), .B(\ab[42][13] ), .CI(\SUMB[41][14] ), 
        .CO(\CARRYB[42][13] ), .S(\SUMB[42][13] ) );
  FA1 S2_43_13 ( .A(\CARRYB[42][13] ), .B(\ab[43][13] ), .CI(\SUMB[42][14] ), 
        .CO(\CARRYB[43][13] ), .S(\SUMB[43][13] ) );
  FA1 S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA1 S2_12_27 ( .A(n663), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), .CO(
        \CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA1 S2_38_16 ( .A(\CARRYB[37][16] ), .B(\ab[38][16] ), .CI(\SUMB[37][17] ), 
        .CO(\CARRYB[38][16] ), .S(\SUMB[38][16] ) );
  FA1 S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA1 S2_15_27 ( .A(\CARRYB[14][27] ), .B(n718), .CI(\SUMB[14][28] ), .CO(
        \CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA1 S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA1P S2_26_19 ( .A(\CARRYB[25][19] ), .B(\ab[26][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA1AP S2_15_29 ( .A(n714), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), .CO(
        \CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA1AP S2_39_15 ( .A(\ab[39][15] ), .B(\CARRYB[38][15] ), .CI(\SUMB[38][16] ), 
        .CO(\CARRYB[39][15] ), .S(\SUMB[39][15] ) );
  FA1P S2_12_31 ( .A(\SUMB[11][32] ), .B(\CARRYB[11][31] ), .CI(n673), .CO(
        \CARRYB[12][31] ), .S(\SUMB[12][31] ) );
  FA1 S2_36_22 ( .A(\ab[36][22] ), .B(\CARRYB[35][22] ), .CI(\SUMB[35][23] ), 
        .CO(\CARRYB[36][22] ), .S(\SUMB[36][22] ) );
  FA1AP S2_21_38 ( .A(\ab[38][21] ), .B(\CARRYB[20][38] ), .CI(\SUMB[20][39] ), 
        .CO(\CARRYB[21][38] ), .S(\SUMB[21][38] ) );
  FA1 S2_37_32 ( .A(\CARRYB[36][32] ), .B(\ab[37][32] ), .CI(\SUMB[36][33] ), 
        .CO(\CARRYB[37][32] ), .S(\SUMB[37][32] ) );
  FA1AP S2_33_34 ( .A(\CARRYB[32][34] ), .B(\ab[34][33] ), .CI(\SUMB[32][35] ), 
        .CO(\CARRYB[33][34] ), .S(\SUMB[33][34] ) );
  FA1A S2_44_29 ( .A(\ab[44][29] ), .B(\CARRYB[43][29] ), .CI(\SUMB[43][30] ), 
        .CO(\CARRYB[44][29] ), .S(\SUMB[44][29] ) );
  FA1AP S2_45_29 ( .A(\ab[45][29] ), .B(\CARRYB[44][29] ), .CI(\SUMB[44][30] ), 
        .CO(\CARRYB[45][29] ), .S(\SUMB[45][29] ) );
  FA1P S1_13_0 ( .A(n2191), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), .CO(
        \CARRYB[13][0] ), .S(\A1[11] ) );
  FA1 S2_23_21 ( .A(\CARRYB[22][21] ), .B(\ab[23][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA1 S2_36_16 ( .A(\ab[36][16] ), .B(\CARRYB[35][16] ), .CI(\SUMB[35][17] ), 
        .CO(\CARRYB[36][16] ), .S(\SUMB[36][16] ) );
  FA1A S2_9_18 ( .A(n560), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), .CO(
        \CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1AP S2_33_23 ( .A(\ab[33][23] ), .B(\CARRYB[32][23] ), .CI(\SUMB[32][24] ), 
        .CO(\CARRYB[33][23] ), .S(\SUMB[33][23] ) );
  FA1P S2_3_34 ( .A(n2276), .B(\CARRYB[2][34] ), .CI(\SUMB[2][35] ), .CO(
        \CARRYB[3][34] ), .S(\SUMB[3][34] ) );
  FA1AP S2_8_23 ( .A(\CARRYB[7][23] ), .B(n533), .CI(\SUMB[7][24] ), .CO(
        \CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1P S2_13_21 ( .A(\CARRYB[12][21] ), .B(n696), .CI(\SUMB[12][22] ), .CO(
        \CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA1A S2_17_19 ( .A(\ab[19][17] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA1 S2_43_8 ( .A(n520), .B(\CARRYB[42][8] ), .CI(\SUMB[42][9] ), .CO(
        \CARRYB[43][8] ), .S(\SUMB[43][8] ) );
  AN2P U2 ( .A(n1350), .B(n2427), .Z(\CARRYB[1][1] ) );
  EOP U3 ( .A(n2427), .B(n1350), .Z(\SUMB[1][1] ) );
  ND3P U4 ( .A(n839), .B(n840), .C(n841), .Z(\CARRYB[38][22] ) );
  ND3P U5 ( .A(n994), .B(n995), .C(n996), .Z(\CARRYB[3][21] ) );
  ND2P U6 ( .A(\CARRYB[11][25] ), .B(n661), .Z(n1168) );
  ND2P U7 ( .A(\CARRYB[11][25] ), .B(\SUMB[11][26] ), .Z(n1167) );
  EO3 U8 ( .A(\CARRYB[39][14] ), .B(\ab[40][14] ), .C(\SUMB[39][15] ), .Z(
        \SUMB[40][14] ) );
  ND2 U9 ( .A(\CARRYB[39][14] ), .B(\SUMB[39][15] ), .Z(n3) );
  ND2 U10 ( .A(\CARRYB[39][14] ), .B(\ab[40][14] ), .Z(n4) );
  ND2 U11 ( .A(\SUMB[39][15] ), .B(\ab[40][14] ), .Z(n5) );
  ND3 U12 ( .A(n3), .B(n4), .C(n5), .Z(\CARRYB[40][14] ) );
  EOP U13 ( .A(\SUMB[35][20] ), .B(n1143), .Z(\SUMB[36][19] ) );
  ND3P U14 ( .A(n1905), .B(n1906), .C(n1907), .Z(\CARRYB[43][15] ) );
  EOP U15 ( .A(\CARRYB[19][26] ), .B(n1147), .Z(\SUMB[20][26] ) );
  EO U16 ( .A(\SUMB[19][27] ), .B(\ab[26][20] ), .Z(n1147) );
  EO U17 ( .A(\SUMB[27][33] ), .B(\ab[32][28] ), .Z(n6) );
  EO U18 ( .A(\CARRYB[27][32] ), .B(n6), .Z(\SUMB[28][32] ) );
  ND2 U19 ( .A(\CARRYB[27][32] ), .B(\SUMB[27][33] ), .Z(n7) );
  ND2 U20 ( .A(\CARRYB[27][32] ), .B(\ab[32][28] ), .Z(n8) );
  ND2 U21 ( .A(\SUMB[27][33] ), .B(\ab[32][28] ), .Z(n9) );
  ND3 U22 ( .A(n7), .B(n8), .C(n9), .Z(\CARRYB[28][32] ) );
  EOP U23 ( .A(\CARRYB[40][13] ), .B(\ab[41][13] ), .Z(n1234) );
  ND3P U24 ( .A(n1235), .B(n1236), .C(n1237), .Z(\CARRYB[41][13] ) );
  ND3 U25 ( .A(n1151), .B(n1152), .C(n1153), .Z(n10) );
  EO U26 ( .A(\CARRYB[36][20] ), .B(\ab[37][20] ), .Z(n11) );
  EO U27 ( .A(\SUMB[36][21] ), .B(n11), .Z(\SUMB[37][20] ) );
  ND2 U28 ( .A(\SUMB[36][21] ), .B(\CARRYB[36][20] ), .Z(n12) );
  ND2 U29 ( .A(\SUMB[36][21] ), .B(\ab[37][20] ), .Z(n13) );
  ND2 U30 ( .A(\CARRYB[36][20] ), .B(\ab[37][20] ), .Z(n14) );
  ND3 U31 ( .A(n12), .B(n13), .C(n14), .Z(\CARRYB[37][20] ) );
  IVDA U32 ( .A(n2175), .Z(n15) );
  ND3 U33 ( .A(n1151), .B(n1152), .C(n1153), .Z(\CARRYB[13][32] ) );
  ND3 U34 ( .A(n1206), .B(n1207), .C(n1208), .Z(\CARRYB[43][27] ) );
  ND2P U35 ( .A(\CARRYB[35][19] ), .B(\ab[36][19] ), .Z(n1146) );
  ND2P U36 ( .A(A[38]), .B(n2040), .Z(n1731) );
  EOP U37 ( .A(\SUMB[44][7] ), .B(n485), .Z(n16) );
  EO U38 ( .A(\CARRYB[44][6] ), .B(n16), .Z(\SUMB[45][6] ) );
  ND2 U39 ( .A(\CARRYB[44][6] ), .B(\SUMB[44][7] ), .Z(n17) );
  ND2 U40 ( .A(\CARRYB[44][6] ), .B(n485), .Z(n18) );
  ND2 U41 ( .A(\SUMB[44][7] ), .B(n485), .Z(n19) );
  ND3 U42 ( .A(n17), .B(n18), .C(n19), .Z(\CARRYB[45][6] ) );
  FA1AP U43 ( .A(\CARRYB[31][14] ), .B(\ab[32][14] ), .CI(\SUMB[31][15] ), .S(
        n20) );
  EOP U44 ( .A(\CARRYB[10][37] ), .B(n656), .Z(n905) );
  EO3P U45 ( .A(\CARRYB[23][31] ), .B(\ab[31][24] ), .C(\SUMB[23][32] ), .Z(
        \SUMB[24][31] ) );
  EO U46 ( .A(\SUMB[20][36] ), .B(\ab[35][21] ), .Z(n1054) );
  EOP U47 ( .A(\CARRYB[37][29] ), .B(\ab[38][29] ), .Z(n794) );
  EOP U48 ( .A(n2226), .B(n2175), .Z(\SUMB[1][37] ) );
  EOP U49 ( .A(\CARRYB[9][37] ), .B(n599), .Z(n1001) );
  ND2P U50 ( .A(\CARRYB[30][14] ), .B(\ab[31][14] ), .Z(n1190) );
  ND2P U51 ( .A(\CARRYB[30][14] ), .B(\SUMB[30][15] ), .Z(n1189) );
  EO U52 ( .A(\SUMB[43][7] ), .B(n1383), .Z(\SUMB[44][6] ) );
  ND2 U53 ( .A(\SUMB[10][20] ), .B(\CARRYB[10][19] ), .Z(n826) );
  ND2 U54 ( .A(\CARRYB[10][19] ), .B(n618), .Z(n828) );
  EO3P U55 ( .A(\CARRYB[34][8] ), .B(n507), .C(\SUMB[34][9] ), .Z(n21) );
  EOP U56 ( .A(\CARRYB[30][10] ), .B(n585), .Z(n22) );
  EOP U57 ( .A(\SUMB[30][11] ), .B(n22), .Z(\SUMB[31][10] ) );
  ND2 U58 ( .A(\SUMB[30][11] ), .B(\CARRYB[30][10] ), .Z(n23) );
  ND2 U59 ( .A(\SUMB[30][11] ), .B(n585), .Z(n24) );
  ND2 U60 ( .A(\CARRYB[30][10] ), .B(n585), .Z(n25) );
  ND3P U61 ( .A(n23), .B(n24), .C(n25), .Z(\CARRYB[31][10] ) );
  EO3 U62 ( .A(\CARRYB[34][8] ), .B(n507), .C(\SUMB[34][9] ), .Z(\SUMB[35][8] ) );
  ND3 U63 ( .A(n1514), .B(n1515), .C(n1516), .Z(\CARRYB[30][10] ) );
  ND3P U64 ( .A(n1538), .B(n1539), .C(n1540), .Z(\CARRYB[6][26] ) );
  ND3P U65 ( .A(n754), .B(n755), .C(n756), .Z(\CARRYB[26][12] ) );
  ND2P U66 ( .A(\SUMB[11][34] ), .B(\CARRYB[11][33] ), .Z(n1419) );
  ND2P U67 ( .A(\SUMB[11][34] ), .B(n653), .Z(n1420) );
  EOP U68 ( .A(\CARRYB[45][21] ), .B(\ab[46][21] ), .Z(n845) );
  ND3P U69 ( .A(n1927), .B(n1928), .C(n1929), .Z(\CARRYB[18][28] ) );
  ND3 U70 ( .A(n1964), .B(n1965), .C(n1966), .Z(\CARRYB[14][42] ) );
  EO U71 ( .A(n1199), .B(\SUMB[21][35] ), .Z(\SUMB[22][34] ) );
  ND3 U72 ( .A(n155), .B(n156), .C(n157), .Z(\CARRYB[33][9] ) );
  EOP U73 ( .A(\SUMB[21][18] ), .B(n1689), .Z(\SUMB[22][17] ) );
  ND3P U74 ( .A(n1850), .B(n1851), .C(n1852), .Z(\CARRYB[46][21] ) );
  EOP U75 ( .A(\CARRYB[28][24] ), .B(\ab[29][24] ), .Z(n1433) );
  EOP U76 ( .A(\SUMB[13][31] ), .B(n983), .Z(\SUMB[14][30] ) );
  EO3 U77 ( .A(\CARRYB[32][13] ), .B(\ab[33][13] ), .C(n20), .Z(\SUMB[33][13] ) );
  ND2 U78 ( .A(\CARRYB[32][13] ), .B(\SUMB[32][14] ), .Z(n26) );
  ND2 U79 ( .A(\CARRYB[32][13] ), .B(\ab[33][13] ), .Z(n27) );
  ND2 U80 ( .A(\SUMB[32][14] ), .B(\ab[33][13] ), .Z(n28) );
  ND3 U81 ( .A(n26), .B(n27), .C(n28), .Z(\CARRYB[33][13] ) );
  FA1AP U82 ( .A(\CARRYB[37][30] ), .B(\ab[38][30] ), .CI(\SUMB[37][31] ), .S(
        n29) );
  EO3 U83 ( .A(\SUMB[7][39] ), .B(n531), .C(\CARRYB[7][38] ), .Z(\SUMB[8][38] ) );
  ND2P U84 ( .A(\SUMB[7][39] ), .B(\CARRYB[7][38] ), .Z(n30) );
  ND2 U85 ( .A(\SUMB[7][39] ), .B(n531), .Z(n31) );
  ND2P U86 ( .A(\CARRYB[7][38] ), .B(n531), .Z(n32) );
  ND3P U87 ( .A(n30), .B(n31), .C(n32), .Z(\CARRYB[8][38] ) );
  EO U88 ( .A(\SUMB[4][41] ), .B(n432), .Z(n33) );
  EO U89 ( .A(\CARRYB[4][40] ), .B(n33), .Z(\SUMB[5][40] ) );
  AN2 U90 ( .A(\ab[25][25] ), .B(n2117), .Z(n2235) );
  EOP U91 ( .A(\CARRYB[22][9] ), .B(n584), .Z(n1904) );
  ND3P U92 ( .A(n1173), .B(n1174), .C(n1175), .Z(\CARRYB[16][11] ) );
  EOP U93 ( .A(\SUMB[41][5] ), .B(n1814), .Z(\SUMB[42][4] ) );
  EOP U94 ( .A(\SUMB[44][4] ), .B(n1703), .Z(\SUMB[45][3] ) );
  EOP U95 ( .A(\SUMB[25][9] ), .B(n1732), .Z(\SUMB[26][8] ) );
  EOP U96 ( .A(\SUMB[22][10] ), .B(n1904), .Z(\SUMB[23][9] ) );
  AN2P U97 ( .A(n2206), .B(n2200), .Z(\CARRYB[1][42] ) );
  EO U98 ( .A(n2200), .B(n2206), .Z(\SUMB[1][42] ) );
  EOP U99 ( .A(\SUMB[1][43] ), .B(n1404), .Z(\SUMB[2][42] ) );
  ND2P U100 ( .A(\SUMB[33][11] ), .B(n590), .Z(n1392) );
  ND2P U101 ( .A(\SUMB[33][11] ), .B(\CARRYB[33][10] ), .Z(n1391) );
  EOP U102 ( .A(\CARRYB[30][13] ), .B(n685), .Z(n1761) );
  EOP U103 ( .A(\CARRYB[45][19] ), .B(\ab[46][19] ), .Z(n1246) );
  EOP U104 ( .A(\SUMB[45][20] ), .B(n1246), .Z(\SUMB[46][19] ) );
  ND3P U105 ( .A(n118), .B(n119), .C(n120), .Z(\CARRYB[15][26] ) );
  ND2P U106 ( .A(n78), .B(n79), .Z(\SUMB[1][32] ) );
  ND2 U107 ( .A(n1108), .B(n1109), .Z(\SUMB[40][15] ) );
  EO3P U108 ( .A(\CARRYB[26][20] ), .B(\ab[27][20] ), .C(\SUMB[26][21] ), .Z(
        \SUMB[27][20] ) );
  AN2 U109 ( .A(n2175), .B(n2226), .Z(\CARRYB[1][37] ) );
  EOP U110 ( .A(n501), .B(\CARRYB[35][7] ), .Z(n34) );
  EOP U111 ( .A(n34), .B(n21), .Z(\SUMB[36][7] ) );
  ND2 U112 ( .A(\CARRYB[34][8] ), .B(n507), .Z(n35) );
  ND2 U113 ( .A(\CARRYB[34][8] ), .B(\SUMB[34][9] ), .Z(n36) );
  ND2 U114 ( .A(n507), .B(\SUMB[34][9] ), .Z(n37) );
  ND3P U115 ( .A(n35), .B(n36), .C(n37), .Z(\CARRYB[35][8] ) );
  ND2 U116 ( .A(n501), .B(\CARRYB[35][7] ), .Z(n38) );
  ND2 U117 ( .A(n501), .B(\SUMB[35][8] ), .Z(n39) );
  ND2 U118 ( .A(\CARRYB[35][7] ), .B(\SUMB[35][8] ), .Z(n40) );
  ND3P U119 ( .A(n38), .B(n39), .C(n40), .Z(\CARRYB[36][7] ) );
  EO3P U120 ( .A(\CARRYB[27][11] ), .B(n628), .C(\SUMB[27][12] ), .Z(
        \SUMB[28][11] ) );
  ND2 U121 ( .A(\CARRYB[27][11] ), .B(\SUMB[27][12] ), .Z(n41) );
  ND2 U122 ( .A(\CARRYB[27][11] ), .B(n628), .Z(n42) );
  ND2 U123 ( .A(\SUMB[27][12] ), .B(n628), .Z(n43) );
  ND3P U124 ( .A(n41), .B(n42), .C(n43), .Z(\CARRYB[28][11] ) );
  EOP U125 ( .A(\CARRYB[1][21] ), .B(n2264), .Z(n44) );
  EOP U126 ( .A(\SUMB[1][22] ), .B(n44), .Z(\SUMB[2][21] ) );
  ND2P U127 ( .A(\SUMB[1][22] ), .B(\CARRYB[1][21] ), .Z(n45) );
  ND2P U128 ( .A(\SUMB[1][22] ), .B(n2264), .Z(n46) );
  ND2 U129 ( .A(\CARRYB[1][21] ), .B(n2264), .Z(n47) );
  ND3P U130 ( .A(n45), .B(n46), .C(n47), .Z(\CARRYB[2][21] ) );
  IVA U131 ( .A(B[0]), .Z(n48) );
  IVAP U132 ( .A(n48), .Z(n49) );
  EOP U133 ( .A(n697), .B(\CARRYB[12][28] ), .Z(n1132) );
  ND3P U134 ( .A(n1391), .B(n1392), .C(n1393), .Z(\CARRYB[34][10] ) );
  ND3P U135 ( .A(n1558), .B(n1559), .C(n1560), .Z(\CARRYB[31][9] ) );
  EOP U136 ( .A(\SUMB[38][6] ), .B(n938), .Z(\SUMB[39][5] ) );
  EOP U137 ( .A(n531), .B(\CARRYB[37][8] ), .Z(n1336) );
  AN2P U138 ( .A(\ab[30][30] ), .B(n243), .Z(n2169) );
  EO3 U139 ( .A(\CARRYB[15][17] ), .B(\ab[17][16] ), .C(\SUMB[15][18] ), .Z(
        \SUMB[16][17] ) );
  EO3 U140 ( .A(\CARRYB[18][37] ), .B(\ab[37][19] ), .C(\SUMB[18][38] ), .Z(
        \SUMB[19][37] ) );
  ND2P U141 ( .A(\CARRYB[18][37] ), .B(\SUMB[18][38] ), .Z(n50) );
  ND2P U142 ( .A(\CARRYB[18][37] ), .B(\ab[37][19] ), .Z(n51) );
  ND2 U143 ( .A(\SUMB[18][38] ), .B(\ab[37][19] ), .Z(n52) );
  ND3P U144 ( .A(n50), .B(n51), .C(n52), .Z(\CARRYB[19][37] ) );
  EO3 U145 ( .A(\SUMB[20][37] ), .B(\ab[36][21] ), .C(\CARRYB[20][36] ), .Z(
        \SUMB[21][36] ) );
  ND2 U146 ( .A(\SUMB[20][37] ), .B(\CARRYB[20][36] ), .Z(n53) );
  ND2 U147 ( .A(\SUMB[20][37] ), .B(\ab[36][21] ), .Z(n54) );
  ND2 U148 ( .A(\CARRYB[20][36] ), .B(\ab[36][21] ), .Z(n55) );
  ND3P U149 ( .A(n53), .B(n54), .C(n55), .Z(\CARRYB[21][36] ) );
  ND3P U150 ( .A(n1259), .B(n1260), .C(n1261), .Z(\CARRYB[35][14] ) );
  EOP U151 ( .A(\CARRYB[9][20] ), .B(n581), .Z(n1778) );
  EO3 U152 ( .A(\SUMB[21][15] ), .B(n700), .C(\CARRYB[21][14] ), .Z(
        \SUMB[22][14] ) );
  EOP U153 ( .A(\CARRYB[21][17] ), .B(\ab[22][17] ), .Z(n1689) );
  EOP U154 ( .A(\CARRYB[7][20] ), .B(n515), .Z(n1764) );
  EOP U155 ( .A(\CARRYB[32][35] ), .B(\ab[35][33] ), .Z(n56) );
  EOP U156 ( .A(\SUMB[32][36] ), .B(n56), .Z(\SUMB[33][35] ) );
  ND2 U157 ( .A(\SUMB[32][36] ), .B(\CARRYB[32][35] ), .Z(n57) );
  ND2 U158 ( .A(\SUMB[32][36] ), .B(\ab[35][33] ), .Z(n58) );
  ND2 U159 ( .A(\CARRYB[32][35] ), .B(\ab[35][33] ), .Z(n59) );
  ND3P U160 ( .A(n57), .B(n58), .C(n59), .Z(\CARRYB[33][35] ) );
  EOP U161 ( .A(\CARRYB[33][35] ), .B(\ab[35][34] ), .Z(n60) );
  EOP U162 ( .A(\SUMB[33][36] ), .B(n60), .Z(\SUMB[34][35] ) );
  ND2 U163 ( .A(\SUMB[33][36] ), .B(\CARRYB[33][35] ), .Z(n61) );
  ND2 U164 ( .A(\SUMB[33][36] ), .B(\ab[35][34] ), .Z(n62) );
  ND2 U165 ( .A(\CARRYB[33][35] ), .B(\ab[35][34] ), .Z(n63) );
  ND3P U166 ( .A(n61), .B(n62), .C(n63), .Z(\CARRYB[34][35] ) );
  EOP U167 ( .A(\SUMB[29][37] ), .B(\ab[36][30] ), .Z(n64) );
  EOP U168 ( .A(\CARRYB[29][36] ), .B(n64), .Z(\SUMB[30][36] ) );
  ND2 U169 ( .A(\CARRYB[29][36] ), .B(\SUMB[29][37] ), .Z(n65) );
  ND2 U170 ( .A(\CARRYB[29][36] ), .B(\ab[36][30] ), .Z(n66) );
  ND2 U171 ( .A(\SUMB[29][37] ), .B(\ab[36][30] ), .Z(n67) );
  ND3 U172 ( .A(n65), .B(n66), .C(n67), .Z(\CARRYB[30][36] ) );
  EOP U173 ( .A(\SUMB[42][32] ), .B(n979), .Z(\SUMB[43][31] ) );
  EOP U174 ( .A(\CARRYB[42][31] ), .B(\ab[43][31] ), .Z(n979) );
  B4I U175 ( .A(n2031), .Z(n2117) );
  EOP U176 ( .A(\CARRYB[40][15] ), .B(\ab[41][15] ), .Z(n1117) );
  ND3P U177 ( .A(n820), .B(n821), .C(n822), .Z(\CARRYB[29][19] ) );
  EOP U178 ( .A(\CARRYB[26][13] ), .B(n682), .Z(n1525) );
  EOP U179 ( .A(\ab[34][22] ), .B(\CARRYB[21][34] ), .Z(n1199) );
  ND3P U180 ( .A(n1783), .B(n1784), .C(n1785), .Z(\CARRYB[25][16] ) );
  EOP U181 ( .A(\SUMB[32][9] ), .B(n1898), .Z(\SUMB[33][8] ) );
  ND3 U182 ( .A(n2147), .B(n2148), .C(n2149), .Z(\CARRYB[45][1] ) );
  EOP U183 ( .A(\CARRYB[41][2] ), .B(n2153), .Z(\SUMB[42][2] ) );
  EOP U184 ( .A(\SUMB[41][3] ), .B(n2265), .Z(n2153) );
  EOP U185 ( .A(\CARRYB[20][15] ), .B(n829), .Z(\SUMB[21][15] ) );
  ND2 U186 ( .A(\SUMB[39][29] ), .B(\ab[40][28] ), .Z(n230) );
  ND2 U187 ( .A(\CARRYB[16][37] ), .B(\SUMB[16][38] ), .Z(n1101) );
  ND3P U188 ( .A(n1821), .B(n1822), .C(n1823), .Z(\CARRYB[21][15] ) );
  EO U189 ( .A(n1336), .B(\SUMB[37][9] ), .Z(\SUMB[38][8] ) );
  EOP U190 ( .A(\SUMB[45][30] ), .B(n1510), .Z(\SUMB[46][29] ) );
  ND2 U191 ( .A(\SUMB[45][30] ), .B(\ab[46][29] ), .Z(n1512) );
  EO3P U192 ( .A(\CARRYB[10][41] ), .B(\ab[41][11] ), .C(\SUMB[10][42] ), .Z(
        \SUMB[11][41] ) );
  EOP U193 ( .A(\CARRYB[43][25] ), .B(\ab[44][25] ), .Z(n68) );
  EOP U194 ( .A(\SUMB[43][26] ), .B(n68), .Z(\SUMB[44][25] ) );
  ND2 U195 ( .A(\CARRYB[39][28] ), .B(\SUMB[39][29] ), .Z(n228) );
  ND2 U196 ( .A(\CARRYB[39][28] ), .B(\ab[40][28] ), .Z(n229) );
  ND3P U197 ( .A(n1486), .B(n1487), .C(n1488), .Z(\CARRYB[7][35] ) );
  ND2P U198 ( .A(n1500), .B(n1501), .Z(\SUMB[14][21] ) );
  ND2P U199 ( .A(n765), .B(\ab[32][14] ), .Z(n2033) );
  EOP U200 ( .A(\CARRYB[31][25] ), .B(\ab[32][25] ), .Z(n760) );
  ND3P U201 ( .A(n776), .B(n777), .C(n778), .Z(\CARRYB[31][25] ) );
  ND3P U202 ( .A(n881), .B(n882), .C(n883), .Z(\CARRYB[26][27] ) );
  AN2P U203 ( .A(n2233), .B(n334), .Z(\CARRYB[1][38] ) );
  ND3P U204 ( .A(n884), .B(n885), .C(n886), .Z(\CARRYB[46][22] ) );
  ND2P U205 ( .A(\ab[43][26] ), .B(\SUMB[42][27] ), .Z(n947) );
  EO3P U206 ( .A(\SUMB[27][36] ), .B(\ab[35][28] ), .C(\CARRYB[27][35] ), .Z(
        \SUMB[28][35] ) );
  ND3P U207 ( .A(n1155), .B(n1156), .C(n1157), .Z(\CARRYB[29][34] ) );
  ND3P U208 ( .A(n1034), .B(n1035), .C(n1036), .Z(\CARRYB[44][25] ) );
  EO U209 ( .A(\CARRYB[47][32] ), .B(\SUMB[47][33] ), .Z(\A1[78] ) );
  ND3P U210 ( .A(n761), .B(n762), .C(n763), .Z(\CARRYB[32][25] ) );
  B5I U211 ( .A(n1731), .Z(n2233) );
  ND2P U212 ( .A(n1082), .B(n1083), .Z(\SUMB[7][35] ) );
  ND2P U213 ( .A(\SUMB[6][36] ), .B(n1081), .Z(n1082) );
  EOP U214 ( .A(n753), .B(\SUMB[26][12] ), .Z(\SUMB[27][11] ) );
  ND3 U215 ( .A(n1200), .B(n1201), .C(n1202), .Z(\CARRYB[21][35] ) );
  EO3P U216 ( .A(\CARRYB[39][28] ), .B(\ab[40][28] ), .C(\SUMB[39][29] ), .Z(
        \SUMB[40][28] ) );
  ND3P U217 ( .A(n2042), .B(n2043), .C(n2044), .Z(\CARRYB[12][45] ) );
  ND3P U218 ( .A(n1243), .B(n1244), .C(n1245), .Z(\CARRYB[4][45] ) );
  EOP U219 ( .A(n942), .B(\SUMB[42][27] ), .Z(\SUMB[43][26] ) );
  EOP U220 ( .A(\CARRYB[45][15] ), .B(\ab[46][15] ), .Z(n1139) );
  ND2 U221 ( .A(\CARRYB[30][19] ), .B(n914), .Z(n915) );
  IV U222 ( .A(\CARRYB[30][19] ), .Z(n913) );
  ND2 U223 ( .A(\SUMB[4][30] ), .B(\CARRYB[4][29] ), .Z(n73) );
  ND2 U224 ( .A(\SUMB[4][30] ), .B(n411), .Z(n74) );
  ND3P U225 ( .A(n1938), .B(n1939), .C(n1940), .Z(\CARRYB[38][34] ) );
  ND3P U226 ( .A(n1967), .B(n1968), .C(n1969), .Z(\CARRYB[15][41] ) );
  ND3P U227 ( .A(n869), .B(n870), .C(n871), .Z(\CARRYB[47][11] ) );
  ND3P U228 ( .A(n943), .B(n944), .C(n945), .Z(\CARRYB[42][27] ) );
  ND2 U229 ( .A(\CARRYB[1][45] ), .B(\SUMB[1][46] ), .Z(n185) );
  ND2 U230 ( .A(\SUMB[1][46] ), .B(n2247), .Z(n187) );
  ND3P U231 ( .A(n2131), .B(n2132), .C(n2133), .Z(\CARRYB[46][0] ) );
  ND3P U232 ( .A(n1861), .B(n1862), .C(n1863), .Z(\CARRYB[35][0] ) );
  ND3P U233 ( .A(n1865), .B(n1866), .C(n1867), .Z(\CARRYB[36][0] ) );
  EO3P U234 ( .A(\CARRYB[1][45] ), .B(n2247), .C(\SUMB[1][46] ), .Z(
        \SUMB[2][45] ) );
  ND3P U235 ( .A(n1654), .B(n1655), .C(n1656), .Z(\CARRYB[7][28] ) );
  ND3 U236 ( .A(n2067), .B(n2068), .C(n2069), .Z(\CARRYB[4][30] ) );
  ND3P U237 ( .A(n1273), .B(n1274), .C(n1275), .Z(\CARRYB[24][37] ) );
  ND3P U238 ( .A(n1457), .B(n1458), .C(n1459), .Z(\CARRYB[2][44] ) );
  AN2P U239 ( .A(\CARRYB[47][1] ), .B(\SUMB[47][2] ), .Z(\A2[48] ) );
  ND3P U240 ( .A(n1978), .B(n1979), .C(n1980), .Z(\CARRYB[30][2] ) );
  ND3P U241 ( .A(n2128), .B(n2129), .C(n2130), .Z(\CARRYB[35][2] ) );
  ND3P U242 ( .A(n1203), .B(n1204), .C(n1205), .Z(\CARRYB[22][34] ) );
  ND2P U243 ( .A(\ab[34][22] ), .B(\SUMB[21][35] ), .Z(n1204) );
  EOP U244 ( .A(\SUMB[45][32] ), .B(\ab[46][31] ), .Z(n69) );
  EOP U245 ( .A(\CARRYB[45][31] ), .B(n69), .Z(\SUMB[46][31] ) );
  ND2 U246 ( .A(\CARRYB[45][31] ), .B(\SUMB[45][32] ), .Z(n70) );
  ND2 U247 ( .A(\CARRYB[45][31] ), .B(\ab[46][31] ), .Z(n71) );
  ND2 U248 ( .A(\SUMB[45][32] ), .B(\ab[46][31] ), .Z(n72) );
  ND3P U249 ( .A(n70), .B(n71), .C(n72), .Z(\CARRYB[46][31] ) );
  EO3 U250 ( .A(\SUMB[4][30] ), .B(n411), .C(\CARRYB[4][29] ), .Z(
        \SUMB[5][29] ) );
  ND2P U251 ( .A(\CARRYB[4][29] ), .B(n411), .Z(n75) );
  ND3P U252 ( .A(n73), .B(n74), .C(n75), .Z(\CARRYB[5][29] ) );
  ND2P U253 ( .A(n2312), .B(n77), .Z(n78) );
  ND2 U254 ( .A(n76), .B(n1621), .Z(n79) );
  IV U255 ( .A(n2312), .Z(n76) );
  IVP U256 ( .A(n1621), .Z(n77) );
  AN2P U257 ( .A(\ab[33][33] ), .B(n243), .Z(n2312) );
  EOP U258 ( .A(\CARRYB[4][28] ), .B(n412), .Z(n80) );
  EOP U259 ( .A(\SUMB[4][29] ), .B(n80), .Z(\SUMB[5][28] ) );
  ND2 U260 ( .A(\SUMB[4][29] ), .B(\CARRYB[4][28] ), .Z(n81) );
  ND2 U261 ( .A(\SUMB[4][29] ), .B(n412), .Z(n82) );
  ND2 U262 ( .A(\CARRYB[4][28] ), .B(n412), .Z(n83) );
  ND3 U263 ( .A(n81), .B(n82), .C(n83), .Z(\CARRYB[5][28] ) );
  ND2 U264 ( .A(\CARRYB[4][40] ), .B(\SUMB[4][41] ), .Z(n84) );
  ND2 U265 ( .A(\CARRYB[4][40] ), .B(n432), .Z(n85) );
  ND2 U266 ( .A(\SUMB[4][41] ), .B(n432), .Z(n86) );
  ND3 U267 ( .A(n84), .B(n85), .C(n86), .Z(\CARRYB[5][40] ) );
  EO3P U268 ( .A(\ab[36][24] ), .B(\CARRYB[23][36] ), .C(\SUMB[23][37] ), .Z(
        \SUMB[24][36] ) );
  EOP U269 ( .A(\ab[35][25] ), .B(\CARRYB[24][35] ), .Z(n87) );
  EOP U270 ( .A(n87), .B(\SUMB[24][36] ), .Z(\SUMB[25][35] ) );
  ND2 U271 ( .A(\ab[36][24] ), .B(\CARRYB[23][36] ), .Z(n88) );
  ND2 U272 ( .A(\ab[36][24] ), .B(\SUMB[23][37] ), .Z(n89) );
  ND2 U273 ( .A(\CARRYB[23][36] ), .B(\SUMB[23][37] ), .Z(n90) );
  ND3 U274 ( .A(n88), .B(n89), .C(n90), .Z(\CARRYB[24][36] ) );
  ND2 U275 ( .A(\ab[35][25] ), .B(\CARRYB[24][35] ), .Z(n91) );
  ND2P U276 ( .A(\ab[35][25] ), .B(\SUMB[24][36] ), .Z(n92) );
  ND2P U277 ( .A(\CARRYB[24][35] ), .B(\SUMB[24][36] ), .Z(n93) );
  ND3P U278 ( .A(n91), .B(n92), .C(n93), .Z(\CARRYB[25][35] ) );
  EO3 U279 ( .A(\CARRYB[24][22] ), .B(\ab[25][22] ), .C(\SUMB[24][23] ), .Z(
        \SUMB[25][22] ) );
  ND2 U280 ( .A(\CARRYB[24][22] ), .B(\SUMB[24][23] ), .Z(n94) );
  ND2 U281 ( .A(\CARRYB[24][22] ), .B(\ab[25][22] ), .Z(n95) );
  ND2 U282 ( .A(\SUMB[24][23] ), .B(\ab[25][22] ), .Z(n96) );
  ND3 U283 ( .A(n94), .B(n95), .C(n96), .Z(\CARRYB[25][22] ) );
  EO3P U284 ( .A(\CARRYB[28][40] ), .B(\ab[40][29] ), .C(\SUMB[28][41] ), .Z(
        \SUMB[29][40] ) );
  ND2 U285 ( .A(\CARRYB[28][40] ), .B(\SUMB[28][41] ), .Z(n97) );
  ND2 U286 ( .A(\CARRYB[28][40] ), .B(\ab[40][29] ), .Z(n98) );
  ND2 U287 ( .A(\SUMB[28][41] ), .B(\ab[40][29] ), .Z(n99) );
  ND3P U288 ( .A(n97), .B(n98), .C(n99), .Z(\CARRYB[29][40] ) );
  EO3P U289 ( .A(\SUMB[14][23] ), .B(n720), .C(\CARRYB[14][22] ), .Z(
        \SUMB[15][22] ) );
  ND2 U290 ( .A(\CARRYB[14][22] ), .B(\SUMB[14][23] ), .Z(n100) );
  ND2 U291 ( .A(\CARRYB[14][22] ), .B(n720), .Z(n101) );
  ND2 U292 ( .A(\SUMB[14][23] ), .B(n720), .Z(n102) );
  ND3 U293 ( .A(n100), .B(n101), .C(n102), .Z(\CARRYB[15][22] ) );
  EO U294 ( .A(\ab[46][22] ), .B(\ab[47][21] ), .Z(n103) );
  EOP U295 ( .A(\CARRYB[21][46] ), .B(n103), .Z(\SUMB[22][46] ) );
  ND2P U296 ( .A(\CARRYB[21][46] ), .B(\ab[46][22] ), .Z(n104) );
  ND2P U297 ( .A(\CARRYB[21][46] ), .B(\ab[47][21] ), .Z(n105) );
  ND2 U298 ( .A(\ab[46][22] ), .B(\ab[47][21] ), .Z(n106) );
  ND3P U299 ( .A(n104), .B(n105), .C(n106), .Z(\CARRYB[22][46] ) );
  EOP U300 ( .A(\SUMB[26][35] ), .B(\ab[34][27] ), .Z(n107) );
  EOP U301 ( .A(\CARRYB[26][34] ), .B(n107), .Z(\SUMB[27][34] ) );
  ND2 U302 ( .A(\CARRYB[26][34] ), .B(\SUMB[26][35] ), .Z(n108) );
  ND2 U303 ( .A(\CARRYB[26][34] ), .B(\ab[34][27] ), .Z(n109) );
  ND2 U304 ( .A(\SUMB[26][35] ), .B(\ab[34][27] ), .Z(n110) );
  ND3P U305 ( .A(n108), .B(n109), .C(n110), .Z(\CARRYB[27][34] ) );
  EO3 U306 ( .A(\CARRYB[19][39] ), .B(\ab[39][20] ), .C(\SUMB[19][40] ), .Z(
        \SUMB[20][39] ) );
  ND2 U307 ( .A(\CARRYB[19][39] ), .B(\SUMB[19][40] ), .Z(n111) );
  ND2 U308 ( .A(\CARRYB[19][39] ), .B(\ab[39][20] ), .Z(n112) );
  ND2 U309 ( .A(\SUMB[19][40] ), .B(\ab[39][20] ), .Z(n113) );
  ND3P U310 ( .A(n111), .B(n112), .C(n113), .Z(\CARRYB[20][39] ) );
  EO3P U311 ( .A(\CARRYB[18][40] ), .B(\ab[40][19] ), .C(\SUMB[18][41] ), .Z(
        \SUMB[19][40] ) );
  EO3P U312 ( .A(\CARRYB[30][35] ), .B(\ab[35][31] ), .C(\SUMB[30][36] ), .Z(
        \SUMB[31][35] ) );
  ND2 U313 ( .A(\CARRYB[30][35] ), .B(\SUMB[30][36] ), .Z(n114) );
  ND2 U314 ( .A(\CARRYB[30][35] ), .B(\ab[35][31] ), .Z(n115) );
  ND2 U315 ( .A(\SUMB[30][36] ), .B(\ab[35][31] ), .Z(n116) );
  ND3P U316 ( .A(n114), .B(n115), .C(n116), .Z(\CARRYB[31][35] ) );
  EOP U317 ( .A(\SUMB[9][28] ), .B(n611), .Z(n117) );
  EOP U318 ( .A(\CARRYB[9][27] ), .B(n117), .Z(\SUMB[10][27] ) );
  EO3 U319 ( .A(\CARRYB[14][26] ), .B(n715), .C(\SUMB[14][27] ), .Z(
        \SUMB[15][26] ) );
  ND2 U320 ( .A(\CARRYB[14][26] ), .B(\SUMB[14][27] ), .Z(n118) );
  ND2 U321 ( .A(\CARRYB[14][26] ), .B(n715), .Z(n119) );
  ND2 U322 ( .A(\SUMB[14][27] ), .B(n715), .Z(n120) );
  EO3P U323 ( .A(\SUMB[45][24] ), .B(\ab[46][23] ), .C(\CARRYB[45][23] ), .Z(
        \SUMB[46][23] ) );
  ND2 U324 ( .A(\CARRYB[45][23] ), .B(\SUMB[45][24] ), .Z(n121) );
  ND2 U325 ( .A(\CARRYB[45][23] ), .B(\ab[46][23] ), .Z(n122) );
  ND2 U326 ( .A(\SUMB[45][24] ), .B(\ab[46][23] ), .Z(n123) );
  ND3 U327 ( .A(n121), .B(n122), .C(n123), .Z(\CARRYB[46][23] ) );
  EOP U328 ( .A(\SUMB[39][18] ), .B(\ab[40][17] ), .Z(n124) );
  EOP U329 ( .A(\CARRYB[39][17] ), .B(n124), .Z(\SUMB[40][17] ) );
  EO U330 ( .A(\CARRYB[26][31] ), .B(\ab[31][27] ), .Z(n125) );
  EO U331 ( .A(\SUMB[26][32] ), .B(n125), .Z(\SUMB[27][31] ) );
  EOP U332 ( .A(\CARRYB[32][17] ), .B(\ab[33][17] ), .Z(n126) );
  EOP U333 ( .A(\SUMB[32][18] ), .B(n126), .Z(\SUMB[33][17] ) );
  ND3P U334 ( .A(n1270), .B(n1271), .C(n1272), .Z(\CARRYB[32][17] ) );
  EO3P U335 ( .A(n2251), .B(\CARRYB[40][2] ), .C(\SUMB[40][3] ), .Z(
        \SUMB[41][2] ) );
  EO U336 ( .A(n2206), .B(\CARRYB[41][1] ), .Z(n127) );
  EO U337 ( .A(n127), .B(\SUMB[41][2] ), .Z(\SUMB[42][1] ) );
  ND2 U338 ( .A(n2251), .B(\CARRYB[40][2] ), .Z(n128) );
  ND2 U339 ( .A(n2251), .B(\SUMB[40][3] ), .Z(n129) );
  ND2 U340 ( .A(\CARRYB[40][2] ), .B(\SUMB[40][3] ), .Z(n130) );
  ND3P U341 ( .A(n128), .B(n129), .C(n130), .Z(\CARRYB[41][2] ) );
  ND2 U342 ( .A(n2206), .B(\CARRYB[41][1] ), .Z(n131) );
  ND2P U343 ( .A(n2206), .B(\SUMB[41][2] ), .Z(n132) );
  ND2P U344 ( .A(\CARRYB[41][1] ), .B(\SUMB[41][2] ), .Z(n133) );
  ND3P U345 ( .A(n131), .B(n132), .C(n133), .Z(\CARRYB[42][1] ) );
  EOP U346 ( .A(\SUMB[33][21] ), .B(\ab[34][20] ), .Z(n134) );
  EOP U347 ( .A(\CARRYB[33][20] ), .B(n134), .Z(\SUMB[34][20] ) );
  ND2 U348 ( .A(\CARRYB[33][20] ), .B(\SUMB[33][21] ), .Z(n135) );
  ND2 U349 ( .A(\CARRYB[33][20] ), .B(\ab[34][20] ), .Z(n136) );
  ND2 U350 ( .A(\SUMB[33][21] ), .B(\ab[34][20] ), .Z(n137) );
  ND3P U351 ( .A(n135), .B(n136), .C(n137), .Z(\CARRYB[34][20] ) );
  EOP U352 ( .A(\CARRYB[34][20] ), .B(\ab[35][20] ), .Z(n930) );
  EO3 U353 ( .A(\CARRYB[4][11] ), .B(n418), .C(\SUMB[4][12] ), .Z(
        \SUMB[5][11] ) );
  ND2 U354 ( .A(\CARRYB[4][11] ), .B(\SUMB[4][12] ), .Z(n138) );
  ND2 U355 ( .A(\CARRYB[4][11] ), .B(n418), .Z(n139) );
  ND2 U356 ( .A(\SUMB[4][12] ), .B(n418), .Z(n140) );
  ND3P U357 ( .A(n138), .B(n139), .C(n140), .Z(\CARRYB[5][11] ) );
  EOP U358 ( .A(\SUMB[10][34] ), .B(n636), .Z(n141) );
  EOP U359 ( .A(\CARRYB[10][33] ), .B(n141), .Z(\SUMB[11][33] ) );
  ND2 U360 ( .A(\CARRYB[10][33] ), .B(\SUMB[10][34] ), .Z(n142) );
  ND2 U361 ( .A(\CARRYB[10][33] ), .B(n636), .Z(n143) );
  ND2 U362 ( .A(\SUMB[10][34] ), .B(n636), .Z(n144) );
  ND3P U363 ( .A(n142), .B(n143), .C(n144), .Z(\CARRYB[11][33] ) );
  EO3P U364 ( .A(\CARRYB[22][43] ), .B(\ab[43][23] ), .C(\SUMB[22][44] ), .Z(
        \SUMB[23][43] ) );
  ND2 U365 ( .A(\CARRYB[22][43] ), .B(\SUMB[22][44] ), .Z(n145) );
  ND2 U366 ( .A(\CARRYB[22][43] ), .B(\ab[43][23] ), .Z(n146) );
  ND2 U367 ( .A(\SUMB[22][44] ), .B(\ab[43][23] ), .Z(n147) );
  ND3P U368 ( .A(n145), .B(n146), .C(n147), .Z(\CARRYB[23][43] ) );
  EO3P U369 ( .A(\CARRYB[44][38] ), .B(\ab[45][38] ), .C(\SUMB[44][39] ), .Z(
        \SUMB[45][38] ) );
  ND2 U370 ( .A(\CARRYB[44][38] ), .B(\SUMB[44][39] ), .Z(n148) );
  ND2 U371 ( .A(\CARRYB[44][38] ), .B(\ab[45][38] ), .Z(n149) );
  ND2 U372 ( .A(\SUMB[44][39] ), .B(\ab[45][38] ), .Z(n150) );
  ND3P U373 ( .A(n148), .B(n149), .C(n150), .Z(\CARRYB[45][38] ) );
  EO3 U374 ( .A(\SUMB[13][35] ), .B(\ab[34][14] ), .C(\CARRYB[13][34] ), .Z(
        \SUMB[14][34] ) );
  ND2 U375 ( .A(\SUMB[13][35] ), .B(\CARRYB[13][34] ), .Z(n151) );
  ND2 U376 ( .A(\SUMB[13][35] ), .B(\ab[34][14] ), .Z(n152) );
  ND2 U377 ( .A(\CARRYB[13][34] ), .B(\ab[34][14] ), .Z(n153) );
  ND3 U378 ( .A(n151), .B(n152), .C(n153), .Z(\CARRYB[14][34] ) );
  EOP U379 ( .A(\SUMB[32][10] ), .B(n558), .Z(n154) );
  EOP U380 ( .A(\CARRYB[32][9] ), .B(n154), .Z(\SUMB[33][9] ) );
  ND2 U381 ( .A(\CARRYB[32][9] ), .B(\SUMB[32][10] ), .Z(n155) );
  ND2 U382 ( .A(\CARRYB[32][9] ), .B(n558), .Z(n156) );
  ND2 U383 ( .A(\SUMB[32][10] ), .B(n558), .Z(n157) );
  ND2 U384 ( .A(\CARRYB[32][17] ), .B(\SUMB[32][18] ), .Z(n158) );
  ND2 U385 ( .A(\CARRYB[32][17] ), .B(\ab[33][17] ), .Z(n159) );
  ND2 U386 ( .A(\SUMB[32][18] ), .B(\ab[33][17] ), .Z(n160) );
  ND3 U387 ( .A(n158), .B(n159), .C(n160), .Z(\CARRYB[33][17] ) );
  EO3 U388 ( .A(\CARRYB[32][41] ), .B(\ab[41][33] ), .C(\SUMB[32][42] ), .Z(
        \SUMB[33][41] ) );
  ND2 U389 ( .A(\CARRYB[32][41] ), .B(\SUMB[32][42] ), .Z(n161) );
  ND2 U390 ( .A(\CARRYB[32][41] ), .B(\ab[41][33] ), .Z(n162) );
  ND2 U391 ( .A(\SUMB[32][42] ), .B(\ab[41][33] ), .Z(n163) );
  ND3P U392 ( .A(n161), .B(n162), .C(n163), .Z(\CARRYB[33][41] ) );
  EO3P U393 ( .A(\ab[40][15] ), .B(\CARRYB[14][40] ), .C(\SUMB[14][41] ), .Z(
        \SUMB[15][40] ) );
  EOP U394 ( .A(\CARRYB[15][39] ), .B(\ab[39][16] ), .Z(n164) );
  EOP U395 ( .A(n164), .B(\SUMB[15][40] ), .Z(\SUMB[16][39] ) );
  ND2 U396 ( .A(\ab[40][15] ), .B(\CARRYB[14][40] ), .Z(n165) );
  ND2 U397 ( .A(\ab[40][15] ), .B(\SUMB[14][41] ), .Z(n166) );
  ND2 U398 ( .A(\CARRYB[14][40] ), .B(\SUMB[14][41] ), .Z(n167) );
  ND3 U399 ( .A(n165), .B(n166), .C(n167), .Z(\CARRYB[15][40] ) );
  ND2 U400 ( .A(\CARRYB[15][39] ), .B(\ab[39][16] ), .Z(n168) );
  ND2P U401 ( .A(\CARRYB[15][39] ), .B(\SUMB[15][40] ), .Z(n169) );
  ND2P U402 ( .A(\ab[39][16] ), .B(\SUMB[15][40] ), .Z(n170) );
  ND3P U403 ( .A(n168), .B(n169), .C(n170), .Z(\CARRYB[16][39] ) );
  ND2 U404 ( .A(\CARRYB[18][40] ), .B(\SUMB[18][41] ), .Z(n171) );
  ND2 U405 ( .A(\CARRYB[18][40] ), .B(\ab[40][19] ), .Z(n172) );
  ND2 U406 ( .A(\SUMB[18][41] ), .B(\ab[40][19] ), .Z(n173) );
  ND3P U407 ( .A(n171), .B(n172), .C(n173), .Z(\CARRYB[19][40] ) );
  EO3P U408 ( .A(\CARRYB[4][39] ), .B(n396), .C(\SUMB[4][40] ), .Z(
        \SUMB[5][39] ) );
  EOP U409 ( .A(n456), .B(\CARRYB[5][38] ), .Z(n174) );
  EOP U410 ( .A(n174), .B(\SUMB[5][39] ), .Z(\SUMB[6][38] ) );
  ND2 U411 ( .A(n396), .B(\CARRYB[4][39] ), .Z(n175) );
  ND2 U412 ( .A(n396), .B(\SUMB[4][40] ), .Z(n176) );
  ND2 U413 ( .A(\CARRYB[4][39] ), .B(\SUMB[4][40] ), .Z(n177) );
  ND3 U414 ( .A(n175), .B(n176), .C(n177), .Z(\CARRYB[5][39] ) );
  ND2 U415 ( .A(n456), .B(\CARRYB[5][38] ), .Z(n178) );
  ND2P U416 ( .A(n456), .B(\SUMB[5][39] ), .Z(n179) );
  ND2P U417 ( .A(\CARRYB[5][38] ), .B(\SUMB[5][39] ), .Z(n180) );
  ND3P U418 ( .A(n178), .B(n179), .C(n180), .Z(\CARRYB[6][38] ) );
  EOP U419 ( .A(\CARRYB[3][43] ), .B(n389), .Z(n181) );
  EOP U420 ( .A(\SUMB[3][44] ), .B(n181), .Z(\SUMB[4][43] ) );
  ND2 U421 ( .A(\SUMB[3][44] ), .B(\CARRYB[3][43] ), .Z(n182) );
  ND2 U422 ( .A(\SUMB[3][44] ), .B(n389), .Z(n183) );
  ND2 U423 ( .A(\CARRYB[3][43] ), .B(n389), .Z(n184) );
  ND3P U424 ( .A(n182), .B(n183), .C(n184), .Z(\CARRYB[4][43] ) );
  ND2P U425 ( .A(\CARRYB[1][45] ), .B(n2247), .Z(n186) );
  ND3P U426 ( .A(n185), .B(n186), .C(n187), .Z(\CARRYB[2][45] ) );
  EOP U427 ( .A(\CARRYB[40][24] ), .B(\ab[41][24] ), .Z(n188) );
  EOP U428 ( .A(\SUMB[40][25] ), .B(n188), .Z(\SUMB[41][24] ) );
  ND2P U429 ( .A(\SUMB[10][28] ), .B(n190), .Z(n191) );
  ND2 U430 ( .A(n189), .B(n860), .Z(n192) );
  ND2P U431 ( .A(n191), .B(n192), .Z(\SUMB[11][27] ) );
  IVDA U432 ( .A(\SUMB[10][28] ), .Y(n189) );
  IV U433 ( .A(n860), .Z(n190) );
  FA1AP U434 ( .A(\CARRYB[11][26] ), .B(n657), .CI(\SUMB[11][27] ), .S(n786)
         );
  EOP U435 ( .A(\SUMB[19][36] ), .B(\ab[35][20] ), .Z(n193) );
  EOP U436 ( .A(\CARRYB[19][35] ), .B(n193), .Z(\SUMB[20][35] ) );
  ND2P U437 ( .A(\CARRYB[19][35] ), .B(\SUMB[19][36] ), .Z(n194) );
  ND2P U438 ( .A(\CARRYB[19][35] ), .B(\ab[35][20] ), .Z(n195) );
  ND2 U439 ( .A(\SUMB[19][36] ), .B(\ab[35][20] ), .Z(n196) );
  ND3P U440 ( .A(n194), .B(n195), .C(n196), .Z(\CARRYB[20][35] ) );
  EOP U441 ( .A(\CARRYB[45][11] ), .B(\ab[46][11] ), .Z(n197) );
  EOP U442 ( .A(\SUMB[45][12] ), .B(n197), .Z(\SUMB[46][11] ) );
  ND2 U443 ( .A(\SUMB[45][12] ), .B(\CARRYB[45][11] ), .Z(n198) );
  ND2 U444 ( .A(\SUMB[45][12] ), .B(\ab[46][11] ), .Z(n199) );
  ND2 U445 ( .A(\CARRYB[45][11] ), .B(\ab[46][11] ), .Z(n200) );
  ND3P U446 ( .A(n198), .B(n199), .C(n200), .Z(\CARRYB[46][11] ) );
  ND2 U447 ( .A(\CARRYB[10][41] ), .B(\ab[41][11] ), .Z(n201) );
  ND2 U448 ( .A(\CARRYB[10][41] ), .B(\SUMB[10][42] ), .Z(n202) );
  ND2 U449 ( .A(\ab[41][11] ), .B(\SUMB[10][42] ), .Z(n203) );
  ND3 U450 ( .A(n201), .B(n202), .C(n203), .Z(\CARRYB[11][41] ) );
  EOP U451 ( .A(\ab[41][12] ), .B(\SUMB[11][42] ), .Z(n204) );
  EOP U452 ( .A(n204), .B(\CARRYB[11][41] ), .Z(\SUMB[12][41] ) );
  ND2 U453 ( .A(\ab[41][12] ), .B(\SUMB[11][42] ), .Z(n205) );
  ND2 U454 ( .A(\ab[41][12] ), .B(\CARRYB[11][41] ), .Z(n206) );
  ND2 U455 ( .A(\SUMB[11][42] ), .B(\CARRYB[11][41] ), .Z(n207) );
  ND3 U456 ( .A(n205), .B(n206), .C(n207), .Z(\CARRYB[12][41] ) );
  EOP U457 ( .A(\CARRYB[21][39] ), .B(\ab[39][22] ), .Z(n208) );
  EOP U458 ( .A(\SUMB[21][40] ), .B(n208), .Z(\SUMB[22][39] ) );
  ND2 U459 ( .A(\SUMB[21][40] ), .B(\CARRYB[21][39] ), .Z(n209) );
  ND2 U460 ( .A(\SUMB[21][40] ), .B(\ab[39][22] ), .Z(n210) );
  ND2 U461 ( .A(\CARRYB[21][39] ), .B(\ab[39][22] ), .Z(n211) );
  ND3P U462 ( .A(n209), .B(n210), .C(n211), .Z(\CARRYB[22][39] ) );
  ND3P U463 ( .A(n1461), .B(n1462), .C(n1463), .Z(\CARRYB[21][39] ) );
  EO U464 ( .A(\SUMB[37][19] ), .B(\ab[38][18] ), .Z(n212) );
  EO U465 ( .A(\CARRYB[37][18] ), .B(n212), .Z(\SUMB[38][18] ) );
  ND2 U466 ( .A(\CARRYB[37][18] ), .B(\SUMB[37][19] ), .Z(n213) );
  ND2 U467 ( .A(\CARRYB[37][18] ), .B(\ab[38][18] ), .Z(n214) );
  ND2 U468 ( .A(\SUMB[37][19] ), .B(\ab[38][18] ), .Z(n215) );
  ND3P U469 ( .A(n213), .B(n214), .C(n215), .Z(\CARRYB[38][18] ) );
  EOP U470 ( .A(\CARRYB[13][36] ), .B(\ab[36][14] ), .Z(n216) );
  EOP U471 ( .A(\SUMB[13][37] ), .B(n216), .Z(\SUMB[14][36] ) );
  EOP U472 ( .A(n738), .B(\SUMB[14][36] ), .Z(\SUMB[15][35] ) );
  ND2 U473 ( .A(\CARRYB[14][35] ), .B(\SUMB[14][36] ), .Z(n744) );
  ND2P U474 ( .A(\ab[35][15] ), .B(\SUMB[14][36] ), .Z(n743) );
  EO U475 ( .A(\SUMB[14][1] ), .B(n333), .Z(n217) );
  EO U476 ( .A(\CARRYB[14][0] ), .B(n217), .Z(\A1[13] ) );
  ND2 U477 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(n218) );
  ND2 U478 ( .A(\CARRYB[14][0] ), .B(n333), .Z(n219) );
  ND2 U479 ( .A(\SUMB[14][1] ), .B(n333), .Z(n220) );
  ND3 U480 ( .A(n218), .B(n219), .C(n220), .Z(\CARRYB[15][0] ) );
  EO3 U481 ( .A(\CARRYB[13][3] ), .B(n341), .C(\SUMB[13][4] ), .Z(
        \SUMB[14][3] ) );
  ND2 U482 ( .A(\CARRYB[13][3] ), .B(\SUMB[13][4] ), .Z(n221) );
  ND2 U483 ( .A(\CARRYB[13][3] ), .B(n341), .Z(n222) );
  ND2 U484 ( .A(\SUMB[13][4] ), .B(n341), .Z(n223) );
  ND3P U485 ( .A(n221), .B(n222), .C(n223), .Z(\CARRYB[14][3] ) );
  EOP U486 ( .A(\SUMB[46][6] ), .B(n303), .Z(n224) );
  EOP U487 ( .A(\CARRYB[46][5] ), .B(n224), .Z(\SUMB[47][5] ) );
  ND2 U488 ( .A(\CARRYB[46][5] ), .B(\SUMB[46][6] ), .Z(n225) );
  ND2 U489 ( .A(\CARRYB[46][5] ), .B(n303), .Z(n226) );
  ND2 U490 ( .A(\SUMB[46][6] ), .B(n303), .Z(n227) );
  ND3 U491 ( .A(n225), .B(n226), .C(n227), .Z(\CARRYB[47][5] ) );
  ND3P U492 ( .A(n1445), .B(n1446), .C(n1447), .Z(\CARRYB[46][5] ) );
  ND3P U493 ( .A(n228), .B(n229), .C(n230), .Z(\CARRYB[40][28] ) );
  ND2 U494 ( .A(\CARRYB[40][28] ), .B(\ab[41][28] ), .Z(n1317) );
  ND2 U495 ( .A(\SUMB[40][29] ), .B(\CARRYB[40][28] ), .Z(n1315) );
  EO3 U496 ( .A(\SUMB[40][29] ), .B(\ab[41][28] ), .C(\CARRYB[40][28] ), .Z(
        \SUMB[41][28] ) );
  EO3P U497 ( .A(\CARRYB[31][42] ), .B(\ab[42][32] ), .C(\SUMB[31][43] ), .Z(
        \SUMB[32][42] ) );
  ND2 U498 ( .A(\CARRYB[31][42] ), .B(\SUMB[31][43] ), .Z(n231) );
  ND2 U499 ( .A(\CARRYB[31][42] ), .B(\ab[42][32] ), .Z(n232) );
  ND2 U500 ( .A(\SUMB[31][43] ), .B(\ab[42][32] ), .Z(n233) );
  ND3 U501 ( .A(n231), .B(n232), .C(n233), .Z(\CARRYB[32][42] ) );
  EO3P U502 ( .A(\CARRYB[23][5] ), .B(n421), .C(\SUMB[23][6] ), .Z(
        \SUMB[24][5] ) );
  ND2 U503 ( .A(\CARRYB[23][5] ), .B(\SUMB[23][6] ), .Z(n234) );
  ND2 U504 ( .A(\CARRYB[23][5] ), .B(n421), .Z(n235) );
  ND2 U505 ( .A(\SUMB[23][6] ), .B(n421), .Z(n236) );
  ND3P U506 ( .A(n234), .B(n235), .C(n236), .Z(\CARRYB[24][5] ) );
  EO3 U507 ( .A(\CARRYB[16][25] ), .B(\ab[25][17] ), .C(\SUMB[16][26] ), .Z(
        \SUMB[17][25] ) );
  ND2 U508 ( .A(\CARRYB[16][25] ), .B(\SUMB[16][26] ), .Z(n237) );
  ND2 U509 ( .A(\CARRYB[16][25] ), .B(\ab[25][17] ), .Z(n238) );
  ND2 U510 ( .A(\SUMB[16][26] ), .B(\ab[25][17] ), .Z(n239) );
  ND3 U511 ( .A(n237), .B(n238), .C(n239), .Z(\CARRYB[17][25] ) );
  ND2 U512 ( .A(\CARRYB[26][31] ), .B(\SUMB[26][32] ), .Z(n240) );
  ND2 U513 ( .A(\CARRYB[26][31] ), .B(\ab[31][27] ), .Z(n241) );
  ND2 U514 ( .A(\SUMB[26][32] ), .B(\ab[31][27] ), .Z(n242) );
  ND3P U515 ( .A(n240), .B(n241), .C(n242), .Z(\CARRYB[27][31] ) );
  ND3P U516 ( .A(n1888), .B(n1889), .C(n1890), .Z(\CARRYB[18][36] ) );
  ND3P U517 ( .A(n1012), .B(n1013), .C(n1014), .Z(\CARRYB[44][16] ) );
  EOP U518 ( .A(n1537), .B(\SUMB[6][26] ), .Z(\SUMB[7][25] ) );
  EOP U519 ( .A(\CARRYB[28][19] ), .B(n819), .Z(\SUMB[29][19] ) );
  EOP U520 ( .A(\SUMB[28][20] ), .B(\ab[29][19] ), .Z(n819) );
  ND3P U521 ( .A(n917), .B(n918), .C(n919), .Z(\CARRYB[3][24] ) );
  EOP U522 ( .A(\SUMB[26][34] ), .B(n949), .Z(\SUMB[27][33] ) );
  EOP U523 ( .A(\CARRYB[26][33] ), .B(\ab[33][27] ), .Z(n949) );
  EOP U524 ( .A(\CARRYB[47][30] ), .B(\SUMB[47][31] ), .Z(\A1[76] ) );
  EOP U525 ( .A(\CARRYB[45][32] ), .B(n1984), .Z(\SUMB[46][32] ) );
  ND3P U526 ( .A(n1952), .B(n1953), .C(n1954), .Z(\CARRYB[20][43] ) );
  B4IP U527 ( .A(n2031), .Z(PRODUCT[0]) );
  EOP U528 ( .A(n2225), .B(n2222), .Z(\SUMB[1][41] ) );
  EOP U529 ( .A(\CARRYB[28][34] ), .B(\ab[34][29] ), .Z(n1154) );
  ND2P U530 ( .A(\CARRYB[13][36] ), .B(\ab[36][14] ), .Z(n739) );
  B5I U531 ( .A(n2422), .Z(n2421) );
  IV U532 ( .A(\ab[47][47] ), .Z(n2422) );
  EOP U533 ( .A(n2171), .B(n2186), .Z(\SUMB[1][28] ) );
  ND2 U534 ( .A(\CARRYB[30][3] ), .B(n2268), .Z(n2021) );
  B3IP U535 ( .A(B[0]), .Z1(n2031), .Z2(n243) );
  ND3P U536 ( .A(n2020), .B(n2021), .C(n2022), .Z(\CARRYB[31][3] ) );
  ND2 U537 ( .A(\SUMB[45][30] ), .B(\CARRYB[45][29] ), .Z(n1511) );
  EOP U538 ( .A(\CARRYB[45][29] ), .B(\ab[46][29] ), .Z(n1510) );
  EO3P U539 ( .A(\CARRYB[15][37] ), .B(\ab[37][16] ), .C(\SUMB[15][38] ), .Z(
        \SUMB[16][37] ) );
  ND3P U540 ( .A(n2046), .B(n2047), .C(n2048), .Z(\CARRYB[38][1] ) );
  ND3P U541 ( .A(n2055), .B(n2056), .C(n2057), .Z(\CARRYB[17][43] ) );
  EOP U542 ( .A(\CARRYB[1][46] ), .B(n852), .Z(\SUMB[2][46] ) );
  AN2P U543 ( .A(A[47]), .B(n2335), .Z(\ab[7][47] ) );
  B4IP U544 ( .A(\ab[2][2] ), .Z(n2324) );
  EOP U545 ( .A(n2257), .B(n2245), .Z(n852) );
  AN2 U546 ( .A(n2196), .B(n2246), .Z(\CARRYB[1][46] ) );
  ND3P U547 ( .A(n853), .B(n854), .C(n855), .Z(\CARRYB[2][46] ) );
  EOP U548 ( .A(\SUMB[14][44] ), .B(\ab[43][15] ), .Z(n1843) );
  ND2P U549 ( .A(\CARRYB[14][43] ), .B(\ab[43][15] ), .Z(n1845) );
  EOP U550 ( .A(\CARRYB[14][43] ), .B(n1843), .Z(\SUMB[15][43] ) );
  ND3P U551 ( .A(n1844), .B(n1845), .C(n1846), .Z(\CARRYB[15][43] ) );
  EOP U552 ( .A(\CARRYB[19][43] ), .B(n1951), .Z(\SUMB[20][43] ) );
  EOP U553 ( .A(\CARRYB[47][43] ), .B(\SUMB[47][44] ), .Z(\A1[89] ) );
  EOP U554 ( .A(\SUMB[3][46] ), .B(n1242), .Z(\SUMB[4][45] ) );
  EOP U555 ( .A(\CARRYB[3][45] ), .B(n360), .Z(n1242) );
  ND3P U556 ( .A(n1615), .B(n1616), .C(n1617), .Z(\CARRYB[4][44] ) );
  EOP U557 ( .A(\CARRYB[47][44] ), .B(\SUMB[47][45] ), .Z(\A1[90] ) );
  AN2 U558 ( .A(\CARRYB[47][41] ), .B(\SUMB[47][42] ), .Z(\A2[88] ) );
  ND3 U559 ( .A(n1697), .B(n1698), .C(n1699), .Z(\CARRYB[25][29] ) );
  ND2 U560 ( .A(\SUMB[3][33] ), .B(n358), .Z(n1112) );
  ND2 U561 ( .A(\SUMB[7][32] ), .B(\CARRYB[7][31] ), .Z(n1060) );
  ND2 U562 ( .A(\CARRYB[27][37] ), .B(\ab[37][28] ), .Z(n1834) );
  ND2 U563 ( .A(\CARRYB[25][24] ), .B(\ab[26][24] ), .Z(n1580) );
  ND2 U564 ( .A(\CARRYB[3][16] ), .B(n359), .Z(n1772) );
  EO U565 ( .A(\SUMB[3][20] ), .B(n834), .Z(\SUMB[4][19] ) );
  EO U566 ( .A(\CARRYB[3][19] ), .B(n2301), .Z(n834) );
  ND2 U567 ( .A(\CARRYB[28][19] ), .B(\SUMB[28][20] ), .Z(n820) );
  ND3 U568 ( .A(n1024), .B(n1025), .C(n1026), .Z(\CARRYB[7][15] ) );
  ND3 U569 ( .A(n953), .B(n954), .C(n955), .Z(\CARRYB[12][12] ) );
  ND2 U570 ( .A(\SUMB[12][12] ), .B(\CARRYB[12][11] ), .Z(n956) );
  ND2 U571 ( .A(\CARRYB[41][28] ), .B(\ab[42][28] ), .Z(n1444) );
  ND2 U572 ( .A(\CARRYB[39][17] ), .B(\ab[40][17] ), .Z(n1378) );
  ND2 U573 ( .A(\CARRYB[45][4] ), .B(n302), .Z(n1639) );
  ND2 U574 ( .A(n2304), .B(\CARRYB[30][4] ), .Z(n2100) );
  ND2 U575 ( .A(\SUMB[41][5] ), .B(n384), .Z(n1816) );
  ND2 U576 ( .A(n2201), .B(\CARRYB[44][1] ), .Z(n2148) );
  ND2 U577 ( .A(\CARRYB[35][2] ), .B(\SUMB[35][3] ), .Z(n2016) );
  EO U578 ( .A(\SUMB[1][45] ), .B(n1456), .Z(\SUMB[2][44] ) );
  ND3 U579 ( .A(n1566), .B(n1567), .C(n1568), .Z(\CARRYB[2][34] ) );
  EO U580 ( .A(n2172), .B(n2188), .Z(\SUMB[1][35] ) );
  ND3 U581 ( .A(n1110), .B(n1111), .C(n1112), .Z(\CARRYB[4][32] ) );
  ND2 U582 ( .A(\CARRYB[3][32] ), .B(n358), .Z(n1111) );
  ND2 U583 ( .A(\CARRYB[3][32] ), .B(\SUMB[3][33] ), .Z(n1110) );
  EO U584 ( .A(n2184), .B(n2178), .Z(\SUMB[1][34] ) );
  ND3 U585 ( .A(n1056), .B(n1057), .C(n1058), .Z(\CARRYB[7][31] ) );
  ND2 U586 ( .A(\SUMB[6][32] ), .B(\CARRYB[6][31] ), .Z(n1056) );
  ND2 U587 ( .A(\SUMB[6][32] ), .B(n469), .Z(n1057) );
  ND2 U588 ( .A(\SUMB[7][32] ), .B(n514), .Z(n1061) );
  ND2 U589 ( .A(\CARRYB[11][45] ), .B(\ab[45][12] ), .Z(n2043) );
  ND2 U590 ( .A(\CARRYB[11][45] ), .B(\SUMB[11][46] ), .Z(n2042) );
  ND2 U591 ( .A(n2281), .B(\SUMB[3][31] ), .Z(n2067) );
  ND3 U592 ( .A(n906), .B(n907), .C(n908), .Z(\CARRYB[11][37] ) );
  ND2 U593 ( .A(\ab[41][15] ), .B(\SUMB[14][42] ), .Z(n1968) );
  ND2 U594 ( .A(\CARRYB[14][41] ), .B(\SUMB[14][42] ), .Z(n1969) );
  EO U595 ( .A(n332), .B(n2185), .Z(\SUMB[1][31] ) );
  ND3 U596 ( .A(n924), .B(n925), .C(n926), .Z(\CARRYB[10][30] ) );
  ND3 U597 ( .A(n1333), .B(n1334), .C(n1335), .Z(\CARRYB[2][28] ) );
  EO U598 ( .A(n2170), .B(n2167), .Z(\SUMB[1][30] ) );
  ND2 U599 ( .A(\SUMB[6][29] ), .B(n471), .Z(n1655) );
  ND3 U600 ( .A(n2036), .B(n2037), .C(n2038), .Z(\CARRYB[6][29] ) );
  ND3 U601 ( .A(n2011), .B(n2012), .C(n2013), .Z(\CARRYB[10][27] ) );
  EO U602 ( .A(\ab[41][15] ), .B(\CARRYB[14][41] ), .Z(n1963) );
  ND2 U603 ( .A(\CARRYB[19][43] ), .B(\SUMB[19][44] ), .Z(n1952) );
  EO U604 ( .A(n2174), .B(n2166), .Z(\SUMB[1][27] ) );
  ND3 U605 ( .A(n1464), .B(n1465), .C(n1466), .Z(\CARRYB[13][26] ) );
  ND2 U606 ( .A(\SUMB[12][27] ), .B(\CARRYB[12][26] ), .Z(n1464) );
  ND2 U607 ( .A(\CARRYB[12][26] ), .B(n680), .Z(n1466) );
  EO U608 ( .A(\CARRYB[15][31] ), .B(n1412), .Z(\SUMB[16][31] ) );
  EO U609 ( .A(\SUMB[15][32] ), .B(\ab[31][16] ), .Z(n1412) );
  ND3 U610 ( .A(n1438), .B(n1439), .C(n1440), .Z(\CARRYB[18][38] ) );
  EO U611 ( .A(\SUMB[19][44] ), .B(\ab[43][20] ), .Z(n1951) );
  ND3 U612 ( .A(n1605), .B(n1606), .C(n1607), .Z(\CARRYB[5][27] ) );
  ND2 U613 ( .A(\CARRYB[4][27] ), .B(\SUMB[4][28] ), .Z(n1605) );
  IVP U614 ( .A(n1660), .Z(n1283) );
  EO U615 ( .A(\CARRYB[9][26] ), .B(n604), .Z(n1582) );
  EO U616 ( .A(\CARRYB[13][30] ), .B(n705), .Z(n983) );
  ND3 U617 ( .A(n1099), .B(n1100), .C(n1101), .Z(\CARRYB[17][37] ) );
  ND2 U618 ( .A(\ab[37][17] ), .B(\SUMB[16][38] ), .Z(n1100) );
  EO U619 ( .A(\CARRYB[18][26] ), .B(n1379), .Z(\SUMB[19][26] ) );
  EO U620 ( .A(\SUMB[18][27] ), .B(\ab[26][19] ), .Z(n1379) );
  EO U621 ( .A(\CARRYB[13][24] ), .B(n703), .Z(n1286) );
  ND2 U622 ( .A(\ab[25][21] ), .B(\SUMB[20][26] ), .Z(n1552) );
  ND3 U623 ( .A(n1406), .B(n1407), .C(n1408), .Z(\CARRYB[22][28] ) );
  ND2 U624 ( .A(\SUMB[21][29] ), .B(\CARRYB[21][28] ), .Z(n1406) );
  ND2 U625 ( .A(\SUMB[21][29] ), .B(\ab[28][22] ), .Z(n1407) );
  EO U626 ( .A(\SUMB[22][24] ), .B(n1281), .Z(\SUMB[23][23] ) );
  ND3 U627 ( .A(n1989), .B(n1990), .C(n1991), .Z(\CARRYB[23][25] ) );
  EO U628 ( .A(\SUMB[1][23] ), .B(n1749), .Z(\SUMB[2][22] ) );
  EO U629 ( .A(n2316), .B(n2179), .Z(\SUMB[1][21] ) );
  ND3 U630 ( .A(n1263), .B(n1264), .C(n1265), .Z(\CARRYB[6][21] ) );
  EO U631 ( .A(\CARRYB[5][21] ), .B(n434), .Z(n1262) );
  ND3 U632 ( .A(n1016), .B(n1017), .C(n1018), .Z(\CARRYB[25][24] ) );
  ND2 U633 ( .A(\CARRYB[24][24] ), .B(\SUMB[24][25] ), .Z(n1016) );
  ND2 U634 ( .A(\CARRYB[24][24] ), .B(\ab[25][24] ), .Z(n1017) );
  EO U635 ( .A(\CARRYB[24][24] ), .B(n1015), .Z(\SUMB[25][24] ) );
  EO U636 ( .A(\SUMB[24][25] ), .B(\ab[25][24] ), .Z(n1015) );
  ND3 U637 ( .A(n878), .B(n879), .C(n880), .Z(\CARRYB[24][27] ) );
  EO U638 ( .A(\SUMB[23][29] ), .B(n1250), .Z(\SUMB[24][28] ) );
  ND3 U639 ( .A(n950), .B(n951), .C(n952), .Z(\CARRYB[27][33] ) );
  EO U640 ( .A(\CARRYB[27][37] ), .B(n1832), .Z(\SUMB[28][37] ) );
  EO U641 ( .A(\SUMB[27][38] ), .B(\ab[37][28] ), .Z(n1832) );
  ND3 U642 ( .A(n1833), .B(n1834), .C(n1835), .Z(\CARRYB[28][37] ) );
  ND3 U643 ( .A(n1840), .B(n1841), .C(n1842), .Z(\CARRYB[29][38] ) );
  EO U644 ( .A(\CARRYB[5][20] ), .B(n429), .Z(n1753) );
  ND3 U645 ( .A(n1804), .B(n1805), .C(n1806), .Z(\CARRYB[6][18] ) );
  ND3 U646 ( .A(n1828), .B(n1829), .C(n1830), .Z(\CARRYB[12][19] ) );
  ND2 U647 ( .A(\SUMB[11][20] ), .B(\CARRYB[11][19] ), .Z(n1828) );
  EO U648 ( .A(\SUMB[11][20] ), .B(n1827), .Z(\SUMB[12][19] ) );
  EO U649 ( .A(\CARRYB[11][19] ), .B(n658), .Z(n1827) );
  ND2 U650 ( .A(\CARRYB[28][19] ), .B(\ab[29][19] ), .Z(n821) );
  ND2 U651 ( .A(\SUMB[26][29] ), .B(\ab[28][27] ), .Z(n1702) );
  EO U652 ( .A(\SUMB[28][35] ), .B(n1154), .Z(\SUMB[29][34] ) );
  EO U653 ( .A(\CARRYB[3][15] ), .B(n367), .Z(n1792) );
  ND3 U654 ( .A(n1793), .B(n1794), .C(n1795), .Z(\CARRYB[4][15] ) );
  EO U655 ( .A(\SUMB[4][17] ), .B(n1774), .Z(\SUMB[5][16] ) );
  EO U656 ( .A(\CARRYB[4][16] ), .B(n400), .Z(n1774) );
  ND3 U657 ( .A(n1643), .B(n1644), .C(n1645), .Z(\CARRYB[6][15] ) );
  ND2 U658 ( .A(\SUMB[5][16] ), .B(n449), .Z(n1644) );
  ND2 U659 ( .A(\SUMB[5][16] ), .B(\CARRYB[5][15] ), .Z(n1643) );
  ND2 U660 ( .A(\CARRYB[5][15] ), .B(n449), .Z(n1645) );
  EO U661 ( .A(\CARRYB[4][17] ), .B(n966), .Z(\SUMB[5][17] ) );
  EO U662 ( .A(\SUMB[4][18] ), .B(n398), .Z(n966) );
  EO U663 ( .A(\CARRYB[5][18] ), .B(n1803), .Z(\SUMB[6][18] ) );
  ND3 U664 ( .A(n1471), .B(n1472), .C(n1473), .Z(\CARRYB[10][17] ) );
  ND2 U665 ( .A(\CARRYB[28][22] ), .B(\ab[29][22] ), .Z(n1647) );
  ND2 U666 ( .A(\CARRYB[28][22] ), .B(\SUMB[28][23] ), .Z(n1646) );
  ND3 U667 ( .A(n1476), .B(n1477), .C(n1478), .Z(\CARRYB[28][26] ) );
  EO U668 ( .A(\SUMB[28][31] ), .B(n1682), .Z(\SUMB[29][30] ) );
  EO U669 ( .A(\CARRYB[28][30] ), .B(\ab[30][29] ), .Z(n1682) );
  ND3 U670 ( .A(n1683), .B(n1684), .C(n1685), .Z(\CARRYB[29][30] ) );
  ND3 U671 ( .A(n1975), .B(n1976), .C(n1977), .Z(\CARRYB[2][13] ) );
  ND2 U672 ( .A(\CARRYB[1][13] ), .B(\SUMB[1][14] ), .Z(n1976) );
  ND2 U673 ( .A(n2266), .B(\SUMB[1][14] ), .Z(n1977) );
  ND3 U674 ( .A(n808), .B(n809), .C(n810), .Z(\CARRYB[16][17] ) );
  ND3 U675 ( .A(n1231), .B(n1232), .C(n1233), .Z(\CARRYB[31][19] ) );
  EO U676 ( .A(n576), .B(n2054), .Z(n2089) );
  EO U677 ( .A(\SUMB[8][16] ), .B(n1633), .Z(\SUMB[9][15] ) );
  EO U678 ( .A(\SUMB[13][14] ), .B(n675), .Z(n1693) );
  EN U679 ( .A(\SUMB[13][14] ), .B(n675), .Z(n1664) );
  ND3 U680 ( .A(n1824), .B(n1825), .C(n1826), .Z(\CARRYB[14][15] ) );
  ND3 U681 ( .A(n1786), .B(n1787), .C(n1788), .Z(\CARRYB[26][15] ) );
  ND2 U682 ( .A(n715), .B(\SUMB[25][16] ), .Z(n1787) );
  ND2 U683 ( .A(\CARRYB[33][25] ), .B(\SUMB[33][26] ), .Z(n1479) );
  ND3 U684 ( .A(n1387), .B(n1388), .C(n1389), .Z(\CARRYB[23][14] ) );
  ND2 U685 ( .A(\CARRYB[22][14] ), .B(n693), .Z(n1388) );
  EO U686 ( .A(n2183), .B(n2180), .Z(\SUMB[1][11] ) );
  ND3 U687 ( .A(n1008), .B(n1009), .C(n1010), .Z(\CARRYB[13][12] ) );
  ND2 U688 ( .A(\CARRYB[12][12] ), .B(n654), .Z(n1009) );
  ND2 U689 ( .A(\SUMB[12][12] ), .B(n635), .Z(n957) );
  EO U690 ( .A(\SUMB[34][15] ), .B(n1258), .Z(\SUMB[35][14] ) );
  ND3 U691 ( .A(n1847), .B(n1848), .C(n1849), .Z(\CARRYB[37][33] ) );
  ND2 U692 ( .A(\CARRYB[36][33] ), .B(\SUMB[36][34] ), .Z(n1847) );
  EO U693 ( .A(\SUMB[17][11] ), .B(n1561), .Z(\SUMB[18][10] ) );
  ND3 U694 ( .A(n1267), .B(n1268), .C(n1269), .Z(\CARRYB[19][10] ) );
  ND3 U695 ( .A(n1708), .B(n1709), .C(n1710), .Z(\CARRYB[24][10] ) );
  ND3 U696 ( .A(n2111), .B(n2112), .C(n2113), .Z(\CARRYB[12][9] ) );
  ND3 U697 ( .A(n1591), .B(n1592), .C(n1593), .Z(\CARRYB[33][11] ) );
  ND2 U698 ( .A(\SUMB[20][12] ), .B(n619), .Z(n1679) );
  ND3 U699 ( .A(n1148), .B(n1149), .C(n1150), .Z(\CARRYB[38][12] ) );
  EO U700 ( .A(\CARRYB[37][22] ), .B(\ab[38][22] ), .Z(n838) );
  EO U701 ( .A(\SUMB[36][28] ), .B(n1037), .Z(\SUMB[37][27] ) );
  EO U702 ( .A(\CARRYB[36][27] ), .B(\ab[37][27] ), .Z(n1037) );
  EO U703 ( .A(\CARRYB[13][8] ), .B(n2093), .Z(\SUMB[14][8] ) );
  EO U704 ( .A(\SUMB[13][9] ), .B(n536), .Z(n2093) );
  ND3 U705 ( .A(n1340), .B(n1341), .C(n1342), .Z(\CARRYB[38][8] ) );
  ND2 U706 ( .A(n531), .B(\SUMB[37][9] ), .Z(n1341) );
  ND3 U707 ( .A(n1875), .B(n1876), .C(n1877), .Z(\CARRYB[23][8] ) );
  ND2 U708 ( .A(\SUMB[22][9] ), .B(n533), .Z(n1876) );
  ND2 U709 ( .A(\SUMB[22][9] ), .B(\CARRYB[22][8] ), .Z(n1875) );
  ND2 U710 ( .A(\CARRYB[23][8] ), .B(\SUMB[23][9] ), .Z(n1918) );
  EO U711 ( .A(\CARRYB[23][10] ), .B(n597), .Z(n1707) );
  EN U712 ( .A(\CARRYB[23][10] ), .B(n597), .Z(n772) );
  ND3 U713 ( .A(n1733), .B(n1734), .C(n1735), .Z(\CARRYB[26][8] ) );
  EO U714 ( .A(\CARRYB[33][10] ), .B(n590), .Z(n1390) );
  ND3 U715 ( .A(n1626), .B(n1627), .C(n1628), .Z(\CARRYB[39][18] ) );
  ND3 U716 ( .A(n1854), .B(n1855), .C(n1856), .Z(\CARRYB[41][36] ) );
  ND2 U717 ( .A(\CARRYB[40][36] ), .B(\SUMB[40][37] ), .Z(n1854) );
  EO U718 ( .A(\CARRYB[40][36] ), .B(n1853), .Z(\SUMB[41][36] ) );
  EO U719 ( .A(\SUMB[40][37] ), .B(\ab[41][36] ), .Z(n1853) );
  ND3 U720 ( .A(n1941), .B(n1942), .C(n1943), .Z(\CARRYB[2][7] ) );
  ND2 U721 ( .A(n338), .B(\SUMB[1][8] ), .Z(n1942) );
  ND2 U722 ( .A(\CARRYB[1][7] ), .B(\SUMB[1][8] ), .Z(n1943) );
  ND3 U723 ( .A(n1972), .B(n1973), .C(n1974), .Z(\CARRYB[14][6] ) );
  EO U724 ( .A(n327), .B(n2244), .Z(\SUMB[1][7] ) );
  ND3 U725 ( .A(n1920), .B(n1921), .C(n1922), .Z(\CARRYB[19][7] ) );
  ND2 U726 ( .A(\SUMB[18][8] ), .B(n497), .Z(n1922) );
  ND2 U727 ( .A(\CARRYB[18][7] ), .B(\SUMB[18][8] ), .Z(n1920) );
  EO U728 ( .A(n1912), .B(\SUMB[23][9] ), .Z(\SUMB[24][8] ) );
  EO U729 ( .A(n534), .B(\CARRYB[23][8] ), .Z(n1912) );
  EO U730 ( .A(\CARRYB[22][8] ), .B(n533), .Z(n1874) );
  EO U731 ( .A(\CARRYB[42][9] ), .B(n586), .Z(n1724) );
  EO U732 ( .A(\SUMB[42][30] ), .B(n1448), .Z(\SUMB[43][29] ) );
  EO U733 ( .A(\CARRYB[42][29] ), .B(\ab[43][29] ), .Z(n1448) );
  ND3 U734 ( .A(n998), .B(n999), .C(n1000), .Z(\CARRYB[42][21] ) );
  EO U735 ( .A(\CARRYB[13][6] ), .B(n1971), .Z(\SUMB[14][6] ) );
  EO U736 ( .A(\SUMB[13][7] ), .B(n452), .Z(n1971) );
  ND3 U737 ( .A(n1934), .B(n1935), .C(n1936), .Z(\CARRYB[22][5] ) );
  ND2 U738 ( .A(n380), .B(\SUMB[21][6] ), .Z(n1935) );
  ND3 U739 ( .A(n1999), .B(n2000), .C(n2001), .Z(\CARRYB[26][7] ) );
  EO U740 ( .A(\SUMB[30][8] ), .B(n1365), .Z(\SUMB[31][7] ) );
  EO U741 ( .A(\CARRYB[30][7] ), .B(n469), .Z(n1365) );
  ND3 U742 ( .A(n2122), .B(n2123), .C(n2124), .Z(\CARRYB[35][5] ) );
  ND3 U743 ( .A(n1923), .B(n1924), .C(n1925), .Z(\CARRYB[42][16] ) );
  ND3 U744 ( .A(n1359), .B(n1360), .C(n1361), .Z(\CARRYB[42][25] ) );
  EO U745 ( .A(\CARRYB[4][6] ), .B(n2160), .Z(\SUMB[5][6] ) );
  EO U746 ( .A(\SUMB[4][7] ), .B(n448), .Z(n2160) );
  ND2 U747 ( .A(\SUMB[38][6] ), .B(n396), .Z(n940) );
  EO U748 ( .A(n285), .B(n2219), .Z(\SUMB[1][5] ) );
  EO U749 ( .A(n1930), .B(\SUMB[21][6] ), .Z(\SUMB[22][5] ) );
  EO U750 ( .A(n380), .B(\CARRYB[21][5] ), .Z(n1930) );
  EO U751 ( .A(\CARRYB[43][12] ), .B(\ab[44][12] ), .Z(n787) );
  ND2 U752 ( .A(\CARRYB[45][14] ), .B(\ab[46][14] ), .Z(n928) );
  ND2 U753 ( .A(\CARRYB[45][14] ), .B(\SUMB[45][15] ), .Z(n927) );
  IVP U754 ( .A(n2324), .Z(n2320) );
  ND2 U755 ( .A(\SUMB[45][5] ), .B(n302), .Z(n1638) );
  ND2 U756 ( .A(n358), .B(\CARRYB[31][4] ), .Z(n2105) );
  ND2 U757 ( .A(\CARRYB[30][3] ), .B(\SUMB[30][4] ), .Z(n2020) );
  ND3 U758 ( .A(n2060), .B(n2061), .C(n2062), .Z(\CARRYB[37][3] ) );
  EO U759 ( .A(\SUMB[45][25] ), .B(n1959), .Z(\SUMB[46][24] ) );
  EO U760 ( .A(\CARRYB[45][24] ), .B(\ab[46][24] ), .Z(n1959) );
  EO U761 ( .A(\SUMB[45][16] ), .B(n1139), .Z(\SUMB[46][15] ) );
  ND3 U762 ( .A(n927), .B(n928), .C(n929), .Z(\CARRYB[46][14] ) );
  EO U763 ( .A(\SUMB[45][19] ), .B(n1425), .Z(\SUMB[46][18] ) );
  EO U764 ( .A(\CARRYB[45][18] ), .B(\ab[46][18] ), .Z(n1425) );
  ND3 U765 ( .A(n1140), .B(n1141), .C(n1142), .Z(\CARRYB[46][15] ) );
  EO U766 ( .A(n1944), .B(\CARRYB[45][16] ), .Z(\SUMB[46][16] ) );
  EO U767 ( .A(\SUMB[45][33] ), .B(\ab[46][32] ), .Z(n1984) );
  ND3 U768 ( .A(n1511), .B(n1512), .C(n1513), .Z(\CARRYB[46][29] ) );
  ND3 U769 ( .A(n1882), .B(n1883), .C(n1884), .Z(\CARRYB[47][25] ) );
  EO U770 ( .A(\CARRYB[47][14] ), .B(\SUMB[47][15] ), .Z(\A1[60] ) );
  ND3 U771 ( .A(n2136), .B(n2137), .C(n2138), .Z(\CARRYB[10][1] ) );
  ND3 U772 ( .A(n2140), .B(n2141), .C(n2142), .Z(\CARRYB[6][1] ) );
  ND2 U773 ( .A(n1063), .B(\CARRYB[34][0] ), .Z(n1861) );
  ND2 U774 ( .A(\CARRYB[34][0] ), .B(\SUMB[34][1] ), .Z(n1863) );
  ND3 U775 ( .A(n1895), .B(n1896), .C(n1897), .Z(\CARRYB[34][1] ) );
  ND2 U776 ( .A(\CARRYB[37][1] ), .B(\SUMB[37][2] ), .Z(n2046) );
  EO U777 ( .A(\CARRYB[9][1] ), .B(n2135), .Z(\SUMB[10][1] ) );
  EO U778 ( .A(\CARRYB[24][1] ), .B(n2049), .Z(\SUMB[25][1] ) );
  EO U779 ( .A(\CARRYB[37][1] ), .B(n2045), .Z(\SUMB[38][1] ) );
  EO U780 ( .A(\SUMB[37][2] ), .B(n2233), .Z(n2045) );
  IVDA U781 ( .A(\ab[20][20] ), .Y(n244), .Z(n245) );
  IVDA U782 ( .A(\ab[25][25] ), .Y(n246), .Z(n247) );
  IVDA U783 ( .A(\ab[4][4] ), .Y(n348), .Z(n349) );
  IVDA U784 ( .A(\ab[19][19] ), .Y(n249), .Z(n250) );
  IVDA U785 ( .A(\ab[5][5] ), .Y(n375), .Z(n376) );
  IVDA U786 ( .A(\ab[6][6] ), .Y(n425), .Z(n426) );
  IVDA U787 ( .A(\ab[36][36] ), .Y(n253), .Z(n254) );
  IVDA U788 ( .A(\ab[46][46] ), .Y(n255), .Z(n256) );
  IVDA U789 ( .A(n2040), .Y(n257), .Z(n1350) );
  IVP U790 ( .A(\ab[26][26] ), .Z(n2371) );
  IVDA U791 ( .A(\ab[18][18] ), .Y(n258), .Z(n259) );
  IVDA U792 ( .A(\ab[14][14] ), .Y(n260), .Z(n261) );
  IVDA U793 ( .A(\ab[45][45] ), .Y(n262), .Z(n263) );
  IVDA U794 ( .A(\ab[12][12] ), .Y(n264), .Z(n265) );
  IVDA U795 ( .A(\ab[24][24] ), .Y(n266), .Z(n267) );
  IVP U796 ( .A(\ab[28][28] ), .Z(n2377) );
  IVDA U797 ( .A(\ab[34][34] ), .Y(n734), .Z(n735) );
  AN2P U798 ( .A(A[16]), .B(A[0]), .Z(n269) );
  AN2P U799 ( .A(A[20]), .B(n2040), .Z(n270) );
  IVP U800 ( .A(\ab[33][33] ), .Z(n2395) );
  IVP U801 ( .A(\ab[38][38] ), .Z(n2407) );
  IVP U802 ( .A(\ab[37][37] ), .Z(n2403) );
  IVP U803 ( .A(\ab[31][31] ), .Z(n2388) );
  IVP U804 ( .A(\ab[30][30] ), .Z(n2385) );
  IVP U805 ( .A(\ab[27][27] ), .Z(n2374) );
  IVDA U806 ( .A(\ab[17][17] ), .Y(n727), .Z(n728) );
  IVDA U807 ( .A(\ab[40][40] ), .Y(n651), .Z(n652) );
  IVP U808 ( .A(\ab[39][39] ), .Z(n2410) );
  IVDA U809 ( .A(\ab[43][43] ), .Y(n736), .Z(n737) );
  IVDA U810 ( .A(\ab[42][42] ), .Y(n649), .Z(n650) );
  IVP U811 ( .A(\ab[32][32] ), .Z(n2391) );
  IVDA U812 ( .A(\ab[23][23] ), .Y(n277), .Z(n278) );
  IVDA U813 ( .A(\ab[44][44] ), .Y(n279), .Z(n280) );
  IVDA U814 ( .A(\ab[9][9] ), .Y(n553), .Z(n554) );
  IVDA U815 ( .A(\ab[13][13] ), .Y(n645), .Z(n646) );
  IVDA U816 ( .A(\ab[22][22] ), .Y(n731), .Z(n732) );
  AN2P U817 ( .A(A[14]), .B(n2320), .Z(n284) );
  AN2P U818 ( .A(\ab[6][6] ), .B(n243), .Z(n285) );
  AN2P U819 ( .A(A[14]), .B(n2117), .Z(n286) );
  AN2P U820 ( .A(A[12]), .B(n2320), .Z(n287) );
  IVDA U821 ( .A(\ab[10][10] ), .Y(n578), .Z(n579) );
  AN2P U822 ( .A(A[11]), .B(PRODUCT[0]), .Z(n289) );
  IVP U823 ( .A(\ab[29][29] ), .Z(n2381) );
  IVDA U824 ( .A(\ab[21][21] ), .Y(n729), .Z(n730) );
  IVP U825 ( .A(\ab[16][16] ), .Z(n2354) );
  IVDA U826 ( .A(\ab[35][35] ), .Y(n299), .Z(n300) );
  AN2P U827 ( .A(n347), .B(n2319), .Z(n301) );
  AN2P U828 ( .A(n256), .B(n349), .Z(n302) );
  AN2P U829 ( .A(n2331), .B(n2421), .Z(n303) );
  AN2P U830 ( .A(n428), .B(n2331), .Z(n304) );
  AN2P U831 ( .A(n2420), .B(n2331), .Z(n305) );
  AN2P U832 ( .A(n428), .B(n2419), .Z(n306) );
  AN2P U833 ( .A(n2398), .B(n554), .Z(n307) );
  AN2P U834 ( .A(A[16]), .B(n265), .Z(n312) );
  IVDAP U835 ( .A(\ab[41][41] ), .Z(n316) );
  AN2P U836 ( .A(A[37]), .B(n2322), .Z(n318) );
  AN2P U837 ( .A(A[16]), .B(n2320), .Z(n319) );
  AN2P U838 ( .A(A[37]), .B(n2117), .Z(n320) );
  IVDA U839 ( .A(\CARRYB[13][13] ), .Y(n321), .Z(n322) );
  AN2P U840 ( .A(A[4]), .B(n2319), .Z(n323) );
  AN2P U841 ( .A(A[15]), .B(n2320), .Z(n324) );
  AN2P U842 ( .A(A[4]), .B(A[0]), .Z(n326) );
  AN2P U843 ( .A(\ab[8][8] ), .B(A[0]), .Z(n327) );
  IVP U844 ( .A(\ab[11][11] ), .Z(n2344) );
  AN2P U845 ( .A(A[21]), .B(PRODUCT[0]), .Z(n331) );
  AN2P U846 ( .A(A[32]), .B(n243), .Z(n332) );
  AN2P U847 ( .A(\ab[15][15] ), .B(n2117), .Z(n333) );
  AN2P U848 ( .A(\ab[39][39] ), .B(PRODUCT[0]), .Z(n334) );
  AN2P U849 ( .A(A[11]), .B(n2320), .Z(n335) );
  AN2P U850 ( .A(A[8]), .B(n2319), .Z(n336) );
  AN2P U851 ( .A(n2353), .B(n2328), .Z(n337) );
  AN2P U852 ( .A(A[7]), .B(n2319), .Z(n338) );
  AN2P U853 ( .A(n2319), .B(n2421), .Z(n339) );
  AN2P U854 ( .A(A[15]), .B(n2328), .Z(n340) );
  AN2P U855 ( .A(n2347), .B(n2325), .Z(n341) );
  AN2P U856 ( .A(A[37]), .B(n2325), .Z(n342) );
  AN2P U857 ( .A(n426), .B(n2319), .Z(n343) );
  AN2P U858 ( .A(n349), .B(n2326), .Z(n344) );
  AN2P U859 ( .A(n579), .B(n2319), .Z(n345) );
  IVDA U860 ( .A(\ab[3][3] ), .Y(n346), .Z(n347) );
  AN2P U861 ( .A(n2336), .B(n2326), .Z(n350) );
  AN2P U862 ( .A(n2345), .B(n2326), .Z(n351) );
  AN2P U863 ( .A(n2335), .B(n2325), .Z(n352) );
  AN2P U864 ( .A(n278), .B(n349), .Z(n353) );
  AN2P U865 ( .A(n2343), .B(n2328), .Z(n354) );
  AN2P U866 ( .A(n2340), .B(n2325), .Z(n355) );
  AN2P U867 ( .A(n2365), .B(n349), .Z(n356) );
  AN2P U868 ( .A(n2334), .B(n2328), .Z(n357) );
  AN2P U869 ( .A(n2389), .B(n2330), .Z(n358) );
  AN2P U870 ( .A(n2352), .B(n349), .Z(n359) );
  AN2P U871 ( .A(A[45]), .B(n349), .Z(n360) );
  AN2P U872 ( .A(n2402), .B(n2330), .Z(n361) );
  AN2P U873 ( .A(A[26]), .B(n349), .Z(n362) );
  AN2P U874 ( .A(n2398), .B(n2330), .Z(n363) );
  AN2P U875 ( .A(n2369), .B(n349), .Z(n364) );
  AN2P U876 ( .A(n2368), .B(n349), .Z(n365) );
  AN2P U877 ( .A(n2363), .B(n349), .Z(n366) );
  AN2P U878 ( .A(n2349), .B(n349), .Z(n367) );
  AN2P U879 ( .A(n2327), .B(n2421), .Z(n368) );
  AN2P U880 ( .A(n428), .B(n2329), .Z(n369) );
  AN2P U881 ( .A(n2405), .B(n2330), .Z(n370) );
  AN2P U882 ( .A(n728), .B(n349), .Z(n371) );
  AN2P U883 ( .A(A[13]), .B(n2329), .Z(n372) );
  AN2P U884 ( .A(n2339), .B(n2329), .Z(n373) );
  AN2P U885 ( .A(n2398), .B(n2332), .Z(n374) );
  IVDA U886 ( .A(\ab[8][8] ), .Y(n377), .Z(n378) );
  AN2P U887 ( .A(n316), .B(n349), .Z(n379) );
  AN2P U888 ( .A(n2364), .B(n376), .Z(n380) );
  AN2P U889 ( .A(n2372), .B(n376), .Z(n381) );
  AN2P U890 ( .A(n2417), .B(n2329), .Z(n382) );
  AN2P U891 ( .A(n2409), .B(n349), .Z(n383) );
  AN2P U892 ( .A(n2414), .B(n349), .Z(n384) );
  AN2P U893 ( .A(n2348), .B(n2329), .Z(n385) );
  AN2P U894 ( .A(n2345), .B(n2329), .Z(n386) );
  AN2P U895 ( .A(n2338), .B(n2329), .Z(n387) );
  AN2P U896 ( .A(n2342), .B(n2329), .Z(n388) );
  AN2P U897 ( .A(n737), .B(n2329), .Z(n389) );
  AN2P U898 ( .A(n2331), .B(n2329), .Z(n390) );
  AN2P U899 ( .A(n378), .B(n2329), .Z(n391) );
  AN2P U900 ( .A(n2382), .B(n2332), .Z(n392) );
  AN2P U901 ( .A(n2333), .B(n2329), .Z(n393) );
  AN2P U902 ( .A(n263), .B(n2331), .Z(n394) );
  AN2P U903 ( .A(n2362), .B(n376), .Z(n395) );
  AN2P U904 ( .A(n2408), .B(n2332), .Z(n396) );
  AN2P U905 ( .A(n2401), .B(n2332), .Z(n397) );
  AN2P U906 ( .A(n2355), .B(n376), .Z(n398) );
  AN2P U907 ( .A(n2399), .B(n2332), .Z(n399) );
  AN2P U908 ( .A(n2352), .B(n376), .Z(n400) );
  AN2P U909 ( .A(n2392), .B(n2332), .Z(n401) );
  AN2P U910 ( .A(n2360), .B(n376), .Z(n402) );
  AN2P U911 ( .A(n2396), .B(n2332), .Z(n403) );
  AN2P U912 ( .A(n2369), .B(n376), .Z(n404) );
  AN2P U913 ( .A(n265), .B(n2331), .Z(n405) );
  AN2P U914 ( .A(n2329), .B(A[47]), .Z(n406) );
  AN2P U915 ( .A(n2389), .B(n2332), .Z(n407) );
  AN2P U916 ( .A(n2367), .B(n376), .Z(n408) );
  AN2P U917 ( .A(n2398), .B(n2334), .Z(n409) );
  AN2P U918 ( .A(n2370), .B(n376), .Z(n410) );
  AN2P U919 ( .A(n2379), .B(n2332), .Z(n411) );
  AN2P U920 ( .A(n2375), .B(n2332), .Z(n412) );
  AN2P U921 ( .A(n2404), .B(n2332), .Z(n413) );
  AN2P U922 ( .A(n2412), .B(n349), .Z(n414) );
  AN2P U923 ( .A(n2356), .B(n376), .Z(n415) );
  AN2P U924 ( .A(n2386), .B(n2332), .Z(n416) );
  AN2P U925 ( .A(n261), .B(n2331), .Z(n417) );
  AN2P U926 ( .A(n2341), .B(n2331), .Z(n418) );
  AN2P U927 ( .A(n2336), .B(n2331), .Z(n419) );
  AN2P U928 ( .A(n2358), .B(n376), .Z(n420) );
  AN2P U929 ( .A(n267), .B(n376), .Z(n421) );
  AN2P U930 ( .A(n2346), .B(n2331), .Z(n422) );
  AN2P U931 ( .A(n2350), .B(n2331), .Z(n423) );
  AN2P U932 ( .A(n2339), .B(n2331), .Z(n424) );
  IVDA U933 ( .A(\ab[7][7] ), .Y(n427), .Z(n428) );
  AN2P U934 ( .A(n2360), .B(n426), .Z(n429) );
  AN2P U935 ( .A(n2369), .B(n426), .Z(n430) );
  AN2P U936 ( .A(n2382), .B(n2334), .Z(n431) );
  AN2P U937 ( .A(n2411), .B(n2331), .Z(n432) );
  AN2P U938 ( .A(n2392), .B(n2334), .Z(n433) );
  AN2P U939 ( .A(n2362), .B(n426), .Z(n434) );
  AN2P U940 ( .A(n2389), .B(n2334), .Z(n435) );
  AN2P U941 ( .A(n2355), .B(n426), .Z(n436) );
  AN2P U942 ( .A(n2337), .B(n2331), .Z(n437) );
  AN2P U943 ( .A(n2366), .B(n426), .Z(n438) );
  AN2P U944 ( .A(n2416), .B(n2331), .Z(n439) );
  AN2P U945 ( .A(n2400), .B(n2334), .Z(n440) );
  AN2P U946 ( .A(n2364), .B(n426), .Z(n441) );
  AN2P U947 ( .A(n2372), .B(n426), .Z(n442) );
  AN2P U948 ( .A(n2399), .B(n2334), .Z(n443) );
  AN2P U949 ( .A(n316), .B(n2331), .Z(n444) );
  AN2P U950 ( .A(n2352), .B(n2333), .Z(n445) );
  AN2P U951 ( .A(n2415), .B(n2331), .Z(n446) );
  AN2P U952 ( .A(n2375), .B(n426), .Z(n447) );
  AN2P U953 ( .A(n2333), .B(n2331), .Z(n448) );
  AN2P U954 ( .A(n2350), .B(n2333), .Z(n449) );
  AN2P U955 ( .A(n2398), .B(n428), .Z(n450) );
  AN2P U956 ( .A(n2370), .B(n426), .Z(n451) );
  AN2P U957 ( .A(n261), .B(n2333), .Z(n452) );
  AN2P U958 ( .A(n280), .B(n2333), .Z(n453) );
  AN2P U959 ( .A(n2413), .B(n2331), .Z(n454) );
  AN2P U960 ( .A(n2378), .B(n2334), .Z(n455) );
  AN2P U961 ( .A(n2404), .B(n2334), .Z(n456) );
  AN2P U962 ( .A(n2419), .B(n2333), .Z(n457) );
  AN2P U963 ( .A(n2411), .B(n2334), .Z(n458) );
  AN2P U964 ( .A(n2396), .B(n2334), .Z(n459) );
  AN2P U965 ( .A(n2358), .B(n426), .Z(n460) );
  AN2P U966 ( .A(n2346), .B(n2333), .Z(n461) );
  AN2P U967 ( .A(n267), .B(n426), .Z(n462) );
  AN2P U968 ( .A(n2408), .B(n2334), .Z(n463) );
  AN2P U969 ( .A(n2356), .B(n426), .Z(n464) );
  AN2P U970 ( .A(n2386), .B(n2334), .Z(n465) );
  AN2P U971 ( .A(n265), .B(n2333), .Z(n466) );
  AN2P U972 ( .A(n2369), .B(n428), .Z(n467) );
  AN2P U973 ( .A(n2370), .B(n428), .Z(n468) );
  AN2P U974 ( .A(n2386), .B(A[7]), .Z(n469) );
  AN2P U975 ( .A(n2360), .B(n428), .Z(n470) );
  AN2P U976 ( .A(n2375), .B(n428), .Z(n471) );
  AN2P U977 ( .A(n2400), .B(n428), .Z(n472) );
  AN2P U978 ( .A(n2415), .B(n2333), .Z(n473) );
  AN2P U979 ( .A(n2415), .B(n428), .Z(n474) );
  AN2P U980 ( .A(n2350), .B(n2335), .Z(n475) );
  AN2P U981 ( .A(n2389), .B(n428), .Z(n476) );
  AN2P U982 ( .A(n2362), .B(n428), .Z(n477) );
  AN2P U983 ( .A(n2413), .B(n2333), .Z(n478) );
  AN2P U984 ( .A(n2352), .B(n2335), .Z(n479) );
  AN2P U985 ( .A(n2346), .B(n2335), .Z(n480) );
  AN2P U986 ( .A(n2396), .B(n2335), .Z(n481) );
  AN2P U987 ( .A(n428), .B(n2333), .Z(n482) );
  AN2P U988 ( .A(n2336), .B(n2333), .Z(n483) );
  AN2P U989 ( .A(n2337), .B(n2333), .Z(n484) );
  AN2P U990 ( .A(n2418), .B(n2333), .Z(n485) );
  AN2P U991 ( .A(n280), .B(n428), .Z(n486) );
  AN2P U992 ( .A(n2333), .B(n2421), .Z(n487) );
  AN2P U993 ( .A(n2355), .B(n2335), .Z(n488) );
  AN2P U994 ( .A(n2382), .B(n428), .Z(n489) );
  AN2P U995 ( .A(n2404), .B(A[7]), .Z(n490) );
  AN2P U996 ( .A(n2341), .B(n2333), .Z(n491) );
  AN2P U997 ( .A(n2411), .B(A[7]), .Z(n492) );
  AN2P U998 ( .A(n316), .B(n2333), .Z(n493) );
  AN2P U999 ( .A(n2418), .B(n428), .Z(n494) );
  AN2P U1000 ( .A(n2366), .B(n428), .Z(n495) );
  AN2P U1001 ( .A(n2339), .B(n2333), .Z(n496) );
  AN2P U1002 ( .A(n2358), .B(n428), .Z(n497) );
  AN2P U1003 ( .A(n2372), .B(n428), .Z(n498) );
  AN2P U1004 ( .A(n316), .B(A[7]), .Z(n499) );
  AN2P U1005 ( .A(n267), .B(n428), .Z(n500) );
  AN2P U1006 ( .A(n2399), .B(A[7]), .Z(n501) );
  AN2P U1007 ( .A(n2378), .B(n428), .Z(n502) );
  AN2P U1008 ( .A(n2336), .B(n2419), .Z(n503) );
  AN2P U1009 ( .A(n2341), .B(n2335), .Z(n504) );
  AN2P U1010 ( .A(n2413), .B(n428), .Z(n505) );
  AN2P U1011 ( .A(n2364), .B(n428), .Z(n506) );
  AN2P U1012 ( .A(n2398), .B(n378), .Z(n507) );
  AN2P U1013 ( .A(n265), .B(n2335), .Z(n508) );
  AN2P U1014 ( .A(n2337), .B(n2335), .Z(n509) );
  AN2P U1015 ( .A(n2392), .B(A[7]), .Z(n510) );
  AN2P U1016 ( .A(n2408), .B(A[7]), .Z(n511) );
  AN2P U1017 ( .A(n2356), .B(n428), .Z(n512) );
  AN2P U1018 ( .A(n261), .B(n2335), .Z(n513) );
  AN2P U1019 ( .A(n2386), .B(n378), .Z(n514) );
  AN2P U1020 ( .A(n2360), .B(n378), .Z(n515) );
  AN2P U1021 ( .A(n280), .B(n2336), .Z(n516) );
  AN2P U1022 ( .A(n2355), .B(n2336), .Z(n517) );
  AN2P U1023 ( .A(n2336), .B(n2335), .Z(n518) );
  AN2P U1024 ( .A(n2356), .B(n2336), .Z(n519) );
  AN2P U1025 ( .A(n2415), .B(n2336), .Z(n520) );
  AN2P U1026 ( .A(n2418), .B(n2336), .Z(n521) );
  AN2P U1027 ( .A(n2396), .B(n378), .Z(n522) );
  AN2P U1028 ( .A(n2370), .B(n378), .Z(n523) );
  AN2P U1029 ( .A(n2372), .B(n378), .Z(n524) );
  AN2P U1030 ( .A(n2352), .B(n2336), .Z(n525) );
  AN2P U1031 ( .A(n2362), .B(n378), .Z(n526) );
  AN2P U1032 ( .A(n2350), .B(n2336), .Z(n527) );
  AN2P U1033 ( .A(n2339), .B(n2335), .Z(n528) );
  AN2P U1034 ( .A(n2389), .B(n378), .Z(n529) );
  AN2P U1035 ( .A(n2375), .B(n378), .Z(n530) );
  AN2P U1036 ( .A(n2404), .B(n378), .Z(n531) );
  AN2P U1037 ( .A(n265), .B(n2336), .Z(n532) );
  AN2P U1038 ( .A(n2366), .B(n378), .Z(n533) );
  AN2P U1039 ( .A(n267), .B(n378), .Z(n534) );
  AN2P U1040 ( .A(n2360), .B(n2338), .Z(n535) );
  AN2P U1041 ( .A(n261), .B(n2336), .Z(n536) );
  AN2P U1042 ( .A(n2392), .B(n378), .Z(n537) );
  AN2P U1043 ( .A(n2369), .B(n378), .Z(n538) );
  AN2P U1044 ( .A(n2364), .B(n378), .Z(n539) );
  AN2P U1045 ( .A(n2358), .B(n378), .Z(n540) );
  AN2P U1046 ( .A(n2382), .B(n378), .Z(n541) );
  AN2P U1047 ( .A(n2341), .B(n2336), .Z(n542) );
  AN2P U1048 ( .A(n2399), .B(n378), .Z(n543) );
  AN2P U1049 ( .A(n2346), .B(n2336), .Z(n544) );
  AN2P U1050 ( .A(n2411), .B(n378), .Z(n545) );
  AN2P U1051 ( .A(n316), .B(n378), .Z(n546) );
  AN2P U1052 ( .A(n2408), .B(n378), .Z(n547) );
  AN2P U1053 ( .A(n2352), .B(n2337), .Z(n548) );
  AN2P U1054 ( .A(n2378), .B(n378), .Z(n549) );
  AN2P U1055 ( .A(n2413), .B(n378), .Z(n550) );
  AN2P U1056 ( .A(n2400), .B(n378), .Z(n551) );
  AN2P U1057 ( .A(n2337), .B(n2336), .Z(n552) );
  AN2P U1058 ( .A(n2396), .B(n554), .Z(n555) );
  AN2P U1059 ( .A(n2358), .B(n2338), .Z(n556) );
  AN2P U1060 ( .A(n2369), .B(n2338), .Z(n557) );
  AN2P U1061 ( .A(n2392), .B(n554), .Z(n558) );
  AN2P U1062 ( .A(n2350), .B(n2337), .Z(n559) );
  AN2P U1063 ( .A(n2356), .B(n2338), .Z(n560) );
  AN2P U1064 ( .A(n2362), .B(n2338), .Z(n561) );
  AN2P U1065 ( .A(n2387), .B(n554), .Z(n562) );
  AN2P U1066 ( .A(n2375), .B(n2338), .Z(n563) );
  AN2P U1067 ( .A(n2370), .B(n2338), .Z(n564) );
  AN2P U1068 ( .A(n2364), .B(n2338), .Z(n565) );
  AN2P U1069 ( .A(n265), .B(n2337), .Z(n566) );
  AN2P U1070 ( .A(n2399), .B(n554), .Z(n567) );
  AN2P U1071 ( .A(A[32]), .B(n554), .Z(n568) );
  AN2P U1072 ( .A(n2400), .B(n554), .Z(n569) );
  AN2P U1073 ( .A(n2408), .B(n554), .Z(n570) );
  AN2P U1074 ( .A(n267), .B(n2338), .Z(n571) );
  AN2P U1075 ( .A(n2346), .B(n2337), .Z(n572) );
  AN2P U1076 ( .A(A[27]), .B(n2338), .Z(n573) );
  AN2P U1077 ( .A(n2355), .B(n2338), .Z(n574) );
  AN2P U1078 ( .A(n2378), .B(n554), .Z(n575) );
  AN2P U1079 ( .A(n261), .B(n2337), .Z(n576) );
  AN2P U1080 ( .A(n2339), .B(n2336), .Z(n577) );
  AN2P U1081 ( .A(n2382), .B(n2340), .Z(n580) );
  AN2P U1082 ( .A(n2360), .B(n579), .Z(n581) );
  AN2P U1083 ( .A(n2398), .B(n2340), .Z(n582) );
  AN2P U1084 ( .A(n2413), .B(n2337), .Z(n583) );
  AN2P U1085 ( .A(n2366), .B(n2338), .Z(n584) );
  AN2P U1086 ( .A(n2386), .B(n2340), .Z(n585) );
  AN2P U1087 ( .A(n2337), .B(n2415), .Z(n586) );
  AN2P U1088 ( .A(n2339), .B(n2337), .Z(n587) );
  AN2P U1089 ( .A(n2350), .B(n579), .Z(n588) );
  AN2P U1090 ( .A(n2404), .B(n554), .Z(n589) );
  AN2P U1091 ( .A(n2396), .B(n2340), .Z(n590) );
  AN2P U1092 ( .A(n2369), .B(n579), .Z(n591) );
  AN2P U1093 ( .A(n2382), .B(n554), .Z(n592) );
  AN2P U1094 ( .A(n2411), .B(n554), .Z(n593) );
  AN2P U1095 ( .A(n2341), .B(n2337), .Z(n594) );
  AN2P U1096 ( .A(n261), .B(n2339), .Z(n595) );
  AN2P U1097 ( .A(n2346), .B(n2339), .Z(n596) );
  AN2P U1098 ( .A(n267), .B(n579), .Z(n597) );
  AN2P U1099 ( .A(A[32]), .B(n2340), .Z(n598) );
  AN2P U1100 ( .A(n2400), .B(n2340), .Z(n599) );
  AN2P U1101 ( .A(n2355), .B(n579), .Z(n600) );
  AN2P U1102 ( .A(n2399), .B(n2340), .Z(n601) );
  AN2P U1103 ( .A(n2356), .B(n579), .Z(n602) );
  AN2P U1104 ( .A(n2366), .B(n579), .Z(n603) );
  AN2P U1105 ( .A(n2370), .B(n579), .Z(n604) );
  AN2P U1106 ( .A(n2378), .B(n2340), .Z(n605) );
  AN2P U1107 ( .A(n2341), .B(n2339), .Z(n606) );
  AN2P U1108 ( .A(n2352), .B(n579), .Z(n607) );
  AN2P U1109 ( .A(n2358), .B(n579), .Z(n608) );
  AN2P U1110 ( .A(n2398), .B(n2343), .Z(n609) );
  AN2P U1111 ( .A(n2375), .B(n2340), .Z(n610) );
  AN2P U1112 ( .A(A[27]), .B(n2340), .Z(n611) );
  AN2P U1113 ( .A(n316), .B(n2337), .Z(n612) );
  AN2P U1114 ( .A(n2404), .B(n2340), .Z(n613) );
  AN2P U1115 ( .A(n2392), .B(n2340), .Z(n614) );
  AN2P U1116 ( .A(n265), .B(n2339), .Z(n615) );
  AN2P U1117 ( .A(n2362), .B(n579), .Z(n616) );
  AN2P U1118 ( .A(n2364), .B(n579), .Z(n617) );
  AN2P U1119 ( .A(n2358), .B(n2342), .Z(n618) );
  AN2P U1120 ( .A(n2362), .B(n2342), .Z(n619) );
  AN2P U1121 ( .A(A[27]), .B(n2343), .Z(n620) );
  AN2P U1122 ( .A(n267), .B(n2342), .Z(n621) );
  AN2P U1123 ( .A(A[32]), .B(n2343), .Z(n622) );
  AN2P U1124 ( .A(n2382), .B(n2343), .Z(n623) );
  AN2P U1125 ( .A(n2352), .B(n2342), .Z(n624) );
  AN2P U1126 ( .A(n261), .B(n2342), .Z(n625) );
  AN2P U1127 ( .A(n2350), .B(n2342), .Z(n626) );
  AN2P U1128 ( .A(n2360), .B(n2342), .Z(n627) );
  AN2P U1129 ( .A(n2375), .B(n2343), .Z(n628) );
  AN2P U1130 ( .A(n2355), .B(n2342), .Z(n629) );
  AN2P U1131 ( .A(n2370), .B(n2343), .Z(n630) );
  AN2P U1132 ( .A(n2387), .B(n2343), .Z(n631) );
  AN2P U1133 ( .A(n2396), .B(n2343), .Z(n632) );
  AN2P U1134 ( .A(n247), .B(n2343), .Z(n633) );
  AN2P U1135 ( .A(n2346), .B(n2342), .Z(n635) );
  AN2P U1136 ( .A(n2392), .B(n2343), .Z(n636) );
  AN2P U1137 ( .A(n2339), .B(n2411), .Z(n637) );
  AN2P U1138 ( .A(n2356), .B(n2342), .Z(n638) );
  AN2P U1139 ( .A(n2378), .B(n2343), .Z(n639) );
  AN2P U1140 ( .A(n2408), .B(n2339), .Z(n640) );
  AN2P U1141 ( .A(n2364), .B(n2342), .Z(n641) );
  AN2P U1142 ( .A(n2366), .B(n2342), .Z(n642) );
  AN2P U1143 ( .A(n2399), .B(n2343), .Z(n643) );
  AN2P U1144 ( .A(n265), .B(n2341), .Z(n644) );
  IVA U1145 ( .A(\ab[15][15] ), .Z(n2351) );
  AN2P U1146 ( .A(n2394), .B(n2345), .Z(n653) );
  AN2P U1147 ( .A(n646), .B(n265), .Z(n654) );
  AN2P U1148 ( .A(A[15]), .B(n265), .Z(n655) );
  AN2P U1149 ( .A(n2341), .B(n2400), .Z(n656) );
  AN2P U1150 ( .A(A[26]), .B(n2345), .Z(n657) );
  AN2P U1151 ( .A(n250), .B(n265), .Z(n658) );
  AN2P U1152 ( .A(n2348), .B(n265), .Z(n659) );
  AN2P U1153 ( .A(n267), .B(n2345), .Z(n660) );
  AN2P U1154 ( .A(A[25]), .B(n2345), .Z(n661) );
  AN2P U1155 ( .A(n2384), .B(n2345), .Z(n662) );
  AN2P U1156 ( .A(A[27]), .B(n2345), .Z(n663) );
  AN2P U1157 ( .A(n259), .B(n265), .Z(n664) );
  AN2P U1158 ( .A(n245), .B(n265), .Z(n665) );
  AN2P U1159 ( .A(n278), .B(n265), .Z(n666) );
  AN2P U1160 ( .A(n2363), .B(n265), .Z(n667) );
  AN2P U1161 ( .A(A[28]), .B(n2345), .Z(n668) );
  AN2P U1162 ( .A(n2390), .B(n2345), .Z(n669) );
  AN2P U1163 ( .A(n2345), .B(n300), .Z(n672) );
  AN2P U1164 ( .A(n2387), .B(n2345), .Z(n673) );
  AN2P U1165 ( .A(n2397), .B(n2345), .Z(n674) );
  AN2P U1166 ( .A(n2348), .B(n2346), .Z(n675) );
  AN2P U1167 ( .A(n2380), .B(n2345), .Z(n676) );
  AN2P U1168 ( .A(A[17]), .B(n265), .Z(n677) );
  AN2P U1169 ( .A(n2365), .B(n265), .Z(n678) );
  AN2P U1170 ( .A(n250), .B(n2346), .Z(n679) );
  AN2P U1171 ( .A(A[26]), .B(n646), .Z(n680) );
  AN2P U1172 ( .A(n2365), .B(n646), .Z(n681) );
  AN2P U1173 ( .A(A[27]), .B(n646), .Z(n682) );
  AN2P U1174 ( .A(A[25]), .B(n646), .Z(n683) );
  AN2P U1175 ( .A(n278), .B(n646), .Z(n684) );
  AN2P U1176 ( .A(n2387), .B(n646), .Z(n685) );
  AN2P U1177 ( .A(n2353), .B(n2346), .Z(n686) );
  AN2P U1178 ( .A(n728), .B(n2346), .Z(n687) );
  AN2P U1179 ( .A(n245), .B(n2346), .Z(n688) );
  AN2P U1180 ( .A(n2380), .B(n646), .Z(n689) );
  AN2P U1181 ( .A(n267), .B(n646), .Z(n690) );
  AN2P U1182 ( .A(A[15]), .B(n2346), .Z(n691) );
  AN2P U1183 ( .A(n2384), .B(n646), .Z(n692) );
  AN2P U1184 ( .A(n278), .B(n2348), .Z(n693) );
  AN2P U1185 ( .A(n646), .B(n2390), .Z(n694) );
  AN2P U1186 ( .A(n259), .B(n2346), .Z(n695) );
  AN2P U1187 ( .A(n2363), .B(n2346), .Z(n696) );
  AN2P U1188 ( .A(A[28]), .B(n646), .Z(n697) );
  AN2P U1189 ( .A(n259), .B(n2347), .Z(n698) );
  AN2P U1190 ( .A(n250), .B(n2347), .Z(n699) );
  AN2P U1191 ( .A(n2365), .B(n2348), .Z(n700) );
  AN2P U1192 ( .A(n2352), .B(n2347), .Z(n701) );
  AN2P U1193 ( .A(n2380), .B(n2348), .Z(n702) );
  AN2P U1194 ( .A(n267), .B(n2348), .Z(n703) );
  AN2P U1195 ( .A(n2363), .B(n2348), .Z(n704) );
  AN2P U1196 ( .A(n2348), .B(n2384), .Z(n705) );
  AN2P U1197 ( .A(n2376), .B(n2348), .Z(n706) );
  AN2P U1198 ( .A(n2350), .B(n2347), .Z(n707) );
  AN2P U1199 ( .A(A[26]), .B(n2348), .Z(n708) );
  AN2P U1200 ( .A(n245), .B(n2347), .Z(n709) );
  AN2P U1201 ( .A(n728), .B(n2347), .Z(n710) );
  AN2P U1202 ( .A(n247), .B(n2348), .Z(n711) );
  AN2P U1203 ( .A(n2373), .B(n2348), .Z(n712) );
  AN2P U1204 ( .A(n259), .B(n2350), .Z(n713) );
  AN2P U1205 ( .A(n2350), .B(n2380), .Z(n714) );
  AN2P U1206 ( .A(n2370), .B(n2350), .Z(n715) );
  AN2P U1207 ( .A(n278), .B(n2350), .Z(n716) );
  AN2P U1208 ( .A(n2355), .B(n2350), .Z(n717) );
  AN2P U1209 ( .A(n2372), .B(n2350), .Z(n718) );
  AN2P U1210 ( .A(n2363), .B(n2350), .Z(n719) );
  AN2P U1211 ( .A(n2365), .B(n2350), .Z(n720) );
  AN2P U1212 ( .A(n2375), .B(n2349), .Z(n721) );
  AN2P U1213 ( .A(n2352), .B(n2350), .Z(n722) );
  AN2P U1214 ( .A(n2369), .B(n2349), .Z(n723) );
  AN2P U1215 ( .A(n245), .B(n2350), .Z(n724) );
  AN2P U1216 ( .A(n250), .B(n2350), .Z(n725) );
  AN2P U1217 ( .A(n267), .B(n2349), .Z(n726) );
  EO U1218 ( .A(\ab[35][15] ), .B(\CARRYB[14][35] ), .Z(n738) );
  ND2 U1219 ( .A(\CARRYB[13][36] ), .B(\SUMB[13][37] ), .Z(n740) );
  ND2 U1220 ( .A(\ab[36][14] ), .B(\SUMB[13][37] ), .Z(n741) );
  ND3 U1221 ( .A(n739), .B(n740), .C(n741), .Z(\CARRYB[14][36] ) );
  ND2 U1222 ( .A(\ab[35][15] ), .B(\CARRYB[14][35] ), .Z(n742) );
  ND3P U1223 ( .A(n742), .B(n743), .C(n744), .Z(\CARRYB[15][35] ) );
  EO U1224 ( .A(\CARRYB[2][41] ), .B(n2286), .Z(n745) );
  EO U1225 ( .A(\SUMB[2][42] ), .B(n745), .Z(\SUMB[3][41] ) );
  ND2 U1226 ( .A(\SUMB[2][42] ), .B(\CARRYB[2][41] ), .Z(n746) );
  ND2 U1227 ( .A(\SUMB[2][42] ), .B(n2286), .Z(n747) );
  ND2 U1228 ( .A(\CARRYB[2][41] ), .B(n2286), .Z(n748) );
  ND3 U1229 ( .A(n746), .B(n747), .C(n748), .Z(\CARRYB[3][41] ) );
  ND2 U1230 ( .A(n1572), .B(n750), .Z(n751) );
  ND2P U1231 ( .A(n749), .B(\SUMB[40][20] ), .Z(n752) );
  ND2P U1232 ( .A(n751), .B(n752), .Z(\SUMB[41][19] ) );
  IVP U1233 ( .A(n1572), .Z(n749) );
  IVP U1234 ( .A(\SUMB[40][20] ), .Z(n750) );
  ND2P U1235 ( .A(\CARRYB[21][32] ), .B(\ab[32][22] ), .Z(n1400) );
  ND2P U1236 ( .A(\SUMB[21][33] ), .B(\CARRYB[21][32] ), .Z(n1398) );
  EOP U1237 ( .A(n1216), .B(\SUMB[25][7] ), .Z(\SUMB[26][6] ) );
  EO U1238 ( .A(n451), .B(\CARRYB[25][6] ), .Z(n1216) );
  EO U1239 ( .A(\SUMB[23][12] ), .B(n1322), .Z(\SUMB[24][11] ) );
  ND2 U1240 ( .A(\CARRYB[45][0] ), .B(\SUMB[45][1] ), .Z(n2131) );
  ND2P U1241 ( .A(\SUMB[43][9] ), .B(n516), .Z(n1291) );
  ND2P U1242 ( .A(\SUMB[43][9] ), .B(\CARRYB[43][8] ), .Z(n1290) );
  ND3 U1243 ( .A(n1576), .B(n1577), .C(n1578), .Z(\CARRYB[37][19] ) );
  ND3 U1244 ( .A(n934), .B(n935), .C(n936), .Z(\CARRYB[18][27] ) );
  EO3P U1245 ( .A(n657), .B(\CARRYB[25][12] ), .C(\SUMB[25][13] ), .Z(
        \SUMB[26][12] ) );
  EO U1246 ( .A(n620), .B(\CARRYB[26][11] ), .Z(n753) );
  ND2 U1247 ( .A(n657), .B(\CARRYB[25][12] ), .Z(n754) );
  ND2 U1248 ( .A(n657), .B(\SUMB[25][13] ), .Z(n755) );
  ND2 U1249 ( .A(\CARRYB[25][12] ), .B(\SUMB[25][13] ), .Z(n756) );
  ND2 U1250 ( .A(n620), .B(\CARRYB[26][11] ), .Z(n757) );
  ND2P U1251 ( .A(n620), .B(\SUMB[26][12] ), .Z(n758) );
  ND2P U1252 ( .A(\CARRYB[26][11] ), .B(\SUMB[26][12] ), .Z(n759) );
  ND3P U1253 ( .A(n757), .B(n758), .C(n759), .Z(\CARRYB[27][11] ) );
  ND2 U1254 ( .A(\ab[25][21] ), .B(\CARRYB[20][25] ), .Z(n1551) );
  EO U1255 ( .A(\ab[25][21] ), .B(\CARRYB[20][25] ), .Z(n1547) );
  EO U1256 ( .A(n1132), .B(\SUMB[12][29] ), .Z(\SUMB[13][28] ) );
  EOP U1257 ( .A(\SUMB[31][26] ), .B(n760), .Z(\SUMB[32][25] ) );
  ND2 U1258 ( .A(\SUMB[31][26] ), .B(\CARRYB[31][25] ), .Z(n761) );
  ND2 U1259 ( .A(\SUMB[31][26] ), .B(\ab[32][25] ), .Z(n762) );
  ND2 U1260 ( .A(\CARRYB[31][25] ), .B(\ab[32][25] ), .Z(n763) );
  ND3 U1261 ( .A(n823), .B(n824), .C(n825), .Z(n764) );
  ND3 U1262 ( .A(n823), .B(n824), .C(n825), .Z(\CARRYB[43][12] ) );
  ND3 U1263 ( .A(n1005), .B(n1006), .C(n1007), .Z(\CARRYB[32][26] ) );
  ND2 U1264 ( .A(n1474), .B(\CARRYB[45][4] ), .Z(n1637) );
  ND3 U1265 ( .A(n1151), .B(n1152), .C(n1153), .Z(n765) );
  EOP U1266 ( .A(\SUMB[45][6] ), .B(n305), .Z(n766) );
  EOP U1267 ( .A(n876), .B(n766), .Z(\SUMB[46][5] ) );
  EO U1268 ( .A(\CARRYB[16][24] ), .B(\ab[24][17] ), .Z(n767) );
  EO U1269 ( .A(\SUMB[16][25] ), .B(n767), .Z(\SUMB[17][24] ) );
  ND2 U1270 ( .A(\SUMB[16][25] ), .B(\CARRYB[16][24] ), .Z(n768) );
  ND2 U1271 ( .A(\SUMB[16][25] ), .B(\ab[24][17] ), .Z(n769) );
  ND2 U1272 ( .A(\CARRYB[16][24] ), .B(\ab[24][17] ), .Z(n770) );
  ND3 U1273 ( .A(n768), .B(n769), .C(n770), .Z(\CARRYB[17][24] ) );
  ND2P U1274 ( .A(n1489), .B(n1707), .Z(n1491) );
  ND3 U1275 ( .A(n1637), .B(n1638), .C(n1639), .Z(\CARRYB[46][4] ) );
  ND3 U1276 ( .A(n1678), .B(n1679), .C(n1680), .Z(\CARRYB[21][11] ) );
  EO3 U1277 ( .A(\SUMB[14][13] ), .B(n655), .C(\CARRYB[14][12] ), .Z(
        \SUMB[15][12] ) );
  IVP U1278 ( .A(n900), .Z(n901) );
  ND3 U1279 ( .A(n931), .B(n932), .C(n933), .Z(\CARRYB[35][20] ) );
  ND3 U1280 ( .A(n1347), .B(n1348), .C(n1349), .Z(n771) );
  ND3 U1281 ( .A(n1347), .B(n1348), .C(n1349), .Z(\CARRYB[40][11] ) );
  ND3 U1282 ( .A(n1092), .B(n1093), .C(n1094), .Z(\CARRYB[25][28] ) );
  EO3P U1283 ( .A(\CARRYB[41][20] ), .B(\ab[42][20] ), .C(\SUMB[41][21] ), .Z(
        \SUMB[42][20] ) );
  ND2 U1284 ( .A(\CARRYB[41][20] ), .B(\SUMB[41][21] ), .Z(n773) );
  ND2 U1285 ( .A(\CARRYB[41][20] ), .B(\ab[42][20] ), .Z(n774) );
  ND2 U1286 ( .A(\SUMB[41][21] ), .B(\ab[42][20] ), .Z(n775) );
  ND3P U1287 ( .A(n773), .B(n774), .C(n775), .Z(\CARRYB[42][20] ) );
  ND3 U1288 ( .A(n1623), .B(n1624), .C(n1625), .Z(\CARRYB[30][26] ) );
  EO3P U1289 ( .A(\SUMB[30][26] ), .B(\ab[31][25] ), .C(\CARRYB[30][25] ), .Z(
        \SUMB[31][25] ) );
  ND2 U1290 ( .A(\SUMB[30][26] ), .B(\CARRYB[30][25] ), .Z(n776) );
  ND2 U1291 ( .A(\SUMB[30][26] ), .B(\ab[31][25] ), .Z(n777) );
  ND2 U1292 ( .A(\CARRYB[30][25] ), .B(\ab[31][25] ), .Z(n778) );
  EO3 U1293 ( .A(\CARRYB[11][16] ), .B(n312), .C(\SUMB[11][17] ), .Z(
        \SUMB[12][16] ) );
  ND2 U1294 ( .A(\CARRYB[11][16] ), .B(\SUMB[11][17] ), .Z(n779) );
  ND2 U1295 ( .A(\CARRYB[11][16] ), .B(n312), .Z(n780) );
  ND2 U1296 ( .A(\SUMB[11][17] ), .B(n312), .Z(n781) );
  ND3 U1297 ( .A(n779), .B(n780), .C(n781), .Z(\CARRYB[12][16] ) );
  EO3 U1298 ( .A(\SUMB[29][11] ), .B(n580), .C(\CARRYB[29][10] ), .Z(n782) );
  EO3P U1299 ( .A(\CARRYB[36][11] ), .B(n656), .C(\SUMB[36][12] ), .Z(
        \SUMB[37][11] ) );
  ND2 U1300 ( .A(\CARRYB[36][11] ), .B(\SUMB[36][12] ), .Z(n783) );
  ND2 U1301 ( .A(\CARRYB[36][11] ), .B(n656), .Z(n784) );
  ND2 U1302 ( .A(\SUMB[36][12] ), .B(n656), .Z(n785) );
  ND3 U1303 ( .A(n783), .B(n784), .C(n785), .Z(\CARRYB[37][11] ) );
  ND3 U1304 ( .A(n1700), .B(n1701), .C(n1702), .Z(\CARRYB[27][28] ) );
  EOP U1305 ( .A(\SUMB[43][13] ), .B(n787), .Z(\SUMB[44][12] ) );
  ND2 U1306 ( .A(\SUMB[43][13] ), .B(n764), .Z(n788) );
  ND2 U1307 ( .A(\SUMB[43][13] ), .B(\ab[44][12] ), .Z(n789) );
  ND2 U1308 ( .A(n764), .B(\ab[44][12] ), .Z(n790) );
  ND3P U1309 ( .A(n788), .B(n789), .C(n790), .Z(\CARRYB[44][12] ) );
  EO3P U1310 ( .A(\SUMB[20][20] ), .B(\ab[21][19] ), .C(\CARRYB[20][19] ), .Z(
        \SUMB[21][19] ) );
  ND2 U1311 ( .A(\SUMB[20][20] ), .B(\CARRYB[20][19] ), .Z(n791) );
  ND2 U1312 ( .A(\SUMB[20][20] ), .B(\ab[21][19] ), .Z(n792) );
  ND2 U1313 ( .A(\CARRYB[20][19] ), .B(\ab[21][19] ), .Z(n793) );
  ND3 U1314 ( .A(n791), .B(n792), .C(n793), .Z(\CARRYB[21][19] ) );
  ND2 U1315 ( .A(\SUMB[6][29] ), .B(\CARRYB[6][28] ), .Z(n1654) );
  ND2P U1316 ( .A(\SUMB[34][25] ), .B(\CARRYB[34][24] ), .Z(n910) );
  EO U1317 ( .A(\SUMB[37][30] ), .B(n794), .Z(\SUMB[38][29] ) );
  ND2 U1318 ( .A(\SUMB[37][30] ), .B(\CARRYB[37][29] ), .Z(n795) );
  ND2 U1319 ( .A(\SUMB[37][30] ), .B(\ab[38][29] ), .Z(n796) );
  ND2 U1320 ( .A(\CARRYB[37][29] ), .B(\ab[38][29] ), .Z(n797) );
  ND3 U1321 ( .A(n795), .B(n796), .C(n797), .Z(\CARRYB[38][29] ) );
  ND2 U1322 ( .A(\SUMB[20][12] ), .B(\CARRYB[20][11] ), .Z(n1678) );
  AN2P U1323 ( .A(n2168), .B(n2190), .Z(\CARRYB[1][18] ) );
  ND3 U1324 ( .A(n1479), .B(n1480), .C(n1481), .Z(\CARRYB[34][25] ) );
  EOP U1325 ( .A(n2243), .B(n2237), .Z(\SUMB[1][44] ) );
  ND3 U1326 ( .A(n1278), .B(n1279), .C(n1280), .Z(\CARRYB[19][25] ) );
  IVA U1327 ( .A(\CARRYB[34][14] ), .Z(n798) );
  IVP U1328 ( .A(n798), .Z(n799) );
  ND2 U1329 ( .A(\SUMB[5][26] ), .B(\CARRYB[5][25] ), .Z(n1530) );
  EOP U1330 ( .A(\CARRYB[23][14] ), .B(n703), .Z(n800) );
  EOP U1331 ( .A(\SUMB[23][15] ), .B(n800), .Z(\SUMB[24][14] ) );
  ND2 U1332 ( .A(\SUMB[23][15] ), .B(\CARRYB[23][14] ), .Z(n801) );
  ND2 U1333 ( .A(\SUMB[23][15] ), .B(n703), .Z(n802) );
  ND2 U1334 ( .A(\CARRYB[23][14] ), .B(n703), .Z(n803) );
  ND3P U1335 ( .A(n801), .B(n802), .C(n803), .Z(\CARRYB[24][14] ) );
  ND3P U1336 ( .A(n1227), .B(n1228), .C(n1229), .Z(\CARRYB[41][11] ) );
  ND2 U1337 ( .A(\SUMB[38][6] ), .B(\CARRYB[38][5] ), .Z(n939) );
  EO3 U1338 ( .A(\CARRYB[38][26] ), .B(\ab[39][26] ), .C(\SUMB[38][27] ), .Z(
        \SUMB[39][26] ) );
  ND2 U1339 ( .A(\CARRYB[38][26] ), .B(\SUMB[38][27] ), .Z(n804) );
  ND2 U1340 ( .A(\CARRYB[38][26] ), .B(\ab[39][26] ), .Z(n805) );
  ND2 U1341 ( .A(\SUMB[38][27] ), .B(\ab[39][26] ), .Z(n806) );
  ND3 U1342 ( .A(n804), .B(n805), .C(n806), .Z(\CARRYB[39][26] ) );
  EO U1343 ( .A(\CARRYB[39][26] ), .B(\ab[40][26] ), .Z(n856) );
  EO U1344 ( .A(\CARRYB[42][11] ), .B(\ab[43][11] ), .Z(n807) );
  EO U1345 ( .A(\SUMB[42][12] ), .B(n807), .Z(\SUMB[43][11] ) );
  ND2 U1346 ( .A(\CARRYB[15][17] ), .B(\SUMB[15][18] ), .Z(n808) );
  ND2 U1347 ( .A(\CARRYB[15][17] ), .B(\ab[17][16] ), .Z(n809) );
  ND2 U1348 ( .A(\SUMB[15][18] ), .B(\ab[17][16] ), .Z(n810) );
  ND2P U1349 ( .A(\CARRYB[6][16] ), .B(n479), .Z(n1182) );
  ND2P U1350 ( .A(\SUMB[6][17] ), .B(\CARRYB[6][16] ), .Z(n1180) );
  ND2P U1351 ( .A(n1314), .B(\ab[34][25] ), .Z(n1480) );
  EOP U1352 ( .A(\CARRYB[12][20] ), .B(n688), .Z(n811) );
  EOP U1353 ( .A(\SUMB[12][21] ), .B(n811), .Z(\SUMB[13][20] ) );
  ND2 U1354 ( .A(\SUMB[12][21] ), .B(\CARRYB[12][20] ), .Z(n812) );
  ND2 U1355 ( .A(\SUMB[12][21] ), .B(n688), .Z(n813) );
  ND2 U1356 ( .A(\CARRYB[12][20] ), .B(n688), .Z(n814) );
  ND3 U1357 ( .A(n812), .B(n813), .C(n814), .Z(\CARRYB[13][20] ) );
  EOP U1358 ( .A(\CARRYB[21][31] ), .B(\ab[31][22] ), .Z(n815) );
  EOP U1359 ( .A(\SUMB[21][32] ), .B(n815), .Z(\SUMB[22][31] ) );
  ND2 U1360 ( .A(\SUMB[21][32] ), .B(\CARRYB[21][31] ), .Z(n816) );
  ND2 U1361 ( .A(\SUMB[21][32] ), .B(\ab[31][22] ), .Z(n817) );
  ND2 U1362 ( .A(\CARRYB[21][31] ), .B(\ab[31][22] ), .Z(n818) );
  ND3 U1363 ( .A(n816), .B(n817), .C(n818), .Z(\CARRYB[22][31] ) );
  ND2 U1364 ( .A(\SUMB[43][19] ), .B(\CARRYB[43][18] ), .Z(n1630) );
  ND2 U1365 ( .A(\CARRYB[43][18] ), .B(\ab[44][18] ), .Z(n1632) );
  ND2 U1366 ( .A(\SUMB[28][20] ), .B(\ab[29][19] ), .Z(n822) );
  EO3 U1367 ( .A(\SUMB[42][13] ), .B(\ab[43][12] ), .C(\CARRYB[42][12] ), .Z(
        \SUMB[43][12] ) );
  ND2 U1368 ( .A(\SUMB[42][13] ), .B(\CARRYB[42][12] ), .Z(n823) );
  ND2 U1369 ( .A(\SUMB[42][13] ), .B(\ab[43][12] ), .Z(n824) );
  ND2 U1370 ( .A(\CARRYB[42][12] ), .B(\ab[43][12] ), .Z(n825) );
  EO3P U1371 ( .A(\SUMB[10][20] ), .B(n618), .C(\CARRYB[10][19] ), .Z(
        \SUMB[11][19] ) );
  ND2P U1372 ( .A(\SUMB[10][20] ), .B(n618), .Z(n827) );
  ND3P U1373 ( .A(n826), .B(n827), .C(n828), .Z(\CARRYB[11][19] ) );
  EOP U1374 ( .A(\SUMB[20][16] ), .B(n719), .Z(n829) );
  ENP U1375 ( .A(n830), .B(n2248), .Z(n1456) );
  ND2 U1376 ( .A(n2237), .B(n2243), .Z(n830) );
  EO3P U1377 ( .A(\SUMB[21][14] ), .B(n681), .C(\CARRYB[21][13] ), .Z(
        \SUMB[22][13] ) );
  ND2 U1378 ( .A(\SUMB[21][14] ), .B(\CARRYB[21][13] ), .Z(n831) );
  ND2 U1379 ( .A(\SUMB[21][14] ), .B(n681), .Z(n832) );
  ND2 U1380 ( .A(\CARRYB[21][13] ), .B(n681), .Z(n833) );
  ND3 U1381 ( .A(n831), .B(n832), .C(n833), .Z(\CARRYB[22][13] ) );
  EO3 U1382 ( .A(\SUMB[15][33] ), .B(\ab[32][16] ), .C(\CARRYB[15][32] ), .Z(
        \SUMB[16][32] ) );
  ND2 U1383 ( .A(\CARRYB[15][32] ), .B(\ab[32][16] ), .Z(n1358) );
  ND2 U1384 ( .A(\SUMB[3][20] ), .B(\CARRYB[3][19] ), .Z(n835) );
  ND2 U1385 ( .A(\SUMB[3][20] ), .B(n2301), .Z(n836) );
  ND2 U1386 ( .A(\CARRYB[3][19] ), .B(n2301), .Z(n837) );
  ND3P U1387 ( .A(n835), .B(n836), .C(n837), .Z(\CARRYB[4][19] ) );
  EOP U1388 ( .A(\SUMB[37][23] ), .B(n838), .Z(\SUMB[38][22] ) );
  ND2 U1389 ( .A(\SUMB[37][23] ), .B(\CARRYB[37][22] ), .Z(n839) );
  ND2 U1390 ( .A(\SUMB[37][23] ), .B(\ab[38][22] ), .Z(n840) );
  ND2 U1391 ( .A(\CARRYB[37][22] ), .B(\ab[38][22] ), .Z(n841) );
  EO3 U1392 ( .A(\CARRYB[31][24] ), .B(\ab[32][24] ), .C(\SUMB[31][25] ), .Z(
        \SUMB[32][24] ) );
  ND2 U1393 ( .A(\CARRYB[31][24] ), .B(\SUMB[31][25] ), .Z(n842) );
  ND2 U1394 ( .A(\CARRYB[31][24] ), .B(\ab[32][24] ), .Z(n843) );
  ND2 U1395 ( .A(\SUMB[31][25] ), .B(\ab[32][24] ), .Z(n844) );
  ND3 U1396 ( .A(n842), .B(n843), .C(n844), .Z(\CARRYB[32][24] ) );
  EO U1397 ( .A(\SUMB[45][22] ), .B(n845), .Z(\SUMB[46][21] ) );
  EO3 U1398 ( .A(\SUMB[19][35] ), .B(\ab[34][20] ), .C(\CARRYB[19][34] ), .Z(
        \SUMB[20][34] ) );
  ND2 U1399 ( .A(\SUMB[19][35] ), .B(\CARRYB[19][34] ), .Z(n846) );
  ND2 U1400 ( .A(\SUMB[19][35] ), .B(\ab[34][20] ), .Z(n847) );
  ND2 U1401 ( .A(\CARRYB[19][34] ), .B(\ab[34][20] ), .Z(n848) );
  ND3 U1402 ( .A(n846), .B(n847), .C(n848), .Z(\CARRYB[20][34] ) );
  EO3P U1403 ( .A(\CARRYB[19][20] ), .B(n2360), .C(\SUMB[19][21] ), .Z(
        \SUMB[20][20] ) );
  ND2 U1404 ( .A(\CARRYB[19][20] ), .B(\SUMB[19][21] ), .Z(n849) );
  ND2 U1405 ( .A(\CARRYB[19][20] ), .B(n2360), .Z(n850) );
  ND2 U1406 ( .A(\SUMB[19][21] ), .B(n2360), .Z(n851) );
  ND3 U1407 ( .A(n849), .B(n850), .C(n851), .Z(\CARRYB[20][20] ) );
  ND2 U1408 ( .A(\CARRYB[1][46] ), .B(n2257), .Z(n853) );
  ND2 U1409 ( .A(\CARRYB[1][46] ), .B(n2245), .Z(n854) );
  ND2 U1410 ( .A(n2257), .B(n2245), .Z(n855) );
  IV U1411 ( .A(\ab[1][1] ), .Z(n2318) );
  EOP U1412 ( .A(\SUMB[39][27] ), .B(n856), .Z(\SUMB[40][26] ) );
  ND2 U1413 ( .A(\SUMB[39][27] ), .B(\CARRYB[39][26] ), .Z(n857) );
  ND2 U1414 ( .A(\SUMB[39][27] ), .B(\ab[40][26] ), .Z(n858) );
  ND2 U1415 ( .A(\CARRYB[39][26] ), .B(\ab[40][26] ), .Z(n859) );
  ND3 U1416 ( .A(n857), .B(n858), .C(n859), .Z(\CARRYB[40][26] ) );
  EOP U1417 ( .A(\CARRYB[10][27] ), .B(n620), .Z(n860) );
  ND2 U1418 ( .A(\SUMB[10][28] ), .B(\CARRYB[10][27] ), .Z(n861) );
  ND2 U1419 ( .A(\SUMB[10][28] ), .B(n620), .Z(n862) );
  ND2 U1420 ( .A(\CARRYB[10][27] ), .B(n620), .Z(n863) );
  ND3P U1421 ( .A(n861), .B(n862), .C(n863), .Z(\CARRYB[11][27] ) );
  EOP U1422 ( .A(\CARRYB[14][21] ), .B(n719), .Z(n1192) );
  ND3P U1423 ( .A(n1395), .B(n1396), .C(n1397), .Z(\CARRYB[33][28] ) );
  ND2 U1424 ( .A(\CARRYB[3][44] ), .B(\SUMB[3][45] ), .Z(n1615) );
  EOP U1425 ( .A(\CARRYB[14][18] ), .B(n713), .Z(n864) );
  EOP U1426 ( .A(\SUMB[14][19] ), .B(n864), .Z(\SUMB[15][18] ) );
  ND2 U1427 ( .A(\SUMB[14][19] ), .B(\CARRYB[14][18] ), .Z(n865) );
  ND2 U1428 ( .A(\SUMB[14][19] ), .B(n713), .Z(n866) );
  ND2 U1429 ( .A(\CARRYB[14][18] ), .B(n713), .Z(n867) );
  ND3 U1430 ( .A(n865), .B(n866), .C(n867), .Z(\CARRYB[15][18] ) );
  ND3 U1431 ( .A(n1042), .B(n1043), .C(n1044), .Z(\CARRYB[14][18] ) );
  AN2 U1432 ( .A(\CARRYB[47][10] ), .B(\SUMB[47][11] ), .Z(\A2[57] ) );
  EOP U1433 ( .A(\CARRYB[46][11] ), .B(\ab[47][11] ), .Z(n868) );
  EOP U1434 ( .A(\SUMB[46][12] ), .B(n868), .Z(\SUMB[47][11] ) );
  ND2 U1435 ( .A(\SUMB[46][12] ), .B(\CARRYB[46][11] ), .Z(n869) );
  ND2 U1436 ( .A(\SUMB[46][12] ), .B(\ab[47][11] ), .Z(n870) );
  ND2 U1437 ( .A(\CARRYB[46][11] ), .B(\ab[47][11] ), .Z(n871) );
  EO U1438 ( .A(\CARRYB[36][12] ), .B(\ab[37][12] ), .Z(n872) );
  EO U1439 ( .A(\SUMB[36][13] ), .B(n872), .Z(\SUMB[37][12] ) );
  ND2 U1440 ( .A(\SUMB[36][13] ), .B(\CARRYB[36][12] ), .Z(n873) );
  ND2 U1441 ( .A(\SUMB[36][13] ), .B(\ab[37][12] ), .Z(n874) );
  ND2 U1442 ( .A(\CARRYB[36][12] ), .B(\ab[37][12] ), .Z(n875) );
  ND3 U1443 ( .A(n873), .B(n874), .C(n875), .Z(\CARRYB[37][12] ) );
  EO3 U1444 ( .A(\SUMB[12][27] ), .B(n680), .C(\CARRYB[12][26] ), .Z(
        \SUMB[13][26] ) );
  EOP U1445 ( .A(\CARRYB[23][27] ), .B(\ab[27][24] ), .Z(n877) );
  EOP U1446 ( .A(\SUMB[23][28] ), .B(n877), .Z(\SUMB[24][27] ) );
  ND2 U1447 ( .A(\SUMB[23][28] ), .B(\CARRYB[23][27] ), .Z(n878) );
  ND2 U1448 ( .A(\SUMB[23][28] ), .B(\ab[27][24] ), .Z(n879) );
  ND2 U1449 ( .A(\CARRYB[23][27] ), .B(\ab[27][24] ), .Z(n880) );
  EO3P U1450 ( .A(\SUMB[25][28] ), .B(\ab[27][26] ), .C(\CARRYB[25][27] ), .Z(
        \SUMB[26][27] ) );
  ND2 U1451 ( .A(\SUMB[25][28] ), .B(\CARRYB[25][27] ), .Z(n881) );
  ND2 U1452 ( .A(\SUMB[25][28] ), .B(\ab[27][26] ), .Z(n882) );
  ND2 U1453 ( .A(\CARRYB[25][27] ), .B(\ab[27][26] ), .Z(n883) );
  EO3 U1454 ( .A(\CARRYB[45][22] ), .B(\ab[46][22] ), .C(\SUMB[45][23] ), .Z(
        \SUMB[46][22] ) );
  ND2 U1455 ( .A(\CARRYB[45][22] ), .B(\SUMB[45][23] ), .Z(n884) );
  ND2 U1456 ( .A(\CARRYB[45][22] ), .B(\ab[46][22] ), .Z(n885) );
  ND2 U1457 ( .A(\SUMB[45][23] ), .B(\ab[46][22] ), .Z(n886) );
  ND2P U1458 ( .A(\SUMB[38][26] ), .B(\ab[39][25] ), .Z(n1354) );
  ND2P U1459 ( .A(\SUMB[38][26] ), .B(\CARRYB[38][25] ), .Z(n1353) );
  ND3P U1460 ( .A(n2086), .B(n2087), .C(n2088), .Z(\CARRYB[8][14] ) );
  AN2P U1461 ( .A(n2419), .B(PRODUCT[0]), .Z(n887) );
  EO3P U1462 ( .A(\SUMB[7][20] ), .B(n540), .C(\CARRYB[7][19] ), .Z(
        \SUMB[8][19] ) );
  ND2 U1463 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Z(n888) );
  ND2 U1464 ( .A(\SUMB[7][20] ), .B(n540), .Z(n889) );
  ND2 U1465 ( .A(\CARRYB[7][19] ), .B(n540), .Z(n890) );
  ND3 U1466 ( .A(n888), .B(n889), .C(n890), .Z(\CARRYB[8][19] ) );
  AN2P U1467 ( .A(n2237), .B(n2243), .Z(n891) );
  IVDA U1468 ( .A(n2173), .Z(n892) );
  AN2 U1469 ( .A(\ab[20][20] ), .B(n243), .Z(n2173) );
  ND2 U1470 ( .A(\SUMB[45][19] ), .B(\CARRYB[45][18] ), .Z(n1426) );
  ND2 U1471 ( .A(\SUMB[45][19] ), .B(\ab[46][18] ), .Z(n1427) );
  EOP U1472 ( .A(n2227), .B(n2223), .Z(\SUMB[1][22] ) );
  EOP U1473 ( .A(\CARRYB[47][21] ), .B(\SUMB[47][22] ), .Z(\A1[67] ) );
  AN2P U1474 ( .A(A[22]), .B(PRODUCT[0]), .Z(n2316) );
  ND2 U1475 ( .A(\SUMB[32][15] ), .B(n894), .Z(n895) );
  ND2 U1476 ( .A(n893), .B(n1027), .Z(n896) );
  ND2 U1477 ( .A(n895), .B(n896), .Z(\SUMB[33][14] ) );
  IVDA U1478 ( .A(\SUMB[32][15] ), .Y(n893) );
  IV U1479 ( .A(n1027), .Z(n894) );
  EO3P U1480 ( .A(\CARRYB[6][26] ), .B(n468), .C(\SUMB[6][27] ), .Z(
        \SUMB[7][26] ) );
  ND2 U1481 ( .A(\CARRYB[6][26] ), .B(\SUMB[6][27] ), .Z(n897) );
  ND2 U1482 ( .A(\CARRYB[6][26] ), .B(n468), .Z(n898) );
  ND2 U1483 ( .A(\SUMB[6][27] ), .B(n468), .Z(n899) );
  ND3 U1484 ( .A(n897), .B(n898), .C(n899), .Z(\CARRYB[7][26] ) );
  IVA U1485 ( .A(\CARRYB[25][18] ), .Z(n900) );
  EO3 U1486 ( .A(\CARRYB[34][26] ), .B(\ab[35][26] ), .C(\SUMB[34][27] ), .Z(
        \SUMB[35][26] ) );
  ND2 U1487 ( .A(\CARRYB[34][26] ), .B(\SUMB[34][27] ), .Z(n902) );
  ND2 U1488 ( .A(\CARRYB[34][26] ), .B(\ab[35][26] ), .Z(n903) );
  ND2 U1489 ( .A(\SUMB[34][27] ), .B(\ab[35][26] ), .Z(n904) );
  ND3P U1490 ( .A(n902), .B(n903), .C(n904), .Z(\CARRYB[35][26] ) );
  EOP U1491 ( .A(\SUMB[10][38] ), .B(n905), .Z(\SUMB[11][37] ) );
  ND2 U1492 ( .A(\SUMB[10][38] ), .B(\CARRYB[10][37] ), .Z(n906) );
  ND2 U1493 ( .A(\SUMB[10][38] ), .B(n656), .Z(n907) );
  ND2 U1494 ( .A(\CARRYB[10][37] ), .B(n656), .Z(n908) );
  EOP U1495 ( .A(\CARRYB[34][24] ), .B(\ab[35][24] ), .Z(n909) );
  EOP U1496 ( .A(\SUMB[34][25] ), .B(n909), .Z(\SUMB[35][24] ) );
  ND2P U1497 ( .A(\SUMB[34][25] ), .B(\ab[35][24] ), .Z(n911) );
  ND2 U1498 ( .A(\CARRYB[34][24] ), .B(\ab[35][24] ), .Z(n912) );
  ND3P U1499 ( .A(n910), .B(n911), .C(n912), .Z(\CARRYB[35][24] ) );
  ND2 U1500 ( .A(\CARRYB[15][31] ), .B(\ab[31][16] ), .Z(n1414) );
  ND2 U1501 ( .A(n913), .B(n1230), .Z(n916) );
  ND2P U1502 ( .A(n915), .B(n916), .Z(\SUMB[31][19] ) );
  IVP U1503 ( .A(n1230), .Z(n914) );
  ND3 U1504 ( .A(n2104), .B(n2105), .C(n2106), .Z(\CARRYB[32][4] ) );
  EO3 U1505 ( .A(\SUMB[2][25] ), .B(n2289), .C(\CARRYB[2][24] ), .Z(
        \SUMB[3][24] ) );
  ND2 U1506 ( .A(\SUMB[2][25] ), .B(\CARRYB[2][24] ), .Z(n917) );
  ND2 U1507 ( .A(\SUMB[2][25] ), .B(n2289), .Z(n918) );
  ND2 U1508 ( .A(\CARRYB[2][24] ), .B(n2289), .Z(n919) );
  EO U1509 ( .A(\SUMB[24][2] ), .B(n2177), .Z(n2049) );
  EO U1510 ( .A(\CARRYB[20][26] ), .B(\ab[26][21] ), .Z(n920) );
  EOP U1511 ( .A(\SUMB[20][27] ), .B(n920), .Z(\SUMB[21][26] ) );
  ND2 U1512 ( .A(\SUMB[20][27] ), .B(\CARRYB[20][26] ), .Z(n921) );
  ND2 U1513 ( .A(\SUMB[20][27] ), .B(\ab[26][21] ), .Z(n922) );
  ND2 U1514 ( .A(\CARRYB[20][26] ), .B(\ab[26][21] ), .Z(n923) );
  ND3P U1515 ( .A(n921), .B(n922), .C(n923), .Z(\CARRYB[21][26] ) );
  EO3P U1516 ( .A(\CARRYB[9][30] ), .B(n580), .C(\SUMB[9][31] ), .Z(
        \SUMB[10][30] ) );
  ND2 U1517 ( .A(\CARRYB[9][30] ), .B(\SUMB[9][31] ), .Z(n924) );
  ND2 U1518 ( .A(\CARRYB[9][30] ), .B(n580), .Z(n925) );
  ND2 U1519 ( .A(\SUMB[9][31] ), .B(n580), .Z(n926) );
  EO3 U1520 ( .A(\CARRYB[45][14] ), .B(\ab[46][14] ), .C(\SUMB[45][15] ), .Z(
        \SUMB[46][14] ) );
  ND2 U1521 ( .A(\SUMB[45][15] ), .B(\ab[46][14] ), .Z(n929) );
  EOP U1522 ( .A(\SUMB[34][21] ), .B(n930), .Z(\SUMB[35][20] ) );
  ND2 U1523 ( .A(\SUMB[34][21] ), .B(\CARRYB[34][20] ), .Z(n931) );
  ND2 U1524 ( .A(\SUMB[34][21] ), .B(\ab[35][20] ), .Z(n932) );
  ND2 U1525 ( .A(\CARRYB[34][20] ), .B(\ab[35][20] ), .Z(n933) );
  EO3P U1526 ( .A(\CARRYB[17][27] ), .B(\ab[27][18] ), .C(\SUMB[17][28] ), .Z(
        \SUMB[18][27] ) );
  ND2 U1527 ( .A(\CARRYB[17][27] ), .B(\SUMB[17][28] ), .Z(n934) );
  ND2 U1528 ( .A(\CARRYB[17][27] ), .B(\ab[27][18] ), .Z(n935) );
  ND2 U1529 ( .A(\SUMB[17][28] ), .B(\ab[27][18] ), .Z(n936) );
  ND3 U1530 ( .A(n1548), .B(n1549), .C(n1550), .Z(\CARRYB[20][26] ) );
  ND3 U1531 ( .A(n1413), .B(n1414), .C(n1415), .Z(\CARRYB[16][31] ) );
  EOP U1532 ( .A(\CARRYB[38][5] ), .B(n396), .Z(n938) );
  ND2 U1533 ( .A(\CARRYB[38][5] ), .B(n396), .Z(n941) );
  ND3P U1534 ( .A(n939), .B(n940), .C(n941), .Z(\CARRYB[39][5] ) );
  EO3P U1535 ( .A(\SUMB[41][28] ), .B(\CARRYB[41][27] ), .C(\ab[42][27] ), .Z(
        \SUMB[42][27] ) );
  EOP U1536 ( .A(\ab[43][26] ), .B(\CARRYB[42][26] ), .Z(n942) );
  ND2 U1537 ( .A(\ab[42][27] ), .B(\CARRYB[41][27] ), .Z(n943) );
  ND2 U1538 ( .A(\ab[42][27] ), .B(\SUMB[41][28] ), .Z(n944) );
  ND2 U1539 ( .A(\CARRYB[41][27] ), .B(\SUMB[41][28] ), .Z(n945) );
  ND2 U1540 ( .A(\ab[43][26] ), .B(\CARRYB[42][26] ), .Z(n946) );
  ND2P U1541 ( .A(\CARRYB[42][26] ), .B(\SUMB[42][27] ), .Z(n948) );
  ND3P U1542 ( .A(n946), .B(n947), .C(n948), .Z(\CARRYB[43][26] ) );
  ND2 U1543 ( .A(\SUMB[26][34] ), .B(\CARRYB[26][33] ), .Z(n950) );
  ND2 U1544 ( .A(\SUMB[26][34] ), .B(\ab[33][27] ), .Z(n951) );
  ND2 U1545 ( .A(\CARRYB[26][33] ), .B(\ab[33][27] ), .Z(n952) );
  EO3P U1546 ( .A(\CARRYB[11][12] ), .B(n265), .C(\SUMB[11][13] ), .Z(
        \SUMB[12][12] ) );
  ND2 U1547 ( .A(\CARRYB[11][12] ), .B(\SUMB[11][13] ), .Z(n953) );
  ND2 U1548 ( .A(\CARRYB[11][12] ), .B(n265), .Z(n954) );
  ND2 U1549 ( .A(\SUMB[11][13] ), .B(n265), .Z(n955) );
  EO3 U1550 ( .A(\SUMB[12][12] ), .B(n635), .C(\CARRYB[12][11] ), .Z(
        \SUMB[13][11] ) );
  ND2P U1551 ( .A(\CARRYB[12][11] ), .B(n635), .Z(n958) );
  ND3P U1552 ( .A(n956), .B(n957), .C(n958), .Z(\CARRYB[13][11] ) );
  EO3 U1553 ( .A(\CARRYB[32][12] ), .B(n653), .C(\SUMB[32][13] ), .Z(
        \SUMB[33][12] ) );
  ND2 U1554 ( .A(\CARRYB[32][12] ), .B(\SUMB[32][13] ), .Z(n959) );
  ND2 U1555 ( .A(\CARRYB[32][12] ), .B(n653), .Z(n960) );
  ND2 U1556 ( .A(\SUMB[32][13] ), .B(n653), .Z(n961) );
  ND3 U1557 ( .A(n959), .B(n960), .C(n961), .Z(\CARRYB[33][12] ) );
  EOP U1558 ( .A(\SUMB[36][10] ), .B(n569), .Z(n962) );
  EOP U1559 ( .A(\CARRYB[36][9] ), .B(n962), .Z(\SUMB[37][9] ) );
  EO3 U1560 ( .A(\SUMB[25][34] ), .B(\ab[33][26] ), .C(\CARRYB[25][33] ), .Z(
        \SUMB[26][33] ) );
  ND2 U1561 ( .A(\SUMB[25][34] ), .B(\CARRYB[25][33] ), .Z(n963) );
  ND2 U1562 ( .A(\SUMB[25][34] ), .B(\ab[33][26] ), .Z(n964) );
  ND2 U1563 ( .A(\CARRYB[25][33] ), .B(\ab[33][26] ), .Z(n965) );
  ND3P U1564 ( .A(n963), .B(n964), .C(n965), .Z(\CARRYB[26][33] ) );
  ND2P U1565 ( .A(\CARRYB[4][17] ), .B(\SUMB[4][18] ), .Z(n967) );
  ND2P U1566 ( .A(\CARRYB[4][17] ), .B(n398), .Z(n968) );
  ND2 U1567 ( .A(\SUMB[4][18] ), .B(n398), .Z(n969) );
  ND3P U1568 ( .A(n967), .B(n968), .C(n969), .Z(\CARRYB[5][17] ) );
  EOP U1569 ( .A(\CARRYB[2][18] ), .B(n2278), .Z(n970) );
  EOP U1570 ( .A(\SUMB[2][19] ), .B(n970), .Z(\SUMB[3][18] ) );
  EOP U1571 ( .A(\CARRYB[27][18] ), .B(\ab[28][18] ), .Z(n971) );
  EOP U1572 ( .A(\SUMB[27][19] ), .B(n971), .Z(\SUMB[28][18] ) );
  ND2 U1573 ( .A(\SUMB[27][19] ), .B(\CARRYB[27][18] ), .Z(n972) );
  ND2 U1574 ( .A(\SUMB[27][19] ), .B(\ab[28][18] ), .Z(n973) );
  ND2 U1575 ( .A(\CARRYB[27][18] ), .B(\ab[28][18] ), .Z(n974) );
  ND3P U1576 ( .A(n972), .B(n973), .C(n974), .Z(\CARRYB[28][18] ) );
  EOP U1577 ( .A(\CARRYB[25][18] ), .B(\ab[26][18] ), .Z(n975) );
  EOP U1578 ( .A(\SUMB[25][19] ), .B(n975), .Z(\SUMB[26][18] ) );
  ND2 U1579 ( .A(\SUMB[25][19] ), .B(n901), .Z(n976) );
  ND2 U1580 ( .A(\SUMB[25][19] ), .B(\ab[26][18] ), .Z(n977) );
  ND2 U1581 ( .A(n901), .B(\ab[26][18] ), .Z(n978) );
  ND3 U1582 ( .A(n976), .B(n977), .C(n978), .Z(\CARRYB[26][18] ) );
  ND3 U1583 ( .A(n1449), .B(n1450), .C(n1451), .Z(\CARRYB[43][29] ) );
  EO U1584 ( .A(\SUMB[13][25] ), .B(n1286), .Z(\SUMB[14][24] ) );
  ND2 U1585 ( .A(\SUMB[42][32] ), .B(\CARRYB[42][31] ), .Z(n980) );
  ND2 U1586 ( .A(\SUMB[42][32] ), .B(\ab[43][31] ), .Z(n981) );
  ND2 U1587 ( .A(\CARRYB[42][31] ), .B(\ab[43][31] ), .Z(n982) );
  ND3P U1588 ( .A(n980), .B(n981), .C(n982), .Z(\CARRYB[43][31] ) );
  ND2 U1589 ( .A(\SUMB[13][31] ), .B(\CARRYB[13][30] ), .Z(n984) );
  ND2 U1590 ( .A(\SUMB[13][31] ), .B(n705), .Z(n985) );
  ND2 U1591 ( .A(\CARRYB[13][30] ), .B(n705), .Z(n986) );
  ND3P U1592 ( .A(n984), .B(n985), .C(n986), .Z(\CARRYB[14][30] ) );
  EO3P U1593 ( .A(\CARRYB[32][6] ), .B(n433), .C(\SUMB[32][7] ), .Z(
        \SUMB[33][6] ) );
  ND2P U1594 ( .A(\CARRYB[32][6] ), .B(\SUMB[32][7] ), .Z(n987) );
  ND2P U1595 ( .A(\CARRYB[32][6] ), .B(n433), .Z(n988) );
  ND2 U1596 ( .A(\SUMB[32][7] ), .B(n433), .Z(n989) );
  ND3P U1597 ( .A(n987), .B(n988), .C(n989), .Z(\CARRYB[33][6] ) );
  EO3P U1598 ( .A(\SUMB[18][10] ), .B(n556), .C(\CARRYB[18][9] ), .Z(
        \SUMB[19][9] ) );
  ND2 U1599 ( .A(\SUMB[18][10] ), .B(\CARRYB[18][9] ), .Z(n990) );
  ND2 U1600 ( .A(\SUMB[18][10] ), .B(n556), .Z(n991) );
  ND2 U1601 ( .A(\CARRYB[18][9] ), .B(n556), .Z(n992) );
  ND3P U1602 ( .A(n990), .B(n991), .C(n992), .Z(\CARRYB[19][9] ) );
  EOP U1603 ( .A(\CARRYB[2][21] ), .B(n2293), .Z(n993) );
  EOP U1604 ( .A(\SUMB[2][22] ), .B(n993), .Z(\SUMB[3][21] ) );
  ND2 U1605 ( .A(\SUMB[2][22] ), .B(\CARRYB[2][21] ), .Z(n994) );
  ND2 U1606 ( .A(\SUMB[2][22] ), .B(n2293), .Z(n995) );
  ND2 U1607 ( .A(\CARRYB[2][21] ), .B(n2293), .Z(n996) );
  EOP U1608 ( .A(\CARRYB[41][21] ), .B(\ab[42][21] ), .Z(n997) );
  EOP U1609 ( .A(\SUMB[41][22] ), .B(n997), .Z(\SUMB[42][21] ) );
  ND2 U1610 ( .A(\SUMB[41][22] ), .B(\CARRYB[41][21] ), .Z(n998) );
  ND2 U1611 ( .A(\SUMB[41][22] ), .B(\ab[42][21] ), .Z(n999) );
  ND2 U1612 ( .A(\CARRYB[41][21] ), .B(\ab[42][21] ), .Z(n1000) );
  EOP U1613 ( .A(\SUMB[9][38] ), .B(n1001), .Z(\SUMB[10][37] ) );
  ND2 U1614 ( .A(\SUMB[9][38] ), .B(\CARRYB[9][37] ), .Z(n1002) );
  ND2 U1615 ( .A(\SUMB[9][38] ), .B(n599), .Z(n1003) );
  ND2 U1616 ( .A(\CARRYB[9][37] ), .B(n599), .Z(n1004) );
  ND3P U1617 ( .A(n1002), .B(n1003), .C(n1004), .Z(\CARRYB[10][37] ) );
  EO3P U1618 ( .A(\CARRYB[31][26] ), .B(\ab[32][26] ), .C(\SUMB[31][27] ), .Z(
        \SUMB[32][26] ) );
  ND2 U1619 ( .A(\CARRYB[31][26] ), .B(\SUMB[31][27] ), .Z(n1005) );
  ND2 U1620 ( .A(\CARRYB[31][26] ), .B(\ab[32][26] ), .Z(n1006) );
  ND2 U1621 ( .A(\SUMB[31][27] ), .B(\ab[32][26] ), .Z(n1007) );
  EO3P U1622 ( .A(\CARRYB[12][12] ), .B(n654), .C(\SUMB[12][13] ), .Z(
        \SUMB[13][12] ) );
  ND2 U1623 ( .A(\CARRYB[12][12] ), .B(\SUMB[12][13] ), .Z(n1008) );
  ND2 U1624 ( .A(\SUMB[12][13] ), .B(n654), .Z(n1010) );
  EOP U1625 ( .A(\CARRYB[43][16] ), .B(\ab[44][16] ), .Z(n1011) );
  EOP U1626 ( .A(\SUMB[43][17] ), .B(n1011), .Z(\SUMB[44][16] ) );
  ND2 U1627 ( .A(\SUMB[43][17] ), .B(\CARRYB[43][16] ), .Z(n1012) );
  ND2 U1628 ( .A(\SUMB[43][17] ), .B(\ab[44][16] ), .Z(n1013) );
  ND2 U1629 ( .A(\CARRYB[43][16] ), .B(\ab[44][16] ), .Z(n1014) );
  ND2 U1630 ( .A(\SUMB[24][25] ), .B(\ab[25][24] ), .Z(n1018) );
  EO3 U1631 ( .A(\CARRYB[42][27] ), .B(\ab[43][27] ), .C(\SUMB[42][28] ), .Z(
        n1019) );
  EO3P U1632 ( .A(\CARRYB[38][29] ), .B(\ab[39][29] ), .C(n29), .Z(
        \SUMB[39][29] ) );
  ND2 U1633 ( .A(\CARRYB[38][29] ), .B(\SUMB[38][30] ), .Z(n1020) );
  ND2 U1634 ( .A(\CARRYB[38][29] ), .B(\ab[39][29] ), .Z(n1021) );
  ND2 U1635 ( .A(\SUMB[38][30] ), .B(\ab[39][29] ), .Z(n1022) );
  ND3 U1636 ( .A(n1020), .B(n1021), .C(n1022), .Z(\CARRYB[39][29] ) );
  EO3 U1637 ( .A(\CARRYB[42][27] ), .B(\ab[43][27] ), .C(\SUMB[42][28] ), .Z(
        \SUMB[43][27] ) );
  ND2 U1638 ( .A(\CARRYB[19][10] ), .B(n581), .Z(n1956) );
  EOP U1639 ( .A(\CARRYB[6][15] ), .B(n475), .Z(n1023) );
  EOP U1640 ( .A(\SUMB[6][16] ), .B(n1023), .Z(\SUMB[7][15] ) );
  ND2 U1641 ( .A(\SUMB[6][16] ), .B(\CARRYB[6][15] ), .Z(n1024) );
  ND2 U1642 ( .A(\SUMB[6][16] ), .B(n475), .Z(n1025) );
  ND2 U1643 ( .A(\CARRYB[6][15] ), .B(n475), .Z(n1026) );
  AN2 U1644 ( .A(\CARRYB[47][24] ), .B(\SUMB[47][25] ), .Z(\A2[71] ) );
  EOP U1645 ( .A(\CARRYB[32][14] ), .B(\ab[33][14] ), .Z(n1027) );
  ND2 U1646 ( .A(\SUMB[32][15] ), .B(\CARRYB[32][14] ), .Z(n1028) );
  ND2 U1647 ( .A(\SUMB[32][15] ), .B(\ab[33][14] ), .Z(n1029) );
  ND2 U1648 ( .A(\CARRYB[32][14] ), .B(\ab[33][14] ), .Z(n1030) );
  ND3P U1649 ( .A(n1028), .B(n1029), .C(n1030), .Z(\CARRYB[33][14] ) );
  ND3P U1650 ( .A(n1398), .B(n1399), .C(n1400), .Z(\CARRYB[22][32] ) );
  EOP U1651 ( .A(n1394), .B(\SUMB[32][29] ), .Z(\SUMB[33][28] ) );
  ND3P U1652 ( .A(n1073), .B(n1074), .C(n1075), .Z(\CARRYB[32][27] ) );
  EO3 U1653 ( .A(\SUMB[11][16] ), .B(n655), .C(\CARRYB[11][15] ), .Z(
        \SUMB[12][15] ) );
  ND2 U1654 ( .A(\SUMB[11][16] ), .B(\CARRYB[11][15] ), .Z(n1031) );
  ND2 U1655 ( .A(\SUMB[11][16] ), .B(n655), .Z(n1032) );
  ND2 U1656 ( .A(\CARRYB[11][15] ), .B(n655), .Z(n1033) );
  ND3 U1657 ( .A(n1031), .B(n1032), .C(n1033), .Z(\CARRYB[12][15] ) );
  ND2 U1658 ( .A(\SUMB[43][26] ), .B(\CARRYB[43][25] ), .Z(n1034) );
  ND2 U1659 ( .A(\SUMB[43][26] ), .B(\ab[44][25] ), .Z(n1035) );
  ND2 U1660 ( .A(\CARRYB[43][25] ), .B(\ab[44][25] ), .Z(n1036) );
  ND2 U1661 ( .A(\SUMB[36][28] ), .B(\CARRYB[36][27] ), .Z(n1038) );
  ND2 U1662 ( .A(\SUMB[36][28] ), .B(\ab[37][27] ), .Z(n1039) );
  ND2 U1663 ( .A(\CARRYB[36][27] ), .B(\ab[37][27] ), .Z(n1040) );
  ND3 U1664 ( .A(n1038), .B(n1039), .C(n1040), .Z(\CARRYB[37][27] ) );
  ND2P U1665 ( .A(n10), .B(\SUMB[13][33] ), .Z(n2032) );
  EOP U1666 ( .A(\SUMB[13][19] ), .B(n698), .Z(n1041) );
  EOP U1667 ( .A(\CARRYB[13][18] ), .B(n1041), .Z(\SUMB[14][18] ) );
  ND2 U1668 ( .A(\CARRYB[13][18] ), .B(\SUMB[13][19] ), .Z(n1042) );
  ND2 U1669 ( .A(\CARRYB[13][18] ), .B(n698), .Z(n1043) );
  ND2 U1670 ( .A(\SUMB[13][19] ), .B(n698), .Z(n1044) );
  ND2P U1671 ( .A(\CARRYB[37][8] ), .B(\SUMB[37][9] ), .Z(n1342) );
  ND2P U1672 ( .A(\SUMB[40][16] ), .B(\ab[41][15] ), .Z(n1119) );
  ND2P U1673 ( .A(\SUMB[40][16] ), .B(n1087), .Z(n1118) );
  EOP U1674 ( .A(n2182), .B(n2177), .Z(\SUMB[1][25] ) );
  EOP U1675 ( .A(\SUMB[30][13] ), .B(n1533), .Z(\SUMB[31][12] ) );
  ND2P U1676 ( .A(\SUMB[23][11] ), .B(n772), .Z(n1490) );
  EO3P U1677 ( .A(\CARRYB[27][8] ), .B(n530), .C(\SUMB[27][9] ), .Z(
        \SUMB[28][8] ) );
  EO3 U1678 ( .A(\CARRYB[29][27] ), .B(\ab[30][27] ), .C(\SUMB[29][28] ), .Z(
        \SUMB[30][27] ) );
  ND2 U1679 ( .A(\CARRYB[29][27] ), .B(\SUMB[29][28] ), .Z(n1045) );
  ND2 U1680 ( .A(\CARRYB[29][27] ), .B(\ab[30][27] ), .Z(n1046) );
  ND2 U1681 ( .A(\SUMB[29][28] ), .B(\ab[30][27] ), .Z(n1047) );
  ND3 U1682 ( .A(n1045), .B(n1046), .C(n1047), .Z(\CARRYB[30][27] ) );
  IV U1683 ( .A(\SUMB[23][11] ), .Z(n1489) );
  AN2 U1684 ( .A(n2165), .B(n2173), .Z(\CARRYB[1][19] ) );
  FA1AP U1685 ( .A(\ab[45][17] ), .B(\CARRYB[44][17] ), .CI(\SUMB[44][18] ), 
        .S(n1048) );
  EOP U1686 ( .A(\CARRYB[16][29] ), .B(\ab[29][17] ), .Z(n1049) );
  EOP U1687 ( .A(\SUMB[16][30] ), .B(n1049), .Z(\SUMB[17][29] ) );
  ND2 U1688 ( .A(\SUMB[16][30] ), .B(\CARRYB[16][29] ), .Z(n1050) );
  ND2 U1689 ( .A(\SUMB[16][30] ), .B(\ab[29][17] ), .Z(n1051) );
  ND2 U1690 ( .A(\CARRYB[16][29] ), .B(\ab[29][17] ), .Z(n1052) );
  ND3 U1691 ( .A(n1050), .B(n1051), .C(n1052), .Z(\CARRYB[17][29] ) );
  EOP U1692 ( .A(\CARRYB[36][29] ), .B(\ab[37][29] ), .Z(n1053) );
  EOP U1693 ( .A(\SUMB[36][30] ), .B(n1053), .Z(\SUMB[37][29] ) );
  EOP U1694 ( .A(\CARRYB[20][35] ), .B(n1054), .Z(\SUMB[21][35] ) );
  EOP U1695 ( .A(\CARRYB[6][31] ), .B(n469), .Z(n1055) );
  EOP U1696 ( .A(\SUMB[6][32] ), .B(n1055), .Z(\SUMB[7][31] ) );
  ND2 U1697 ( .A(\CARRYB[6][31] ), .B(n469), .Z(n1058) );
  EOP U1698 ( .A(\CARRYB[7][31] ), .B(n514), .Z(n1059) );
  EOP U1699 ( .A(\SUMB[7][32] ), .B(n1059), .Z(\SUMB[8][31] ) );
  ND2 U1700 ( .A(\CARRYB[7][31] ), .B(n514), .Z(n1062) );
  ND3P U1701 ( .A(n1060), .B(n1061), .C(n1062), .Z(\CARRYB[8][31] ) );
  IVDA U1702 ( .A(n2184), .Z(n1063) );
  AN2 U1703 ( .A(A[35]), .B(PRODUCT[0]), .Z(n2184) );
  EO3 U1704 ( .A(\SUMB[28][16] ), .B(n714), .C(\CARRYB[28][15] ), .Z(
        \SUMB[29][15] ) );
  ND2 U1705 ( .A(\SUMB[28][16] ), .B(\CARRYB[28][15] ), .Z(n1064) );
  ND2 U1706 ( .A(\SUMB[28][16] ), .B(n714), .Z(n1065) );
  ND2 U1707 ( .A(\CARRYB[28][15] ), .B(n714), .Z(n1066) );
  ND3P U1708 ( .A(n1064), .B(n1065), .C(n1066), .Z(\CARRYB[29][15] ) );
  EO3 U1709 ( .A(\SUMB[34][13] ), .B(n672), .C(\CARRYB[34][12] ), .Z(
        \SUMB[35][12] ) );
  ND2 U1710 ( .A(\SUMB[34][13] ), .B(\CARRYB[34][12] ), .Z(n1067) );
  ND2 U1711 ( .A(\SUMB[34][13] ), .B(n672), .Z(n1068) );
  ND2 U1712 ( .A(\CARRYB[34][12] ), .B(n672), .Z(n1069) );
  ND3 U1713 ( .A(n1067), .B(n1068), .C(n1069), .Z(\CARRYB[35][12] ) );
  IVA U1714 ( .A(\CARRYB[3][36] ), .Z(n1070) );
  IV U1715 ( .A(n1070), .Z(n1071) );
  EOP U1716 ( .A(\CARRYB[31][27] ), .B(\ab[32][27] ), .Z(n1072) );
  EOP U1717 ( .A(\SUMB[31][28] ), .B(n1072), .Z(\SUMB[32][27] ) );
  ND2 U1718 ( .A(\SUMB[31][28] ), .B(\CARRYB[31][27] ), .Z(n1073) );
  ND2 U1719 ( .A(\SUMB[31][28] ), .B(\ab[32][27] ), .Z(n1074) );
  ND2 U1720 ( .A(\CARRYB[31][27] ), .B(\ab[32][27] ), .Z(n1075) );
  EOP U1721 ( .A(\CARRYB[14][32] ), .B(\ab[32][15] ), .Z(n1076) );
  EOP U1722 ( .A(\SUMB[14][33] ), .B(n1076), .Z(\SUMB[15][32] ) );
  ND2 U1723 ( .A(\SUMB[14][33] ), .B(\CARRYB[14][32] ), .Z(n1077) );
  ND2 U1724 ( .A(\SUMB[14][33] ), .B(\ab[32][15] ), .Z(n1078) );
  ND2 U1725 ( .A(\CARRYB[14][32] ), .B(\ab[32][15] ), .Z(n1079) );
  ND3P U1726 ( .A(n1077), .B(n1078), .C(n1079), .Z(\CARRYB[15][32] ) );
  ND2 U1727 ( .A(n1080), .B(n1485), .Z(n1083) );
  IVDA U1728 ( .A(\SUMB[6][36] ), .Y(n1080) );
  IV U1729 ( .A(n1485), .Z(n1081) );
  EO3 U1730 ( .A(\CARRYB[34][11] ), .B(n609), .C(\SUMB[34][12] ), .Z(
        \SUMB[35][11] ) );
  ND2 U1731 ( .A(\CARRYB[34][11] ), .B(\SUMB[34][12] ), .Z(n1084) );
  ND2 U1732 ( .A(\CARRYB[34][11] ), .B(n609), .Z(n1085) );
  ND2 U1733 ( .A(\SUMB[34][12] ), .B(n609), .Z(n1086) );
  ND3 U1734 ( .A(n1084), .B(n1085), .C(n1086), .Z(\CARRYB[35][11] ) );
  ND2 U1735 ( .A(n435), .B(\SUMB[5][33] ), .Z(n1599) );
  ND3 U1736 ( .A(n1737), .B(n1738), .C(n1739), .Z(n1087) );
  ND3 U1737 ( .A(n1737), .B(n1738), .C(n1739), .Z(\CARRYB[40][15] ) );
  EO3 U1738 ( .A(\CARRYB[15][33] ), .B(\ab[33][16] ), .C(\SUMB[15][34] ), .Z(
        \SUMB[16][33] ) );
  ND2 U1739 ( .A(\CARRYB[15][33] ), .B(\SUMB[15][34] ), .Z(n1088) );
  ND2 U1740 ( .A(\CARRYB[15][33] ), .B(\ab[33][16] ), .Z(n1089) );
  ND2 U1741 ( .A(\SUMB[15][34] ), .B(\ab[33][16] ), .Z(n1090) );
  ND3 U1742 ( .A(n1088), .B(n1089), .C(n1090), .Z(\CARRYB[16][33] ) );
  EOP U1743 ( .A(\CARRYB[24][28] ), .B(\ab[28][25] ), .Z(n1091) );
  EOP U1744 ( .A(\SUMB[24][29] ), .B(n1091), .Z(\SUMB[25][28] ) );
  ND2 U1745 ( .A(\SUMB[24][29] ), .B(\CARRYB[24][28] ), .Z(n1092) );
  ND2 U1746 ( .A(\SUMB[24][29] ), .B(\ab[28][25] ), .Z(n1093) );
  ND2 U1747 ( .A(\CARRYB[24][28] ), .B(\ab[28][25] ), .Z(n1094) );
  EO3P U1748 ( .A(\ab[38][16] ), .B(\CARRYB[15][38] ), .C(\SUMB[15][39] ), .Z(
        \SUMB[16][38] ) );
  EOP U1749 ( .A(\ab[37][17] ), .B(\CARRYB[16][37] ), .Z(n1095) );
  EOP U1750 ( .A(n1095), .B(\SUMB[16][38] ), .Z(\SUMB[17][37] ) );
  ND2 U1751 ( .A(\ab[38][16] ), .B(\CARRYB[15][38] ), .Z(n1096) );
  ND2 U1752 ( .A(\ab[38][16] ), .B(\SUMB[15][39] ), .Z(n1097) );
  ND2 U1753 ( .A(\CARRYB[15][38] ), .B(\SUMB[15][39] ), .Z(n1098) );
  ND3P U1754 ( .A(n1096), .B(n1097), .C(n1098), .Z(\CARRYB[16][38] ) );
  ND2 U1755 ( .A(\ab[37][17] ), .B(\CARRYB[16][37] ), .Z(n1099) );
  EOP U1756 ( .A(\CARRYB[18][36] ), .B(\ab[36][19] ), .Z(n1102) );
  EOP U1757 ( .A(\SUMB[18][37] ), .B(n1102), .Z(\SUMB[19][36] ) );
  ND2 U1758 ( .A(\SUMB[18][37] ), .B(\CARRYB[18][36] ), .Z(n1103) );
  ND2 U1759 ( .A(\SUMB[18][37] ), .B(\ab[36][19] ), .Z(n1104) );
  ND2 U1760 ( .A(\CARRYB[18][36] ), .B(\ab[36][19] ), .Z(n1105) );
  ND3P U1761 ( .A(n1103), .B(n1104), .C(n1105), .Z(\CARRYB[19][36] ) );
  EO U1762 ( .A(\SUMB[33][11] ), .B(n1390), .Z(\SUMB[34][10] ) );
  AN2 U1763 ( .A(n2240), .B(n2235), .Z(\CARRYB[1][24] ) );
  ND2P U1764 ( .A(\CARRYB[39][11] ), .B(\ab[40][11] ), .Z(n1348) );
  ND2P U1765 ( .A(\CARRYB[39][11] ), .B(\SUMB[39][12] ), .Z(n1347) );
  EOP U1766 ( .A(\SUMB[7][21] ), .B(n1764), .Z(\SUMB[8][20] ) );
  ND2 U1767 ( .A(\SUMB[39][16] ), .B(n1107), .Z(n1108) );
  ND2 U1768 ( .A(n1106), .B(n1736), .Z(n1109) );
  IVDA U1769 ( .A(\SUMB[39][16] ), .Y(n1106) );
  IV U1770 ( .A(n1736), .Z(n1107) );
  EO3 U1771 ( .A(\CARRYB[3][32] ), .B(n358), .C(\SUMB[3][33] ), .Z(
        \SUMB[4][32] ) );
  EOP U1772 ( .A(\CARRYB[7][18] ), .B(n519), .Z(n1113) );
  EOP U1773 ( .A(\SUMB[7][19] ), .B(n1113), .Z(\SUMB[8][18] ) );
  ND2 U1774 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Z(n1114) );
  ND2 U1775 ( .A(\SUMB[7][19] ), .B(n519), .Z(n1115) );
  ND2 U1776 ( .A(\CARRYB[7][18] ), .B(n519), .Z(n1116) );
  ND3P U1777 ( .A(n1114), .B(n1115), .C(n1116), .Z(\CARRYB[8][18] ) );
  EOP U1778 ( .A(\SUMB[40][16] ), .B(n1117), .Z(\SUMB[41][15] ) );
  ND2 U1779 ( .A(n1087), .B(\ab[41][15] ), .Z(n1120) );
  ND3P U1780 ( .A(n1118), .B(n1119), .C(n1120), .Z(\CARRYB[41][15] ) );
  EOP U1781 ( .A(\CARRYB[39][16] ), .B(\ab[40][16] ), .Z(n1121) );
  EOP U1782 ( .A(\SUMB[39][17] ), .B(n1121), .Z(\SUMB[40][16] ) );
  ND2 U1783 ( .A(\SUMB[39][17] ), .B(\CARRYB[39][16] ), .Z(n1122) );
  ND2 U1784 ( .A(\SUMB[39][17] ), .B(\ab[40][16] ), .Z(n1123) );
  ND2 U1785 ( .A(\CARRYB[39][16] ), .B(\ab[40][16] ), .Z(n1124) );
  ND3 U1786 ( .A(n1122), .B(n1123), .C(n1124), .Z(\CARRYB[40][16] ) );
  ND2 U1787 ( .A(\CARRYB[30][9] ), .B(n562), .Z(n1559) );
  EO3 U1788 ( .A(\SUMB[9][37] ), .B(n601), .C(\CARRYB[9][36] ), .Z(
        \SUMB[10][36] ) );
  ND2 U1789 ( .A(\SUMB[9][37] ), .B(\CARRYB[9][36] ), .Z(n1125) );
  ND2 U1790 ( .A(\SUMB[9][37] ), .B(n601), .Z(n1126) );
  ND2 U1791 ( .A(\CARRYB[9][36] ), .B(n601), .Z(n1127) );
  ND3 U1792 ( .A(n1125), .B(n1126), .C(n1127), .Z(\CARRYB[10][36] ) );
  EO U1793 ( .A(n1212), .B(\CARRYB[36][4] ), .Z(\SUMB[37][4] ) );
  EOP U1794 ( .A(\CARRYB[23][32] ), .B(\ab[32][24] ), .Z(n1128) );
  EOP U1795 ( .A(\SUMB[23][33] ), .B(n1128), .Z(\SUMB[24][32] ) );
  ND2 U1796 ( .A(\SUMB[23][33] ), .B(\CARRYB[23][32] ), .Z(n1129) );
  ND2 U1797 ( .A(\SUMB[23][33] ), .B(\ab[32][24] ), .Z(n1130) );
  ND2 U1798 ( .A(\CARRYB[23][32] ), .B(\ab[32][24] ), .Z(n1131) );
  ND3P U1799 ( .A(n1129), .B(n1130), .C(n1131), .Z(\CARRYB[24][32] ) );
  ND3 U1800 ( .A(n1319), .B(n1320), .C(n1321), .Z(\CARRYB[40][5] ) );
  EO3 U1801 ( .A(\CARRYB[15][14] ), .B(n701), .C(\SUMB[15][15] ), .Z(
        \SUMB[16][14] ) );
  EO3P U1802 ( .A(n676), .B(\CARRYB[11][29] ), .C(\SUMB[11][30] ), .Z(
        \SUMB[12][29] ) );
  ND2 U1803 ( .A(n676), .B(\CARRYB[11][29] ), .Z(n1133) );
  ND2 U1804 ( .A(n676), .B(\SUMB[11][30] ), .Z(n1134) );
  ND2 U1805 ( .A(\CARRYB[11][29] ), .B(\SUMB[11][30] ), .Z(n1135) );
  ND3P U1806 ( .A(n1133), .B(n1134), .C(n1135), .Z(\CARRYB[12][29] ) );
  ND2 U1807 ( .A(n697), .B(\CARRYB[12][28] ), .Z(n1136) );
  ND2P U1808 ( .A(n697), .B(\SUMB[12][29] ), .Z(n1137) );
  ND2P U1809 ( .A(\CARRYB[12][28] ), .B(\SUMB[12][29] ), .Z(n1138) );
  ND3P U1810 ( .A(n1136), .B(n1137), .C(n1138), .Z(\CARRYB[13][28] ) );
  ND2 U1811 ( .A(\SUMB[45][16] ), .B(\CARRYB[45][15] ), .Z(n1140) );
  ND2 U1812 ( .A(\SUMB[45][16] ), .B(\ab[46][15] ), .Z(n1141) );
  ND2 U1813 ( .A(\CARRYB[45][15] ), .B(\ab[46][15] ), .Z(n1142) );
  EOP U1814 ( .A(\CARRYB[35][19] ), .B(\ab[36][19] ), .Z(n1143) );
  ND2P U1815 ( .A(\SUMB[35][20] ), .B(\CARRYB[35][19] ), .Z(n1144) );
  ND2P U1816 ( .A(\SUMB[35][20] ), .B(\ab[36][19] ), .Z(n1145) );
  ND3P U1817 ( .A(n1144), .B(n1145), .C(n1146), .Z(\CARRYB[36][19] ) );
  ND2P U1818 ( .A(\CARRYB[36][19] ), .B(\ab[37][19] ), .Z(n1577) );
  ND2 U1819 ( .A(\CARRYB[20][25] ), .B(\SUMB[20][26] ), .Z(n1553) );
  EO U1820 ( .A(n1547), .B(\SUMB[20][26] ), .Z(\SUMB[21][25] ) );
  ND2P U1821 ( .A(\CARRYB[23][20] ), .B(\ab[24][20] ), .Z(n1188) );
  AN2 U1822 ( .A(n2222), .B(n2225), .Z(\CARRYB[1][41] ) );
  EO3P U1823 ( .A(\SUMB[37][13] ), .B(\ab[38][12] ), .C(\CARRYB[37][12] ), .Z(
        \SUMB[38][12] ) );
  ND2 U1824 ( .A(\SUMB[37][13] ), .B(\CARRYB[37][12] ), .Z(n1148) );
  ND2 U1825 ( .A(\SUMB[37][13] ), .B(\ab[38][12] ), .Z(n1149) );
  ND2 U1826 ( .A(\CARRYB[37][12] ), .B(\ab[38][12] ), .Z(n1150) );
  ND3 U1827 ( .A(n1255), .B(n1256), .C(n1257), .Z(\CARRYB[37][13] ) );
  ND2 U1828 ( .A(\CARRYB[25][15] ), .B(\SUMB[25][16] ), .Z(n1788) );
  EO3 U1829 ( .A(\SUMB[12][33] ), .B(n694), .C(\CARRYB[12][32] ), .Z(
        \SUMB[13][32] ) );
  ND2P U1830 ( .A(\CARRYB[12][32] ), .B(\SUMB[12][33] ), .Z(n1151) );
  ND2P U1831 ( .A(\CARRYB[12][32] ), .B(n694), .Z(n1152) );
  ND2P U1832 ( .A(\SUMB[12][33] ), .B(n694), .Z(n1153) );
  ND2 U1833 ( .A(\SUMB[31][5] ), .B(\CARRYB[31][4] ), .Z(n2106) );
  ND2 U1834 ( .A(\SUMB[28][35] ), .B(\CARRYB[28][34] ), .Z(n1155) );
  ND2 U1835 ( .A(\SUMB[28][35] ), .B(\ab[34][29] ), .Z(n1156) );
  ND2 U1836 ( .A(\CARRYB[28][34] ), .B(\ab[34][29] ), .Z(n1157) );
  ND2 U1837 ( .A(\CARRYB[27][35] ), .B(\SUMB[27][36] ), .Z(n1158) );
  ND2 U1838 ( .A(\CARRYB[27][35] ), .B(\ab[35][28] ), .Z(n1159) );
  ND2 U1839 ( .A(\SUMB[27][36] ), .B(\ab[35][28] ), .Z(n1160) );
  ND3 U1840 ( .A(n1158), .B(n1159), .C(n1160), .Z(\CARRYB[28][35] ) );
  EO3P U1841 ( .A(\CARRYB[13][32] ), .B(\ab[32][14] ), .C(\SUMB[13][33] ), .Z(
        \SUMB[14][32] ) );
  EO3 U1842 ( .A(\CARRYB[15][29] ), .B(\ab[29][16] ), .C(\SUMB[15][30] ), .Z(
        \SUMB[16][29] ) );
  AN2 U1843 ( .A(n2221), .B(n2205), .Z(\CARRYB[1][39] ) );
  EO3 U1844 ( .A(\SUMB[45][11] ), .B(\ab[46][10] ), .C(\CARRYB[45][10] ), .Z(
        \SUMB[46][10] ) );
  ND2 U1845 ( .A(\CARRYB[45][10] ), .B(\SUMB[45][11] ), .Z(n1161) );
  ND2 U1846 ( .A(\CARRYB[45][10] ), .B(\ab[46][10] ), .Z(n1162) );
  ND2 U1847 ( .A(\SUMB[45][11] ), .B(\ab[46][10] ), .Z(n1163) );
  ND3 U1848 ( .A(n1161), .B(n1162), .C(n1163), .Z(\CARRYB[46][10] ) );
  EO3 U1849 ( .A(\CARRYB[28][14] ), .B(n702), .C(\SUMB[28][15] ), .Z(
        \SUMB[29][14] ) );
  ND2 U1850 ( .A(\CARRYB[28][14] ), .B(\SUMB[28][15] ), .Z(n1164) );
  ND2 U1851 ( .A(\CARRYB[28][14] ), .B(n702), .Z(n1165) );
  ND2 U1852 ( .A(\SUMB[28][15] ), .B(n702), .Z(n1166) );
  ND3 U1853 ( .A(n1164), .B(n1165), .C(n1166), .Z(\CARRYB[29][14] ) );
  EO3 U1854 ( .A(\CARRYB[11][25] ), .B(n661), .C(\SUMB[11][26] ), .Z(
        \SUMB[12][25] ) );
  ND2 U1855 ( .A(\SUMB[11][26] ), .B(n661), .Z(n1169) );
  ND3P U1856 ( .A(n1167), .B(n1168), .C(n1169), .Z(\CARRYB[12][25] ) );
  EO3 U1857 ( .A(\CARRYB[40][4] ), .B(n379), .C(\SUMB[40][5] ), .Z(
        \SUMB[41][4] ) );
  ND2P U1858 ( .A(\CARRYB[40][4] ), .B(\SUMB[40][5] ), .Z(n1170) );
  ND2 U1859 ( .A(\CARRYB[40][4] ), .B(n379), .Z(n1171) );
  ND2P U1860 ( .A(\SUMB[40][5] ), .B(n379), .Z(n1172) );
  ND3P U1861 ( .A(n1170), .B(n1171), .C(n1172), .Z(\CARRYB[41][4] ) );
  EO3 U1862 ( .A(\SUMB[15][12] ), .B(n624), .C(\CARRYB[15][11] ), .Z(
        \SUMB[16][11] ) );
  ND2 U1863 ( .A(\SUMB[15][12] ), .B(\CARRYB[15][11] ), .Z(n1173) );
  ND2 U1864 ( .A(\SUMB[15][12] ), .B(n624), .Z(n1174) );
  ND2 U1865 ( .A(\CARRYB[15][11] ), .B(n624), .Z(n1175) );
  EOP U1866 ( .A(\CARRYB[16][11] ), .B(n629), .Z(n1176) );
  EOP U1867 ( .A(\SUMB[16][12] ), .B(n1176), .Z(\SUMB[17][11] ) );
  ND2 U1868 ( .A(\SUMB[16][12] ), .B(\CARRYB[16][11] ), .Z(n1177) );
  ND2 U1869 ( .A(\SUMB[16][12] ), .B(n629), .Z(n1178) );
  ND2 U1870 ( .A(\CARRYB[16][11] ), .B(n629), .Z(n1179) );
  ND3P U1871 ( .A(n1177), .B(n1178), .C(n1179), .Z(\CARRYB[17][11] ) );
  EO3 U1872 ( .A(\SUMB[6][17] ), .B(n479), .C(\CARRYB[6][16] ), .Z(
        \SUMB[7][16] ) );
  ND2 U1873 ( .A(\SUMB[6][17] ), .B(n479), .Z(n1181) );
  ND3P U1874 ( .A(n1180), .B(n1181), .C(n1182), .Z(\CARRYB[7][16] ) );
  EO U1875 ( .A(n1908), .B(\CARRYB[43][15] ), .Z(\SUMB[44][15] ) );
  ND3 U1876 ( .A(n1618), .B(n1619), .C(n1620), .Z(\CARRYB[23][24] ) );
  AN2P U1877 ( .A(n2179), .B(n2316), .Z(\CARRYB[1][21] ) );
  ND2 U1878 ( .A(\SUMB[21][15] ), .B(\CARRYB[21][14] ), .Z(n1183) );
  ND2 U1879 ( .A(\SUMB[21][15] ), .B(n700), .Z(n1184) );
  ND2 U1880 ( .A(\CARRYB[21][14] ), .B(n700), .Z(n1185) );
  ND3P U1881 ( .A(n1183), .B(n1184), .C(n1185), .Z(\CARRYB[22][14] ) );
  EO3 U1882 ( .A(\SUMB[23][21] ), .B(\ab[24][20] ), .C(\CARRYB[23][20] ), .Z(
        \SUMB[24][20] ) );
  ND2 U1883 ( .A(\SUMB[23][21] ), .B(\CARRYB[23][20] ), .Z(n1186) );
  ND2 U1884 ( .A(\SUMB[23][21] ), .B(\ab[24][20] ), .Z(n1187) );
  ND3P U1885 ( .A(n1186), .B(n1187), .C(n1188), .Z(\CARRYB[24][20] ) );
  ND2 U1886 ( .A(\CARRYB[8][15] ), .B(n559), .Z(n1636) );
  AN2P U1887 ( .A(n2202), .B(n2204), .Z(\CARRYB[1][43] ) );
  EO3 U1888 ( .A(\SUMB[30][15] ), .B(\ab[31][14] ), .C(\CARRYB[30][14] ), .Z(
        \SUMB[31][14] ) );
  ND2 U1889 ( .A(\SUMB[30][15] ), .B(\ab[31][14] ), .Z(n1191) );
  ND3P U1890 ( .A(n1189), .B(n1190), .C(n1191), .Z(\CARRYB[31][14] ) );
  EOP U1891 ( .A(\SUMB[14][22] ), .B(n1192), .Z(\SUMB[15][21] ) );
  ND2 U1892 ( .A(\SUMB[14][22] ), .B(\CARRYB[14][21] ), .Z(n1193) );
  ND2 U1893 ( .A(\SUMB[14][22] ), .B(n719), .Z(n1194) );
  ND2 U1894 ( .A(\CARRYB[14][21] ), .B(n719), .Z(n1195) );
  ND3P U1895 ( .A(n1193), .B(n1194), .C(n1195), .Z(\CARRYB[15][21] ) );
  ND3P U1896 ( .A(n1503), .B(n1504), .C(n1505), .Z(\CARRYB[14][21] ) );
  EO3P U1897 ( .A(\SUMB[43][27] ), .B(\ab[44][26] ), .C(\CARRYB[43][26] ), .Z(
        \SUMB[44][26] ) );
  ND2 U1898 ( .A(n1019), .B(\CARRYB[43][26] ), .Z(n1196) );
  ND2 U1899 ( .A(n1019), .B(\ab[44][26] ), .Z(n1197) );
  ND2 U1900 ( .A(\CARRYB[43][26] ), .B(\ab[44][26] ), .Z(n1198) );
  ND3P U1901 ( .A(n1196), .B(n1197), .C(n1198), .Z(\CARRYB[44][26] ) );
  ND2 U1902 ( .A(\ab[35][21] ), .B(\CARRYB[20][35] ), .Z(n1200) );
  ND2 U1903 ( .A(\ab[35][21] ), .B(\SUMB[20][36] ), .Z(n1201) );
  ND2 U1904 ( .A(\CARRYB[20][35] ), .B(\SUMB[20][36] ), .Z(n1202) );
  ND2 U1905 ( .A(\ab[34][22] ), .B(\CARRYB[21][34] ), .Z(n1203) );
  ND2P U1906 ( .A(\CARRYB[21][34] ), .B(\SUMB[21][35] ), .Z(n1205) );
  ND2 U1907 ( .A(\CARRYB[5][32] ), .B(\SUMB[5][33] ), .Z(n1600) );
  ND2 U1908 ( .A(\CARRYB[42][27] ), .B(\SUMB[42][28] ), .Z(n1206) );
  ND2 U1909 ( .A(\CARRYB[42][27] ), .B(\ab[43][27] ), .Z(n1207) );
  ND2 U1910 ( .A(\SUMB[42][28] ), .B(\ab[43][27] ), .Z(n1208) );
  EO3P U1911 ( .A(\CARRYB[22][28] ), .B(\ab[28][23] ), .C(\SUMB[22][29] ), .Z(
        \SUMB[23][28] ) );
  EO3P U1912 ( .A(n2300), .B(\CARRYB[35][4] ), .C(\SUMB[35][5] ), .Z(
        \SUMB[36][4] ) );
  ND2 U1913 ( .A(n2300), .B(\CARRYB[35][4] ), .Z(n1209) );
  ND2 U1914 ( .A(n2300), .B(\SUMB[35][5] ), .Z(n1210) );
  ND2 U1915 ( .A(\CARRYB[35][4] ), .B(\SUMB[35][5] ), .Z(n1211) );
  ND3P U1916 ( .A(n1209), .B(n1210), .C(n1211), .Z(\CARRYB[36][4] ) );
  EOP U1917 ( .A(n361), .B(\SUMB[36][5] ), .Z(n1212) );
  ND2 U1918 ( .A(n361), .B(\SUMB[36][5] ), .Z(n1213) );
  ND2 U1919 ( .A(n361), .B(\CARRYB[36][4] ), .Z(n1214) );
  ND2 U1920 ( .A(\SUMB[36][5] ), .B(\CARRYB[36][4] ), .Z(n1215) );
  ND3P U1921 ( .A(n1213), .B(n1214), .C(n1215), .Z(\CARRYB[37][4] ) );
  EO3P U1922 ( .A(\CARRYB[24][7] ), .B(n467), .C(\SUMB[24][8] ), .Z(
        \SUMB[25][7] ) );
  ND2 U1923 ( .A(\CARRYB[24][7] ), .B(n467), .Z(n1217) );
  ND2 U1924 ( .A(\CARRYB[24][7] ), .B(\SUMB[24][8] ), .Z(n1218) );
  ND2 U1925 ( .A(n467), .B(\SUMB[24][8] ), .Z(n1219) );
  ND3P U1926 ( .A(n1217), .B(n1218), .C(n1219), .Z(\CARRYB[25][7] ) );
  ND2P U1927 ( .A(n451), .B(\CARRYB[25][6] ), .Z(n1220) );
  ND2P U1928 ( .A(n451), .B(\SUMB[25][7] ), .Z(n1221) );
  ND2P U1929 ( .A(\CARRYB[25][6] ), .B(\SUMB[25][7] ), .Z(n1222) );
  ND3P U1930 ( .A(n1220), .B(n1221), .C(n1222), .Z(\CARRYB[26][6] ) );
  EO3P U1931 ( .A(\CARRYB[19][8] ), .B(n515), .C(\SUMB[19][9] ), .Z(
        \SUMB[20][8] ) );
  ND2 U1932 ( .A(\CARRYB[19][8] ), .B(\SUMB[19][9] ), .Z(n1223) );
  ND2 U1933 ( .A(\CARRYB[19][8] ), .B(n515), .Z(n1224) );
  ND2 U1934 ( .A(\SUMB[19][9] ), .B(n515), .Z(n1225) );
  ND3P U1935 ( .A(n1223), .B(n1224), .C(n1225), .Z(\CARRYB[20][8] ) );
  ND3 U1936 ( .A(n1442), .B(n1443), .C(n1444), .Z(\CARRYB[42][28] ) );
  EOP U1937 ( .A(\CARRYB[40][11] ), .B(\ab[41][11] ), .Z(n1226) );
  EOP U1938 ( .A(n1226), .B(\SUMB[40][12] ), .Z(\SUMB[41][11] ) );
  ND2 U1939 ( .A(\SUMB[40][12] ), .B(n771), .Z(n1227) );
  ND2 U1940 ( .A(\SUMB[40][12] ), .B(\ab[41][11] ), .Z(n1228) );
  ND2 U1941 ( .A(n771), .B(\ab[41][11] ), .Z(n1229) );
  ND2 U1942 ( .A(n451), .B(\CARRYB[5][26] ), .Z(n1538) );
  EOP U1943 ( .A(\SUMB[30][20] ), .B(\ab[31][19] ), .Z(n1230) );
  ND2 U1944 ( .A(\CARRYB[30][19] ), .B(\SUMB[30][20] ), .Z(n1231) );
  ND2 U1945 ( .A(\CARRYB[30][19] ), .B(\ab[31][19] ), .Z(n1232) );
  ND2 U1946 ( .A(\SUMB[30][20] ), .B(\ab[31][19] ), .Z(n1233) );
  EOP U1947 ( .A(\SUMB[40][14] ), .B(n1234), .Z(\SUMB[41][13] ) );
  ND2 U1948 ( .A(\SUMB[40][14] ), .B(\CARRYB[40][13] ), .Z(n1235) );
  ND2 U1949 ( .A(\SUMB[40][14] ), .B(\ab[41][13] ), .Z(n1236) );
  ND2 U1950 ( .A(\CARRYB[40][13] ), .B(\ab[41][13] ), .Z(n1237) );
  EOP U1951 ( .A(\CARRYB[2][45] ), .B(n2290), .Z(n1238) );
  EOP U1952 ( .A(\SUMB[2][46] ), .B(n1238), .Z(\SUMB[3][45] ) );
  ND2 U1953 ( .A(\SUMB[2][46] ), .B(\CARRYB[2][45] ), .Z(n1239) );
  ND2 U1954 ( .A(\SUMB[2][46] ), .B(n2290), .Z(n1240) );
  ND2 U1955 ( .A(\CARRYB[2][45] ), .B(n2290), .Z(n1241) );
  ND3P U1956 ( .A(n1239), .B(n1240), .C(n1241), .Z(\CARRYB[3][45] ) );
  ND2 U1957 ( .A(\SUMB[3][46] ), .B(\CARRYB[3][45] ), .Z(n1243) );
  ND2 U1958 ( .A(\SUMB[3][46] ), .B(n360), .Z(n1244) );
  ND2 U1959 ( .A(\CARRYB[3][45] ), .B(n360), .Z(n1245) );
  ND3 U1960 ( .A(n1573), .B(n1574), .C(n1575), .Z(\CARRYB[41][19] ) );
  ND2 U1961 ( .A(\SUMB[45][20] ), .B(\CARRYB[45][19] ), .Z(n1247) );
  ND2 U1962 ( .A(\SUMB[45][20] ), .B(\ab[46][19] ), .Z(n1248) );
  ND2 U1963 ( .A(\CARRYB[45][19] ), .B(\ab[46][19] ), .Z(n1249) );
  ND3P U1964 ( .A(n1247), .B(n1248), .C(n1249), .Z(\CARRYB[46][19] ) );
  EOP U1965 ( .A(\CARRYB[23][28] ), .B(\ab[28][24] ), .Z(n1250) );
  ND2 U1966 ( .A(\SUMB[23][29] ), .B(\CARRYB[23][28] ), .Z(n1251) );
  ND2 U1967 ( .A(\SUMB[23][29] ), .B(\ab[28][24] ), .Z(n1252) );
  ND2 U1968 ( .A(\CARRYB[23][28] ), .B(\ab[28][24] ), .Z(n1253) );
  ND3P U1969 ( .A(n1251), .B(n1252), .C(n1253), .Z(\CARRYB[24][28] ) );
  EOP U1970 ( .A(\CARRYB[36][13] ), .B(\ab[37][13] ), .Z(n1254) );
  EOP U1971 ( .A(\SUMB[36][14] ), .B(n1254), .Z(\SUMB[37][13] ) );
  ND2 U1972 ( .A(\SUMB[36][14] ), .B(\CARRYB[36][13] ), .Z(n1255) );
  ND2 U1973 ( .A(\SUMB[36][14] ), .B(\ab[37][13] ), .Z(n1256) );
  ND2 U1974 ( .A(\CARRYB[36][13] ), .B(\ab[37][13] ), .Z(n1257) );
  EOP U1975 ( .A(\CARRYB[34][14] ), .B(\ab[35][14] ), .Z(n1258) );
  ND2 U1976 ( .A(\SUMB[34][15] ), .B(n799), .Z(n1259) );
  ND2 U1977 ( .A(\SUMB[34][15] ), .B(\ab[35][14] ), .Z(n1260) );
  ND2 U1978 ( .A(n799), .B(\ab[35][14] ), .Z(n1261) );
  EOP U1979 ( .A(\SUMB[5][22] ), .B(n1262), .Z(\SUMB[6][21] ) );
  ND2 U1980 ( .A(\SUMB[5][22] ), .B(\CARRYB[5][21] ), .Z(n1263) );
  ND2 U1981 ( .A(\SUMB[5][22] ), .B(n434), .Z(n1264) );
  ND2 U1982 ( .A(\CARRYB[5][21] ), .B(n434), .Z(n1265) );
  EOP U1983 ( .A(\CARRYB[18][10] ), .B(n608), .Z(n1266) );
  EOP U1984 ( .A(\SUMB[18][11] ), .B(n1266), .Z(\SUMB[19][10] ) );
  ND2 U1985 ( .A(\SUMB[18][11] ), .B(\CARRYB[18][10] ), .Z(n1267) );
  ND2 U1986 ( .A(\SUMB[18][11] ), .B(n608), .Z(n1268) );
  ND2 U1987 ( .A(\CARRYB[18][10] ), .B(n608), .Z(n1269) );
  EO3 U1988 ( .A(\CARRYB[31][17] ), .B(\ab[32][17] ), .C(\SUMB[31][18] ), .Z(
        \SUMB[32][17] ) );
  ND2 U1989 ( .A(\CARRYB[31][17] ), .B(\SUMB[31][18] ), .Z(n1270) );
  ND2 U1990 ( .A(\CARRYB[31][17] ), .B(\ab[32][17] ), .Z(n1271) );
  ND2 U1991 ( .A(\SUMB[31][18] ), .B(\ab[32][17] ), .Z(n1272) );
  ND3P U1992 ( .A(n2032), .B(n2033), .C(n2034), .Z(\CARRYB[14][32] ) );
  EO3 U1993 ( .A(\CARRYB[23][37] ), .B(\ab[37][24] ), .C(\SUMB[23][38] ), .Z(
        \SUMB[24][37] ) );
  ND2 U1994 ( .A(\CARRYB[23][37] ), .B(\SUMB[23][38] ), .Z(n1273) );
  ND2 U1995 ( .A(\CARRYB[23][37] ), .B(\ab[37][24] ), .Z(n1274) );
  ND2 U1996 ( .A(\SUMB[23][38] ), .B(\ab[37][24] ), .Z(n1275) );
  IVDA U1997 ( .A(n2246), .Z(n1276) );
  ND2P U1998 ( .A(n1490), .B(n1491), .Z(\SUMB[24][10] ) );
  AN2P U1999 ( .A(n2187), .B(n2193), .Z(\CARRYB[1][16] ) );
  EOP U2000 ( .A(\CARRYB[18][25] ), .B(\ab[25][19] ), .Z(n1277) );
  EOP U2001 ( .A(\SUMB[18][26] ), .B(n1277), .Z(\SUMB[19][25] ) );
  ND2 U2002 ( .A(\SUMB[18][26] ), .B(\CARRYB[18][25] ), .Z(n1278) );
  ND2 U2003 ( .A(\SUMB[18][26] ), .B(\ab[25][19] ), .Z(n1279) );
  ND2 U2004 ( .A(\CARRYB[18][25] ), .B(\ab[25][19] ), .Z(n1280) );
  EOP U2005 ( .A(\CARRYB[22][23] ), .B(n2366), .Z(n1281) );
  ND2 U2006 ( .A(n786), .B(n1283), .Z(n1284) );
  ND2 U2007 ( .A(n1282), .B(n1660), .Z(n1285) );
  ND2P U2008 ( .A(n1284), .B(n1285), .Z(\SUMB[13][25] ) );
  IVDA U2009 ( .A(n786), .Y(n1282) );
  ND2 U2010 ( .A(\SUMB[13][25] ), .B(\CARRYB[13][24] ), .Z(n1287) );
  ND2 U2011 ( .A(\SUMB[13][25] ), .B(n703), .Z(n1288) );
  ND2 U2012 ( .A(\CARRYB[13][24] ), .B(n703), .Z(n1289) );
  ND3P U2013 ( .A(n1287), .B(n1288), .C(n1289), .Z(\CARRYB[14][24] ) );
  EO3 U2014 ( .A(\SUMB[43][9] ), .B(n516), .C(\CARRYB[43][8] ), .Z(
        \SUMB[44][8] ) );
  ND2 U2015 ( .A(\CARRYB[43][8] ), .B(n516), .Z(n1292) );
  ND3P U2016 ( .A(n1290), .B(n1291), .C(n1292), .Z(\CARRYB[44][8] ) );
  EOP U2017 ( .A(\CARRYB[21][15] ), .B(n720), .Z(n1293) );
  EOP U2018 ( .A(\SUMB[21][16] ), .B(n1293), .Z(\SUMB[22][15] ) );
  ND2 U2019 ( .A(\SUMB[21][16] ), .B(\CARRYB[21][15] ), .Z(n1294) );
  ND2 U2020 ( .A(\SUMB[21][16] ), .B(n720), .Z(n1295) );
  ND2 U2021 ( .A(\CARRYB[21][15] ), .B(n720), .Z(n1296) );
  ND3 U2022 ( .A(n1294), .B(n1295), .C(n1296), .Z(\CARRYB[22][15] ) );
  EO3 U2023 ( .A(\CARRYB[9][35] ), .B(n582), .C(\SUMB[9][36] ), .Z(
        \SUMB[10][35] ) );
  ND2 U2024 ( .A(\CARRYB[9][35] ), .B(\SUMB[9][36] ), .Z(n1297) );
  ND2 U2025 ( .A(\CARRYB[9][35] ), .B(n582), .Z(n1298) );
  ND2 U2026 ( .A(\SUMB[9][36] ), .B(n582), .Z(n1299) );
  ND3 U2027 ( .A(n1297), .B(n1298), .C(n1299), .Z(\CARRYB[10][35] ) );
  EO3 U2028 ( .A(\CARRYB[11][34] ), .B(n674), .C(\SUMB[11][35] ), .Z(
        \SUMB[12][34] ) );
  ND2 U2029 ( .A(\CARRYB[11][34] ), .B(\SUMB[11][35] ), .Z(n1300) );
  ND2 U2030 ( .A(\CARRYB[11][34] ), .B(n674), .Z(n1301) );
  ND2 U2031 ( .A(\SUMB[11][35] ), .B(n674), .Z(n1302) );
  ND3 U2032 ( .A(n1300), .B(n1301), .C(n1302), .Z(\CARRYB[12][34] ) );
  EOP U2033 ( .A(\SUMB[19][34] ), .B(\ab[33][20] ), .Z(n1303) );
  EOP U2034 ( .A(\CARRYB[19][33] ), .B(n1303), .Z(\SUMB[20][33] ) );
  EO3P U2035 ( .A(\CARRYB[25][30] ), .B(\ab[30][26] ), .C(\SUMB[25][31] ), .Z(
        \SUMB[26][30] ) );
  ND2 U2036 ( .A(\CARRYB[25][30] ), .B(\SUMB[25][31] ), .Z(n1304) );
  ND2 U2037 ( .A(\CARRYB[25][30] ), .B(\ab[30][26] ), .Z(n1305) );
  ND2 U2038 ( .A(\SUMB[25][31] ), .B(\ab[30][26] ), .Z(n1306) );
  ND3 U2039 ( .A(n1304), .B(n1305), .C(n1306), .Z(\CARRYB[26][30] ) );
  ND3 U2040 ( .A(n1797), .B(n1798), .C(n1799), .Z(\CARRYB[40][10] ) );
  ND2 U2041 ( .A(\CARRYB[30][9] ), .B(n782), .Z(n1558) );
  ND2 U2042 ( .A(n782), .B(n562), .Z(n1560) );
  EO3 U2043 ( .A(\CARRYB[29][25] ), .B(\ab[30][25] ), .C(\SUMB[29][26] ), .Z(
        \SUMB[30][25] ) );
  ND2P U2044 ( .A(\CARRYB[29][25] ), .B(\SUMB[29][26] ), .Z(n1307) );
  ND2P U2045 ( .A(\CARRYB[29][25] ), .B(\ab[30][25] ), .Z(n1308) );
  ND2 U2046 ( .A(\SUMB[29][26] ), .B(\ab[30][25] ), .Z(n1309) );
  ND3P U2047 ( .A(n1307), .B(n1308), .C(n1309), .Z(\CARRYB[30][25] ) );
  EOP U2048 ( .A(\SUMB[14][32] ), .B(\ab[31][15] ), .Z(n1310) );
  EOP U2049 ( .A(\CARRYB[14][31] ), .B(n1310), .Z(\SUMB[15][31] ) );
  ND2 U2050 ( .A(\CARRYB[14][31] ), .B(\SUMB[14][32] ), .Z(n1311) );
  ND2 U2051 ( .A(\CARRYB[14][31] ), .B(\ab[31][15] ), .Z(n1312) );
  ND2 U2052 ( .A(\SUMB[14][32] ), .B(\ab[31][15] ), .Z(n1313) );
  ND3P U2053 ( .A(n1311), .B(n1312), .C(n1313), .Z(\CARRYB[15][31] ) );
  FA1A U2054 ( .A(\ab[33][25] ), .B(\CARRYB[32][25] ), .CI(\SUMB[32][26] ), 
        .CO(n1314) );
  ND2 U2055 ( .A(\CARRYB[15][31] ), .B(\SUMB[15][32] ), .Z(n1413) );
  EO3P U2056 ( .A(\CARRYB[12][2] ), .B(n2266), .C(\SUMB[12][3] ), .Z(
        \SUMB[13][2] ) );
  ND2 U2057 ( .A(\SUMB[40][29] ), .B(\ab[41][28] ), .Z(n1316) );
  ND3P U2058 ( .A(n1315), .B(n1316), .C(n1317), .Z(\CARRYB[41][28] ) );
  ND2 U2059 ( .A(\SUMB[39][18] ), .B(\CARRYB[39][17] ), .Z(n1376) );
  ND2 U2060 ( .A(\SUMB[39][18] ), .B(\ab[40][17] ), .Z(n1377) );
  AN2 U2061 ( .A(\ab[23][23] ), .B(n2117), .Z(n2227) );
  IV U2062 ( .A(n1740), .Z(n1741) );
  EOP U2063 ( .A(\CARRYB[39][5] ), .B(n432), .Z(n1318) );
  EOP U2064 ( .A(\SUMB[39][6] ), .B(n1318), .Z(\SUMB[40][5] ) );
  ND2 U2065 ( .A(\SUMB[39][6] ), .B(\CARRYB[39][5] ), .Z(n1319) );
  ND2 U2066 ( .A(\SUMB[39][6] ), .B(n432), .Z(n1320) );
  ND2 U2067 ( .A(\CARRYB[39][5] ), .B(n432), .Z(n1321) );
  EOP U2068 ( .A(\CARRYB[23][11] ), .B(n621), .Z(n1322) );
  ND2 U2069 ( .A(\SUMB[23][12] ), .B(\CARRYB[23][11] ), .Z(n1323) );
  ND2 U2070 ( .A(\SUMB[23][12] ), .B(n621), .Z(n1324) );
  ND2 U2071 ( .A(\CARRYB[23][11] ), .B(n621), .Z(n1325) );
  ND3 U2072 ( .A(n1323), .B(n1324), .C(n1325), .Z(\CARRYB[24][11] ) );
  IV U2073 ( .A(\CARRYB[9][20] ), .Z(n1740) );
  ND2 U2074 ( .A(\SUMB[42][12] ), .B(\CARRYB[42][11] ), .Z(n1326) );
  ND2 U2075 ( .A(\SUMB[42][12] ), .B(\ab[43][11] ), .Z(n1327) );
  ND2 U2076 ( .A(\CARRYB[42][11] ), .B(\ab[43][11] ), .Z(n1328) );
  ND3 U2077 ( .A(n1326), .B(n1327), .C(n1328), .Z(\CARRYB[43][11] ) );
  EO U2078 ( .A(\CARRYB[40][12] ), .B(\ab[41][12] ), .Z(n1329) );
  EO U2079 ( .A(\SUMB[40][13] ), .B(n1329), .Z(\SUMB[41][12] ) );
  ND2 U2080 ( .A(\SUMB[40][13] ), .B(\CARRYB[40][12] ), .Z(n1330) );
  ND2 U2081 ( .A(\SUMB[40][13] ), .B(\ab[41][12] ), .Z(n1331) );
  ND2 U2082 ( .A(\CARRYB[40][12] ), .B(\ab[41][12] ), .Z(n1332) );
  ND3P U2083 ( .A(n1330), .B(n1331), .C(n1332), .Z(\CARRYB[41][12] ) );
  EO3P U2084 ( .A(\SUMB[1][29] ), .B(n2210), .C(\CARRYB[1][28] ), .Z(
        \SUMB[2][28] ) );
  ND2 U2085 ( .A(\SUMB[1][29] ), .B(\CARRYB[1][28] ), .Z(n1333) );
  ND2 U2086 ( .A(\SUMB[1][29] ), .B(n2210), .Z(n1334) );
  ND2 U2087 ( .A(\CARRYB[1][28] ), .B(n2210), .Z(n1335) );
  EO U2088 ( .A(\SUMB[9][27] ), .B(n1582), .Z(\SUMB[10][26] ) );
  ND2 U2089 ( .A(n569), .B(\CARRYB[36][9] ), .Z(n1337) );
  ND2 U2090 ( .A(n569), .B(\SUMB[36][10] ), .Z(n1338) );
  ND2 U2091 ( .A(\CARRYB[36][9] ), .B(\SUMB[36][10] ), .Z(n1339) );
  ND3P U2092 ( .A(n1337), .B(n1338), .C(n1339), .Z(\CARRYB[37][9] ) );
  ND2 U2093 ( .A(n531), .B(\CARRYB[37][8] ), .Z(n1340) );
  EOP U2094 ( .A(\CARRYB[23][25] ), .B(\ab[25][24] ), .Z(n1343) );
  EOP U2095 ( .A(\SUMB[23][26] ), .B(n1343), .Z(\SUMB[24][25] ) );
  ND2 U2096 ( .A(\SUMB[23][26] ), .B(\CARRYB[23][25] ), .Z(n1344) );
  ND2 U2097 ( .A(\SUMB[23][26] ), .B(\ab[25][24] ), .Z(n1345) );
  ND2 U2098 ( .A(\CARRYB[23][25] ), .B(\ab[25][24] ), .Z(n1346) );
  ND3P U2099 ( .A(n1344), .B(n1345), .C(n1346), .Z(\CARRYB[24][25] ) );
  EO3 U2100 ( .A(\CARRYB[39][11] ), .B(\ab[40][11] ), .C(\SUMB[39][12] ), .Z(
        \SUMB[40][11] ) );
  ND2 U2101 ( .A(\SUMB[39][12] ), .B(\ab[40][11] ), .Z(n1349) );
  AN2 U2102 ( .A(\CARRYB[47][0] ), .B(\SUMB[47][1] ), .Z(\A2[47] ) );
  ND3 U2103 ( .A(n1657), .B(n1658), .C(n1659), .Z(\CARRYB[27][20] ) );
  EOP U2104 ( .A(\CARRYB[2][28] ), .B(n2284), .Z(n1351) );
  EOP U2105 ( .A(\SUMB[2][29] ), .B(n1351), .Z(\SUMB[3][28] ) );
  AN2P U2106 ( .A(A[28]), .B(n2327), .Z(n2284) );
  EOP U2107 ( .A(\CARRYB[38][25] ), .B(\ab[39][25] ), .Z(n1352) );
  EOP U2108 ( .A(\SUMB[38][26] ), .B(n1352), .Z(\SUMB[39][25] ) );
  ND2 U2109 ( .A(\CARRYB[38][25] ), .B(\ab[39][25] ), .Z(n1355) );
  ND3P U2110 ( .A(n1353), .B(n1354), .C(n1355), .Z(\CARRYB[39][25] ) );
  ND2 U2111 ( .A(\SUMB[15][33] ), .B(\CARRYB[15][32] ), .Z(n1356) );
  ND2 U2112 ( .A(\SUMB[15][33] ), .B(\ab[32][16] ), .Z(n1357) );
  ND3 U2113 ( .A(n1356), .B(n1357), .C(n1358), .Z(\CARRYB[16][32] ) );
  EO3 U2114 ( .A(\SUMB[24][30] ), .B(\ab[29][25] ), .C(\CARRYB[24][29] ), .Z(
        \SUMB[25][29] ) );
  ND2P U2115 ( .A(\CARRYB[6][25] ), .B(\SUMB[6][26] ), .Z(n1543) );
  ND2P U2116 ( .A(n467), .B(\SUMB[6][26] ), .Z(n1542) );
  EO3 U2117 ( .A(\CARRYB[41][25] ), .B(\ab[42][25] ), .C(\SUMB[41][26] ), .Z(
        \SUMB[42][25] ) );
  ND2 U2118 ( .A(\CARRYB[41][25] ), .B(\SUMB[41][26] ), .Z(n1359) );
  ND2 U2119 ( .A(\CARRYB[41][25] ), .B(\ab[42][25] ), .Z(n1360) );
  ND2 U2120 ( .A(\SUMB[41][26] ), .B(\ab[42][25] ), .Z(n1361) );
  ND2 U2121 ( .A(\CARRYB[23][31] ), .B(\SUMB[23][32] ), .Z(n1362) );
  ND2 U2122 ( .A(\CARRYB[23][31] ), .B(\ab[31][24] ), .Z(n1363) );
  ND2 U2123 ( .A(\SUMB[23][32] ), .B(\ab[31][24] ), .Z(n1364) );
  ND3 U2124 ( .A(n1362), .B(n1363), .C(n1364), .Z(\CARRYB[24][31] ) );
  ND2 U2125 ( .A(\SUMB[30][8] ), .B(\CARRYB[30][7] ), .Z(n1366) );
  ND2 U2126 ( .A(\SUMB[30][8] ), .B(n469), .Z(n1367) );
  ND2 U2127 ( .A(\CARRYB[30][7] ), .B(n469), .Z(n1368) );
  ND3 U2128 ( .A(n1366), .B(n1367), .C(n1368), .Z(\CARRYB[31][7] ) );
  EOP U2129 ( .A(\SUMB[43][4] ), .B(n2285), .Z(n1369) );
  EOP U2130 ( .A(\CARRYB[43][3] ), .B(n1369), .Z(\SUMB[44][3] ) );
  ND2 U2131 ( .A(\CARRYB[43][3] ), .B(\SUMB[43][4] ), .Z(n1370) );
  ND2 U2132 ( .A(\CARRYB[43][3] ), .B(n2285), .Z(n1371) );
  ND2 U2133 ( .A(\SUMB[43][4] ), .B(n2285), .Z(n1372) );
  ND3P U2134 ( .A(n1370), .B(n1371), .C(n1372), .Z(\CARRYB[44][3] ) );
  ND2 U2135 ( .A(\SUMB[14][13] ), .B(\CARRYB[14][12] ), .Z(n1373) );
  ND2 U2136 ( .A(\SUMB[14][13] ), .B(n655), .Z(n1374) );
  ND2 U2137 ( .A(\CARRYB[14][12] ), .B(n655), .Z(n1375) );
  ND3P U2138 ( .A(n1373), .B(n1374), .C(n1375), .Z(\CARRYB[15][12] ) );
  ND3 U2139 ( .A(n1518), .B(n1519), .C(n1520), .Z(\CARRYB[24][33] ) );
  AN2P U2140 ( .A(\ab[43][43] ), .B(PRODUCT[0]), .Z(n2200) );
  EOP U2141 ( .A(\SUMB[25][16] ), .B(n1782), .Z(\SUMB[26][15] ) );
  ND2P U2142 ( .A(\CARRYB[32][1] ), .B(\SUMB[32][2] ), .Z(n1893) );
  ND2P U2143 ( .A(n2181), .B(\CARRYB[32][1] ), .Z(n1891) );
  EO3 U2144 ( .A(\CARRYB[21][32] ), .B(\ab[32][22] ), .C(\SUMB[21][33] ), .Z(
        \SUMB[22][32] ) );
  ND3P U2145 ( .A(n1376), .B(n1377), .C(n1378), .Z(\CARRYB[40][17] ) );
  ND2P U2146 ( .A(\CARRYB[18][26] ), .B(\SUMB[18][27] ), .Z(n1380) );
  ND2P U2147 ( .A(\CARRYB[18][26] ), .B(\ab[26][19] ), .Z(n1381) );
  ND2 U2148 ( .A(\SUMB[18][27] ), .B(\ab[26][19] ), .Z(n1382) );
  ND3P U2149 ( .A(n1380), .B(n1381), .C(n1382), .Z(\CARRYB[19][26] ) );
  ND2 U2150 ( .A(\CARRYB[26][23] ), .B(\SUMB[26][24] ), .Z(n1686) );
  AN2 U2151 ( .A(n2314), .B(n2312), .Z(\CARRYB[1][32] ) );
  EOP U2152 ( .A(\CARRYB[43][6] ), .B(n453), .Z(n1383) );
  ND2P U2153 ( .A(\SUMB[43][7] ), .B(\CARRYB[43][6] ), .Z(n1384) );
  ND2P U2154 ( .A(\SUMB[43][7] ), .B(n453), .Z(n1385) );
  ND2 U2155 ( .A(\CARRYB[43][6] ), .B(n453), .Z(n1386) );
  ND3P U2156 ( .A(n1384), .B(n1385), .C(n1386), .Z(\CARRYB[44][6] ) );
  EO3P U2157 ( .A(\SUMB[22][15] ), .B(n693), .C(\CARRYB[22][14] ), .Z(
        \SUMB[23][14] ) );
  ND2 U2158 ( .A(\CARRYB[22][14] ), .B(\SUMB[22][15] ), .Z(n1387) );
  ND2 U2159 ( .A(\SUMB[22][15] ), .B(n693), .Z(n1389) );
  ND2 U2160 ( .A(\CARRYB[33][10] ), .B(n590), .Z(n1393) );
  ND2 U2161 ( .A(\SUMB[39][11] ), .B(\CARRYB[39][10] ), .Z(n1797) );
  ND2 U2162 ( .A(\SUMB[39][11] ), .B(n637), .Z(n1798) );
  EOP U2163 ( .A(\CARRYB[32][28] ), .B(\ab[33][28] ), .Z(n1394) );
  ND2 U2164 ( .A(\SUMB[32][29] ), .B(\CARRYB[32][28] ), .Z(n1395) );
  ND2 U2165 ( .A(\SUMB[32][29] ), .B(\ab[33][28] ), .Z(n1396) );
  ND2 U2166 ( .A(\CARRYB[32][28] ), .B(\ab[33][28] ), .Z(n1397) );
  ND2 U2167 ( .A(\SUMB[21][33] ), .B(\ab[32][22] ), .Z(n1399) );
  ND2 U2168 ( .A(\SUMB[19][34] ), .B(\CARRYB[19][33] ), .Z(n1401) );
  ND2 U2169 ( .A(\SUMB[19][34] ), .B(\ab[33][20] ), .Z(n1402) );
  ND2 U2170 ( .A(\CARRYB[19][33] ), .B(\ab[33][20] ), .Z(n1403) );
  ND3 U2171 ( .A(n1401), .B(n1402), .C(n1403), .Z(\CARRYB[20][33] ) );
  EOP U2172 ( .A(\CARRYB[1][42] ), .B(n2265), .Z(n1404) );
  AN2P U2173 ( .A(n2220), .B(n2224), .Z(\CARRYB[1][26] ) );
  ND3 U2174 ( .A(n2050), .B(n2051), .C(n2052), .Z(\CARRYB[25][1] ) );
  EOP U2175 ( .A(\CARRYB[21][28] ), .B(\ab[28][22] ), .Z(n1405) );
  EOP U2176 ( .A(\SUMB[21][29] ), .B(n1405), .Z(\SUMB[22][28] ) );
  ND2 U2177 ( .A(\CARRYB[21][28] ), .B(\ab[28][22] ), .Z(n1408) );
  ND2 U2178 ( .A(\CARRYB[22][28] ), .B(\SUMB[22][29] ), .Z(n1409) );
  ND2 U2179 ( .A(\CARRYB[22][28] ), .B(\ab[28][23] ), .Z(n1410) );
  ND2 U2180 ( .A(\SUMB[22][29] ), .B(\ab[28][23] ), .Z(n1411) );
  ND3P U2181 ( .A(n1409), .B(n1410), .C(n1411), .Z(\CARRYB[23][28] ) );
  ND2 U2182 ( .A(\SUMB[15][32] ), .B(\ab[31][16] ), .Z(n1415) );
  ND3 U2183 ( .A(n1704), .B(n1705), .C(n1706), .Z(\CARRYB[45][3] ) );
  EO3P U2184 ( .A(\CARRYB[4][37] ), .B(n397), .C(\SUMB[4][38] ), .Z(
        \SUMB[5][37] ) );
  ND2 U2185 ( .A(\CARRYB[4][37] ), .B(\SUMB[4][38] ), .Z(n1416) );
  ND2 U2186 ( .A(\CARRYB[4][37] ), .B(n397), .Z(n1417) );
  ND2 U2187 ( .A(\SUMB[4][38] ), .B(n397), .Z(n1418) );
  ND3 U2188 ( .A(n1416), .B(n1417), .C(n1418), .Z(\CARRYB[5][37] ) );
  EO3P U2189 ( .A(\SUMB[11][34] ), .B(n653), .C(\CARRYB[11][33] ), .Z(
        \SUMB[12][33] ) );
  ND2P U2190 ( .A(\CARRYB[11][33] ), .B(n653), .Z(n1421) );
  ND3P U2191 ( .A(n1419), .B(n1420), .C(n1421), .Z(\CARRYB[12][33] ) );
  ND2 U2192 ( .A(\CARRYB[26][20] ), .B(\ab[27][20] ), .Z(n1658) );
  EO3P U2193 ( .A(\CARRYB[42][7] ), .B(n474), .C(\SUMB[42][8] ), .Z(
        \SUMB[43][7] ) );
  ND2 U2194 ( .A(\CARRYB[42][7] ), .B(\SUMB[42][8] ), .Z(n1422) );
  ND2 U2195 ( .A(\CARRYB[42][7] ), .B(n474), .Z(n1423) );
  ND2 U2196 ( .A(\SUMB[42][8] ), .B(n474), .Z(n1424) );
  ND3 U2197 ( .A(n1422), .B(n1423), .C(n1424), .Z(\CARRYB[43][7] ) );
  ND2 U2198 ( .A(\CARRYB[45][18] ), .B(\ab[46][18] ), .Z(n1428) );
  ND3P U2199 ( .A(n1426), .B(n1427), .C(n1428), .Z(\CARRYB[46][18] ) );
  EOP U2200 ( .A(\CARRYB[35][21] ), .B(\ab[36][21] ), .Z(n1429) );
  EOP U2201 ( .A(n1429), .B(\SUMB[35][22] ), .Z(\SUMB[36][21] ) );
  ND2 U2202 ( .A(\SUMB[35][22] ), .B(\CARRYB[35][21] ), .Z(n1430) );
  ND2 U2203 ( .A(\SUMB[35][22] ), .B(\ab[36][21] ), .Z(n1431) );
  ND2 U2204 ( .A(\CARRYB[35][21] ), .B(\ab[36][21] ), .Z(n1432) );
  ND3 U2205 ( .A(n1430), .B(n1431), .C(n1432), .Z(\CARRYB[36][21] ) );
  EOP U2206 ( .A(\SUMB[28][25] ), .B(n1433), .Z(\SUMB[29][24] ) );
  ND2 U2207 ( .A(\SUMB[28][25] ), .B(\CARRYB[28][24] ), .Z(n1434) );
  ND2 U2208 ( .A(\SUMB[28][25] ), .B(\ab[29][24] ), .Z(n1435) );
  ND2 U2209 ( .A(\CARRYB[28][24] ), .B(\ab[29][24] ), .Z(n1436) );
  ND3 U2210 ( .A(n1434), .B(n1435), .C(n1436), .Z(\CARRYB[29][24] ) );
  EOP U2211 ( .A(\CARRYB[17][38] ), .B(\ab[38][18] ), .Z(n1437) );
  EOP U2212 ( .A(\SUMB[17][39] ), .B(n1437), .Z(\SUMB[18][38] ) );
  ND2 U2213 ( .A(\SUMB[17][39] ), .B(\CARRYB[17][38] ), .Z(n1438) );
  ND2 U2214 ( .A(\SUMB[17][39] ), .B(\ab[38][18] ), .Z(n1439) );
  ND2 U2215 ( .A(\CARRYB[17][38] ), .B(\ab[38][18] ), .Z(n1440) );
  EOP U2216 ( .A(\CARRYB[41][28] ), .B(\ab[42][28] ), .Z(n1441) );
  EOP U2217 ( .A(\SUMB[41][29] ), .B(n1441), .Z(\SUMB[42][28] ) );
  ND2 U2218 ( .A(\SUMB[41][29] ), .B(\CARRYB[41][28] ), .Z(n1442) );
  ND2 U2219 ( .A(\SUMB[41][29] ), .B(\ab[42][28] ), .Z(n1443) );
  ND3P U2220 ( .A(n1996), .B(n1997), .C(n1998), .Z(\CARRYB[11][13] ) );
  ND2 U2221 ( .A(\SUMB[45][6] ), .B(\CARRYB[45][5] ), .Z(n1445) );
  ND2 U2222 ( .A(\SUMB[45][6] ), .B(n305), .Z(n1446) );
  ND2 U2223 ( .A(\CARRYB[45][5] ), .B(n305), .Z(n1447) );
  AN2 U2224 ( .A(n2188), .B(n2172), .Z(\CARRYB[1][35] ) );
  ND2 U2225 ( .A(\SUMB[42][30] ), .B(\CARRYB[42][29] ), .Z(n1449) );
  ND2 U2226 ( .A(\SUMB[42][30] ), .B(\ab[43][29] ), .Z(n1450) );
  ND2 U2227 ( .A(\CARRYB[42][29] ), .B(\ab[43][29] ), .Z(n1451) );
  EOP U2228 ( .A(\CARRYB[25][37] ), .B(\ab[37][26] ), .Z(n1452) );
  EOP U2229 ( .A(\SUMB[25][38] ), .B(n1452), .Z(\SUMB[26][37] ) );
  ND2 U2230 ( .A(\SUMB[25][38] ), .B(\CARRYB[25][37] ), .Z(n1453) );
  ND2 U2231 ( .A(\SUMB[25][38] ), .B(\ab[37][26] ), .Z(n1454) );
  ND2 U2232 ( .A(\CARRYB[25][37] ), .B(\ab[37][26] ), .Z(n1455) );
  ND3P U2233 ( .A(n1453), .B(n1454), .C(n1455), .Z(\CARRYB[26][37] ) );
  ND2 U2234 ( .A(\SUMB[1][45] ), .B(n891), .Z(n1457) );
  ND2 U2235 ( .A(\SUMB[1][45] ), .B(n2248), .Z(n1458) );
  ND2 U2236 ( .A(n891), .B(n2248), .Z(n1459) );
  EOP U2237 ( .A(\SUMB[20][40] ), .B(\ab[39][21] ), .Z(n1460) );
  EOP U2238 ( .A(\CARRYB[20][39] ), .B(n1460), .Z(\SUMB[21][39] ) );
  ND2 U2239 ( .A(\CARRYB[20][39] ), .B(\SUMB[20][40] ), .Z(n1461) );
  ND2 U2240 ( .A(\CARRYB[20][39] ), .B(\ab[39][21] ), .Z(n1462) );
  ND2 U2241 ( .A(\SUMB[20][40] ), .B(\ab[39][21] ), .Z(n1463) );
  ND2 U2242 ( .A(\SUMB[12][27] ), .B(n680), .Z(n1465) );
  EO3 U2243 ( .A(\SUMB[26][23] ), .B(\ab[27][22] ), .C(\CARRYB[26][22] ), .Z(
        \SUMB[27][22] ) );
  ND2 U2244 ( .A(\CARRYB[26][22] ), .B(\SUMB[26][23] ), .Z(n1467) );
  ND2 U2245 ( .A(\CARRYB[26][22] ), .B(\ab[27][22] ), .Z(n1468) );
  ND2 U2246 ( .A(\SUMB[26][23] ), .B(\ab[27][22] ), .Z(n1469) );
  ND3 U2247 ( .A(n1467), .B(n1468), .C(n1469), .Z(\CARRYB[27][22] ) );
  ND3 U2248 ( .A(n1694), .B(n1695), .C(n1696), .Z(\CARRYB[14][13] ) );
  ND2 U2249 ( .A(\CARRYB[5][29] ), .B(\SUMB[5][30] ), .Z(n2036) );
  ND2 U2250 ( .A(\CARRYB[5][29] ), .B(n455), .Z(n2037) );
  EO U2251 ( .A(\CARRYB[9][17] ), .B(n600), .Z(n1470) );
  EO U2252 ( .A(\SUMB[9][18] ), .B(n1470), .Z(\SUMB[10][17] ) );
  ND2 U2253 ( .A(\SUMB[9][18] ), .B(\CARRYB[9][17] ), .Z(n1471) );
  ND2 U2254 ( .A(\SUMB[9][18] ), .B(n600), .Z(n1472) );
  ND2 U2255 ( .A(\CARRYB[9][17] ), .B(n600), .Z(n1473) );
  FA1AP U2256 ( .A(\CARRYB[44][5] ), .B(n394), .CI(\SUMB[44][6] ), .CO(n876), 
        .S(n1474) );
  EOP U2257 ( .A(\CARRYB[27][26] ), .B(\ab[28][26] ), .Z(n1475) );
  EOP U2258 ( .A(\SUMB[27][27] ), .B(n1475), .Z(\SUMB[28][26] ) );
  ND2 U2259 ( .A(\SUMB[27][27] ), .B(\CARRYB[27][26] ), .Z(n1476) );
  ND2 U2260 ( .A(\SUMB[27][27] ), .B(\ab[28][26] ), .Z(n1477) );
  ND2 U2261 ( .A(\CARRYB[27][26] ), .B(\ab[28][26] ), .Z(n1478) );
  EO3P U2262 ( .A(\CARRYB[33][25] ), .B(\ab[34][25] ), .C(\SUMB[33][26] ), .Z(
        \SUMB[34][25] ) );
  ND2 U2263 ( .A(\SUMB[33][26] ), .B(\ab[34][25] ), .Z(n1481) );
  AN2 U2264 ( .A(n2167), .B(n2170), .Z(\CARRYB[1][30] ) );
  EO3 U2265 ( .A(\CARRYB[43][24] ), .B(\ab[44][24] ), .C(\SUMB[43][25] ), .Z(
        \SUMB[44][24] ) );
  ND2 U2266 ( .A(\CARRYB[43][24] ), .B(\SUMB[43][25] ), .Z(n1482) );
  ND2 U2267 ( .A(\CARRYB[43][24] ), .B(\ab[44][24] ), .Z(n1483) );
  ND2 U2268 ( .A(\SUMB[43][25] ), .B(\ab[44][24] ), .Z(n1484) );
  ND3P U2269 ( .A(n1482), .B(n1483), .C(n1484), .Z(\CARRYB[44][24] ) );
  EOP U2270 ( .A(\CARRYB[6][35] ), .B(n450), .Z(n1485) );
  ND2 U2271 ( .A(\SUMB[6][36] ), .B(\CARRYB[6][35] ), .Z(n1486) );
  ND2 U2272 ( .A(\SUMB[6][36] ), .B(n450), .Z(n1487) );
  ND2 U2273 ( .A(\CARRYB[6][35] ), .B(n450), .Z(n1488) );
  ND2 U2274 ( .A(\SUMB[3][31] ), .B(\CARRYB[3][30] ), .Z(n2069) );
  EOP U2275 ( .A(n2066), .B(\CARRYB[3][30] ), .Z(\SUMB[4][30] ) );
  ND3P U2276 ( .A(n2063), .B(n2064), .C(n2065), .Z(\CARRYB[3][30] ) );
  EO3 U2277 ( .A(\CARRYB[41][26] ), .B(\ab[42][26] ), .C(\SUMB[41][27] ), .Z(
        \SUMB[42][26] ) );
  ND2 U2278 ( .A(\CARRYB[41][26] ), .B(\SUMB[41][27] ), .Z(n1492) );
  ND2 U2279 ( .A(\CARRYB[41][26] ), .B(\ab[42][26] ), .Z(n1493) );
  ND2 U2280 ( .A(\SUMB[41][27] ), .B(\ab[42][26] ), .Z(n1494) );
  ND3P U2281 ( .A(n1492), .B(n1493), .C(n1494), .Z(\CARRYB[42][26] ) );
  EO3P U2282 ( .A(n2181), .B(\CARRYB[32][1] ), .C(\SUMB[32][2] ), .Z(
        \SUMB[33][1] ) );
  ND3 U2283 ( .A(n1746), .B(n1747), .C(n1748), .Z(\CARRYB[12][14] ) );
  ND3 U2284 ( .A(n2008), .B(n2009), .C(n2010), .Z(\CARRYB[3][28] ) );
  EO3 U2285 ( .A(\SUMB[21][34] ), .B(\ab[33][22] ), .C(\CARRYB[21][33] ), .Z(
        \SUMB[22][33] ) );
  ND2 U2286 ( .A(\SUMB[21][34] ), .B(\CARRYB[21][33] ), .Z(n1495) );
  ND2 U2287 ( .A(\SUMB[21][34] ), .B(\ab[33][22] ), .Z(n1496) );
  ND2 U2288 ( .A(\CARRYB[21][33] ), .B(\ab[33][22] ), .Z(n1497) );
  ND3 U2289 ( .A(n1495), .B(n1496), .C(n1497), .Z(\CARRYB[22][33] ) );
  ND2 U2290 ( .A(\SUMB[13][22] ), .B(n1499), .Z(n1500) );
  ND2 U2291 ( .A(n1498), .B(n1502), .Z(n1501) );
  IVDA U2292 ( .A(\SUMB[13][22] ), .Y(n1498) );
  IV U2293 ( .A(n1502), .Z(n1499) );
  EOP U2294 ( .A(\CARRYB[13][21] ), .B(n704), .Z(n1502) );
  ND2 U2295 ( .A(\SUMB[13][22] ), .B(\CARRYB[13][21] ), .Z(n1503) );
  ND2 U2296 ( .A(\SUMB[13][22] ), .B(n704), .Z(n1504) );
  ND2 U2297 ( .A(\CARRYB[13][21] ), .B(n704), .Z(n1505) );
  ND3 U2298 ( .A(n1807), .B(n1808), .C(n1809), .Z(\CARRYB[3][18] ) );
  EOP U2299 ( .A(\SUMB[35][36] ), .B(\ab[36][35] ), .Z(n1506) );
  EOP U2300 ( .A(\CARRYB[35][35] ), .B(n1506), .Z(\SUMB[36][35] ) );
  ND2 U2301 ( .A(\CARRYB[35][35] ), .B(\SUMB[35][36] ), .Z(n1507) );
  ND2 U2302 ( .A(\CARRYB[35][35] ), .B(\ab[36][35] ), .Z(n1508) );
  ND2 U2303 ( .A(\SUMB[35][36] ), .B(\ab[36][35] ), .Z(n1509) );
  ND3P U2304 ( .A(n1507), .B(n1508), .C(n1509), .Z(\CARRYB[36][35] ) );
  ND2 U2305 ( .A(\CARRYB[45][29] ), .B(\ab[46][29] ), .Z(n1513) );
  ND2 U2306 ( .A(\CARRYB[29][10] ), .B(\SUMB[29][11] ), .Z(n1514) );
  ND2 U2307 ( .A(\CARRYB[29][10] ), .B(n580), .Z(n1515) );
  ND2 U2308 ( .A(\SUMB[29][11] ), .B(n580), .Z(n1516) );
  ND3 U2309 ( .A(n1672), .B(n1673), .C(n1674), .Z(\CARRYB[20][32] ) );
  ND2 U2310 ( .A(n451), .B(\SUMB[5][27] ), .Z(n1539) );
  ND2 U2311 ( .A(\CARRYB[5][26] ), .B(\SUMB[5][27] ), .Z(n1540) );
  EOP U2312 ( .A(\CARRYB[23][33] ), .B(\ab[33][24] ), .Z(n1517) );
  EOP U2313 ( .A(\SUMB[23][34] ), .B(n1517), .Z(\SUMB[24][33] ) );
  ND2 U2314 ( .A(\SUMB[23][34] ), .B(\CARRYB[23][33] ), .Z(n1518) );
  ND2 U2315 ( .A(\SUMB[23][34] ), .B(\ab[33][24] ), .Z(n1519) );
  ND2 U2316 ( .A(\CARRYB[23][33] ), .B(\ab[33][24] ), .Z(n1520) );
  EOP U2317 ( .A(\CARRYB[7][28] ), .B(n530), .Z(n1521) );
  EOP U2318 ( .A(\SUMB[7][29] ), .B(n1521), .Z(\SUMB[8][28] ) );
  ND2 U2319 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Z(n1522) );
  ND2 U2320 ( .A(\SUMB[7][29] ), .B(n530), .Z(n1523) );
  ND2 U2321 ( .A(\CARRYB[7][28] ), .B(n530), .Z(n1524) );
  ND3P U2322 ( .A(n1522), .B(n1523), .C(n1524), .Z(\CARRYB[8][28] ) );
  EOP U2323 ( .A(\SUMB[26][14] ), .B(n1525), .Z(\SUMB[27][13] ) );
  ND2 U2324 ( .A(\SUMB[26][14] ), .B(\CARRYB[26][13] ), .Z(n1526) );
  ND2 U2325 ( .A(\SUMB[26][14] ), .B(n682), .Z(n1527) );
  ND2 U2326 ( .A(\CARRYB[26][13] ), .B(n682), .Z(n1528) );
  ND3 U2327 ( .A(n1526), .B(n1527), .C(n1528), .Z(\CARRYB[27][13] ) );
  EOP U2328 ( .A(\CARRYB[5][25] ), .B(n430), .Z(n1529) );
  EOP U2329 ( .A(\SUMB[5][26] ), .B(n1529), .Z(\SUMB[6][25] ) );
  ND2P U2330 ( .A(\SUMB[5][26] ), .B(n430), .Z(n1531) );
  ND2 U2331 ( .A(\CARRYB[5][25] ), .B(n430), .Z(n1532) );
  ND3P U2332 ( .A(n1530), .B(n1531), .C(n1532), .Z(\CARRYB[6][25] ) );
  EOP U2333 ( .A(\CARRYB[30][12] ), .B(n673), .Z(n1533) );
  ND2 U2334 ( .A(\SUMB[30][13] ), .B(\CARRYB[30][12] ), .Z(n1534) );
  ND2 U2335 ( .A(\SUMB[30][13] ), .B(n673), .Z(n1535) );
  ND2 U2336 ( .A(\CARRYB[30][12] ), .B(n673), .Z(n1536) );
  ND3 U2337 ( .A(n1534), .B(n1535), .C(n1536), .Z(\CARRYB[31][12] ) );
  EO3P U2338 ( .A(n451), .B(\CARRYB[5][26] ), .C(\SUMB[5][27] ), .Z(
        \SUMB[6][26] ) );
  EOP U2339 ( .A(\CARRYB[6][25] ), .B(n467), .Z(n1537) );
  ND2 U2340 ( .A(n467), .B(\CARRYB[6][25] ), .Z(n1541) );
  ND3P U2341 ( .A(n1541), .B(n1542), .C(n1543), .Z(\CARRYB[7][25] ) );
  EO3P U2342 ( .A(\CARRYB[41][10] ), .B(\ab[42][10] ), .C(\SUMB[41][11] ), .Z(
        \SUMB[42][10] ) );
  ND2 U2343 ( .A(\CARRYB[41][10] ), .B(\SUMB[41][11] ), .Z(n1544) );
  ND2 U2344 ( .A(\CARRYB[41][10] ), .B(\ab[42][10] ), .Z(n1545) );
  ND2 U2345 ( .A(\SUMB[41][11] ), .B(\ab[42][10] ), .Z(n1546) );
  ND3P U2346 ( .A(n1544), .B(n1545), .C(n1546), .Z(\CARRYB[42][10] ) );
  ND2 U2347 ( .A(\ab[26][20] ), .B(\CARRYB[19][26] ), .Z(n1548) );
  ND2 U2348 ( .A(\ab[26][20] ), .B(\SUMB[19][27] ), .Z(n1549) );
  ND2 U2349 ( .A(\CARRYB[19][26] ), .B(\SUMB[19][27] ), .Z(n1550) );
  ND3P U2350 ( .A(n1551), .B(n1552), .C(n1553), .Z(\CARRYB[21][25] ) );
  EO3 U2351 ( .A(\SUMB[3][32] ), .B(n2304), .C(\CARRYB[3][31] ), .Z(
        \SUMB[4][31] ) );
  ND2 U2352 ( .A(\CARRYB[3][31] ), .B(\SUMB[3][32] ), .Z(n1554) );
  ND2 U2353 ( .A(\CARRYB[3][31] ), .B(n2304), .Z(n1555) );
  ND2 U2354 ( .A(\SUMB[3][32] ), .B(n2304), .Z(n1556) );
  ND3 U2355 ( .A(n1554), .B(n1555), .C(n1556), .Z(\CARRYB[4][31] ) );
  EOP U2356 ( .A(n782), .B(n562), .Z(n1557) );
  EOP U2357 ( .A(\CARRYB[30][9] ), .B(n1557), .Z(\SUMB[31][9] ) );
  EOP U2358 ( .A(\CARRYB[17][10] ), .B(n602), .Z(n1561) );
  ND2 U2359 ( .A(\SUMB[17][11] ), .B(\CARRYB[17][10] ), .Z(n1562) );
  ND2 U2360 ( .A(\SUMB[17][11] ), .B(n602), .Z(n1563) );
  ND2 U2361 ( .A(\CARRYB[17][10] ), .B(n602), .Z(n1564) );
  ND3P U2362 ( .A(n1562), .B(n1563), .C(n1564), .Z(\CARRYB[18][10] ) );
  AN2P U2363 ( .A(\ab[17][17] ), .B(n2117), .Z(n2193) );
  EO3P U2364 ( .A(\SUMB[1][35] ), .B(\CARRYB[1][34] ), .C(n2213), .Z(
        \SUMB[2][34] ) );
  EOP U2365 ( .A(n2275), .B(\CARRYB[2][33] ), .Z(n1565) );
  EOP U2366 ( .A(n1565), .B(\SUMB[2][34] ), .Z(\SUMB[3][33] ) );
  ND2 U2367 ( .A(\SUMB[1][35] ), .B(\CARRYB[1][34] ), .Z(n1566) );
  ND2 U2368 ( .A(\SUMB[1][35] ), .B(n2213), .Z(n1567) );
  ND2 U2369 ( .A(\CARRYB[1][34] ), .B(n2213), .Z(n1568) );
  ND2 U2370 ( .A(n2275), .B(\CARRYB[2][33] ), .Z(n1569) );
  ND2 U2371 ( .A(n2275), .B(\SUMB[2][34] ), .Z(n1570) );
  ND2 U2372 ( .A(\CARRYB[2][33] ), .B(\SUMB[2][34] ), .Z(n1571) );
  ND3P U2373 ( .A(n1569), .B(n1570), .C(n1571), .Z(\CARRYB[3][33] ) );
  EOP U2374 ( .A(\CARRYB[40][19] ), .B(\ab[41][19] ), .Z(n1572) );
  ND2 U2375 ( .A(\SUMB[40][20] ), .B(\CARRYB[40][19] ), .Z(n1573) );
  ND2 U2376 ( .A(\SUMB[40][20] ), .B(\ab[41][19] ), .Z(n1574) );
  ND2 U2377 ( .A(\CARRYB[40][19] ), .B(\ab[41][19] ), .Z(n1575) );
  EO3P U2378 ( .A(\CARRYB[36][19] ), .B(\ab[37][19] ), .C(\SUMB[36][20] ), .Z(
        \SUMB[37][19] ) );
  ND2 U2379 ( .A(\CARRYB[36][19] ), .B(\SUMB[36][20] ), .Z(n1576) );
  ND2 U2380 ( .A(\SUMB[36][20] ), .B(\ab[37][19] ), .Z(n1578) );
  EO3P U2381 ( .A(\CARRYB[25][24] ), .B(\ab[26][24] ), .C(\SUMB[25][25] ), .Z(
        \SUMB[26][24] ) );
  ND2 U2382 ( .A(\CARRYB[25][24] ), .B(\SUMB[25][25] ), .Z(n1579) );
  ND2 U2383 ( .A(\SUMB[25][25] ), .B(\ab[26][24] ), .Z(n1581) );
  ND3P U2384 ( .A(n1579), .B(n1580), .C(n1581), .Z(\CARRYB[26][24] ) );
  EO3P U2385 ( .A(\CARRYB[36][33] ), .B(\ab[37][33] ), .C(\SUMB[36][34] ), .Z(
        \SUMB[37][33] ) );
  EOP U2386 ( .A(n320), .B(n2197), .Z(\SUMB[1][36] ) );
  ND3 U2387 ( .A(n2107), .B(n2108), .C(n2109), .Z(\CARRYB[18][8] ) );
  ND2 U2388 ( .A(\SUMB[9][27] ), .B(\CARRYB[9][26] ), .Z(n1583) );
  ND2 U2389 ( .A(\SUMB[9][27] ), .B(n604), .Z(n1584) );
  ND2 U2390 ( .A(\CARRYB[9][26] ), .B(n604), .Z(n1585) );
  ND3 U2391 ( .A(n1583), .B(n1584), .C(n1585), .Z(\CARRYB[10][26] ) );
  ND2P U2392 ( .A(\CARRYB[4][21] ), .B(n395), .Z(n1813) );
  ND2P U2393 ( .A(\CARRYB[3][16] ), .B(\SUMB[3][17] ), .Z(n1771) );
  EOP U2394 ( .A(n2246), .B(n2196), .Z(\SUMB[1][46] ) );
  EOP U2395 ( .A(\CARRYB[2][22] ), .B(n2292), .Z(n1586) );
  EOP U2396 ( .A(\SUMB[2][23] ), .B(n1586), .Z(\SUMB[3][22] ) );
  ND2 U2397 ( .A(\SUMB[2][23] ), .B(\CARRYB[2][22] ), .Z(n1587) );
  ND2 U2398 ( .A(\SUMB[2][23] ), .B(n2292), .Z(n1588) );
  ND2 U2399 ( .A(\CARRYB[2][22] ), .B(n2292), .Z(n1589) );
  ND3 U2400 ( .A(n1587), .B(n1588), .C(n1589), .Z(\CARRYB[3][22] ) );
  EOP U2401 ( .A(\CARRYB[32][11] ), .B(n636), .Z(n1590) );
  EOP U2402 ( .A(\SUMB[32][12] ), .B(n1590), .Z(\SUMB[33][11] ) );
  ND2 U2403 ( .A(\SUMB[32][12] ), .B(\CARRYB[32][11] ), .Z(n1591) );
  ND2 U2404 ( .A(\SUMB[32][12] ), .B(n636), .Z(n1592) );
  ND2 U2405 ( .A(\CARRYB[32][11] ), .B(n636), .Z(n1593) );
  EO3P U2406 ( .A(n401), .B(\CARRYB[4][33] ), .C(\SUMB[4][34] ), .Z(
        \SUMB[5][33] ) );
  EOP U2407 ( .A(n435), .B(\CARRYB[5][32] ), .Z(n1594) );
  EOP U2408 ( .A(n1594), .B(\SUMB[5][33] ), .Z(\SUMB[6][32] ) );
  ND2 U2409 ( .A(n401), .B(\CARRYB[4][33] ), .Z(n1595) );
  ND2 U2410 ( .A(n401), .B(\SUMB[4][34] ), .Z(n1596) );
  ND2 U2411 ( .A(\CARRYB[4][33] ), .B(\SUMB[4][34] ), .Z(n1597) );
  ND3 U2412 ( .A(n1595), .B(n1596), .C(n1597), .Z(\CARRYB[5][33] ) );
  ND2 U2413 ( .A(n435), .B(\CARRYB[5][32] ), .Z(n1598) );
  ND3P U2414 ( .A(n1598), .B(n1599), .C(n1600), .Z(\CARRYB[6][32] ) );
  EO3 U2415 ( .A(\CARRYB[9][32] ), .B(n598), .C(\SUMB[9][33] ), .Z(
        \SUMB[10][32] ) );
  ND2 U2416 ( .A(\CARRYB[9][32] ), .B(\SUMB[9][33] ), .Z(n1601) );
  ND2 U2417 ( .A(\CARRYB[9][32] ), .B(n598), .Z(n1602) );
  ND2 U2418 ( .A(\SUMB[9][33] ), .B(n598), .Z(n1603) );
  ND3P U2419 ( .A(n1601), .B(n1602), .C(n1603), .Z(\CARRYB[10][32] ) );
  EOP U2420 ( .A(\SUMB[4][28] ), .B(n381), .Z(n1604) );
  EOP U2421 ( .A(\CARRYB[4][27] ), .B(n1604), .Z(\SUMB[5][27] ) );
  ND2P U2422 ( .A(\CARRYB[4][27] ), .B(n381), .Z(n1606) );
  ND2 U2423 ( .A(\SUMB[4][28] ), .B(n381), .Z(n1607) );
  ND3 U2424 ( .A(n1815), .B(n1816), .C(n1817), .Z(\CARRYB[42][4] ) );
  ND2 U2425 ( .A(\SUMB[41][5] ), .B(\CARRYB[41][4] ), .Z(n1815) );
  ND2 U2426 ( .A(\CARRYB[22][23] ), .B(\SUMB[22][24] ), .Z(n1608) );
  ND2 U2427 ( .A(\CARRYB[22][23] ), .B(n2366), .Z(n1609) );
  ND2 U2428 ( .A(\SUMB[22][24] ), .B(n2366), .Z(n1610) );
  ND3P U2429 ( .A(n1608), .B(n1609), .C(n1610), .Z(\CARRYB[23][23] ) );
  EO3 U2430 ( .A(\SUMB[26][22] ), .B(\ab[27][21] ), .C(\CARRYB[26][21] ), .Z(
        \SUMB[27][21] ) );
  EO3P U2431 ( .A(\CARRYB[8][34] ), .B(n555), .C(\SUMB[8][35] ), .Z(
        \SUMB[9][34] ) );
  ND2 U2432 ( .A(\CARRYB[8][34] ), .B(\SUMB[8][35] ), .Z(n1611) );
  ND2 U2433 ( .A(\CARRYB[8][34] ), .B(n555), .Z(n1612) );
  ND2 U2434 ( .A(\SUMB[8][35] ), .B(n555), .Z(n1613) );
  ND3 U2435 ( .A(n1611), .B(n1612), .C(n1613), .Z(\CARRYB[9][34] ) );
  EOP U2436 ( .A(\SUMB[3][45] ), .B(n382), .Z(n1614) );
  EOP U2437 ( .A(\CARRYB[3][44] ), .B(n1614), .Z(\SUMB[4][44] ) );
  ND2P U2438 ( .A(\CARRYB[3][44] ), .B(n382), .Z(n1616) );
  ND2 U2439 ( .A(\SUMB[3][45] ), .B(n382), .Z(n1617) );
  ND2P U2440 ( .A(n2281), .B(\CARRYB[3][30] ), .Z(n2068) );
  EO3 U2441 ( .A(\CARRYB[22][24] ), .B(\ab[24][23] ), .C(\SUMB[22][25] ), .Z(
        \SUMB[23][24] ) );
  ND2 U2442 ( .A(\CARRYB[22][24] ), .B(\SUMB[22][25] ), .Z(n1618) );
  ND2 U2443 ( .A(\CARRYB[22][24] ), .B(\ab[24][23] ), .Z(n1619) );
  ND2 U2444 ( .A(\SUMB[22][25] ), .B(\ab[24][23] ), .Z(n1620) );
  NR2P U2445 ( .A(n2391), .B(n2318), .Z(n1621) );
  NR2 U2446 ( .A(n2391), .B(n2318), .Z(n2314) );
  EOP U2447 ( .A(\CARRYB[29][26] ), .B(\ab[30][26] ), .Z(n1622) );
  EOP U2448 ( .A(\SUMB[29][27] ), .B(n1622), .Z(\SUMB[30][26] ) );
  ND2 U2449 ( .A(\SUMB[29][27] ), .B(\CARRYB[29][26] ), .Z(n1623) );
  ND2 U2450 ( .A(\SUMB[29][27] ), .B(\ab[30][26] ), .Z(n1624) );
  ND2 U2451 ( .A(\CARRYB[29][26] ), .B(\ab[30][26] ), .Z(n1625) );
  ND3 U2452 ( .A(n1858), .B(n1859), .C(n1860), .Z(\CARRYB[39][4] ) );
  EOP U2453 ( .A(\CARRYB[17][8] ), .B(n519), .Z(n1926) );
  ND3P U2454 ( .A(n1931), .B(n1932), .C(n1933), .Z(\CARRYB[21][6] ) );
  EO3P U2455 ( .A(\CARRYB[34][5] ), .B(n374), .C(\SUMB[34][6] ), .Z(
        \SUMB[35][5] ) );
  EO3P U2456 ( .A(\CARRYB[38][18] ), .B(\ab[39][18] ), .C(\SUMB[38][19] ), .Z(
        \SUMB[39][18] ) );
  ND2 U2457 ( .A(\CARRYB[38][18] ), .B(\SUMB[38][19] ), .Z(n1626) );
  ND2 U2458 ( .A(\CARRYB[38][18] ), .B(\ab[39][18] ), .Z(n1627) );
  ND2 U2459 ( .A(\SUMB[38][19] ), .B(\ab[39][18] ), .Z(n1628) );
  EOP U2460 ( .A(n2224), .B(n2220), .Z(\SUMB[1][26] ) );
  EOP U2461 ( .A(\CARRYB[43][18] ), .B(\ab[44][18] ), .Z(n1629) );
  EOP U2462 ( .A(\SUMB[43][19] ), .B(n1629), .Z(\SUMB[44][18] ) );
  ND2P U2463 ( .A(\SUMB[43][19] ), .B(\ab[44][18] ), .Z(n1631) );
  ND3P U2464 ( .A(n1630), .B(n1631), .C(n1632), .Z(\CARRYB[44][18] ) );
  ND3 U2465 ( .A(n1661), .B(n1662), .C(n1663), .Z(\CARRYB[13][25] ) );
  EOP U2466 ( .A(\CARRYB[8][15] ), .B(n559), .Z(n1633) );
  ND2 U2467 ( .A(\SUMB[8][16] ), .B(\CARRYB[8][15] ), .Z(n1634) );
  ND2 U2468 ( .A(\SUMB[8][16] ), .B(n559), .Z(n1635) );
  ND3P U2469 ( .A(n1634), .B(n1635), .C(n1636), .Z(\CARRYB[9][15] ) );
  EO3 U2470 ( .A(\CARRYB[45][4] ), .B(n302), .C(n1474), .Z(\SUMB[46][4] ) );
  EO3 U2471 ( .A(\CARRYB[34][7] ), .B(n450), .C(\SUMB[34][8] ), .Z(
        \SUMB[35][7] ) );
  ND2 U2472 ( .A(\CARRYB[34][7] ), .B(\SUMB[34][8] ), .Z(n1640) );
  ND2 U2473 ( .A(\CARRYB[34][7] ), .B(n450), .Z(n1641) );
  ND2 U2474 ( .A(\SUMB[34][8] ), .B(n450), .Z(n1642) );
  ND3P U2475 ( .A(n1640), .B(n1641), .C(n1642), .Z(\CARRYB[35][7] ) );
  EO3 U2476 ( .A(\SUMB[5][16] ), .B(n449), .C(\CARRYB[5][15] ), .Z(
        \SUMB[6][15] ) );
  ND2 U2477 ( .A(\CARRYB[45][0] ), .B(n887), .Z(n2132) );
  EO3 U2478 ( .A(\CARRYB[28][22] ), .B(\ab[29][22] ), .C(\SUMB[28][23] ), .Z(
        \SUMB[29][22] ) );
  ND2 U2479 ( .A(\SUMB[28][23] ), .B(\ab[29][22] ), .Z(n1648) );
  ND3P U2480 ( .A(n1646), .B(n1647), .C(n1648), .Z(\CARRYB[29][22] ) );
  EOP U2481 ( .A(\SUMB[13][16] ), .B(n1681), .Z(\SUMB[14][15] ) );
  EOP U2482 ( .A(\CARRYB[16][10] ), .B(n600), .Z(n1649) );
  EOP U2483 ( .A(\SUMB[16][11] ), .B(n1649), .Z(\SUMB[17][10] ) );
  ND2 U2484 ( .A(\SUMB[16][11] ), .B(\CARRYB[16][10] ), .Z(n1650) );
  ND2 U2485 ( .A(\SUMB[16][11] ), .B(n600), .Z(n1651) );
  ND2 U2486 ( .A(\CARRYB[16][10] ), .B(n600), .Z(n1652) );
  ND3P U2487 ( .A(n1650), .B(n1651), .C(n1652), .Z(\CARRYB[17][10] ) );
  EOP U2488 ( .A(\CARRYB[6][28] ), .B(n471), .Z(n1653) );
  EOP U2489 ( .A(\SUMB[6][29] ), .B(n1653), .Z(\SUMB[7][28] ) );
  ND2 U2490 ( .A(\CARRYB[6][28] ), .B(n471), .Z(n1656) );
  ND2 U2491 ( .A(\CARRYB[26][20] ), .B(\SUMB[26][21] ), .Z(n1657) );
  ND2 U2492 ( .A(\SUMB[26][21] ), .B(\ab[27][20] ), .Z(n1659) );
  EOP U2493 ( .A(\CARRYB[12][25] ), .B(n683), .Z(n1660) );
  ND2 U2494 ( .A(\SUMB[12][26] ), .B(\CARRYB[12][25] ), .Z(n1661) );
  ND2 U2495 ( .A(\SUMB[12][26] ), .B(n683), .Z(n1662) );
  ND2 U2496 ( .A(\CARRYB[12][25] ), .B(n683), .Z(n1663) );
  ND2P U2497 ( .A(n321), .B(n1693), .Z(n1676) );
  ND2 U2498 ( .A(n2201), .B(\SUMB[44][2] ), .Z(n2147) );
  AN2 U2499 ( .A(n347), .B(A[1]), .Z(n2423) );
  ND2P U2500 ( .A(n322), .B(n1664), .Z(n1675) );
  EO3 U2501 ( .A(\CARRYB[12][10] ), .B(n596), .C(\SUMB[12][11] ), .Z(
        \SUMB[13][10] ) );
  ND2 U2502 ( .A(\CARRYB[12][10] ), .B(\SUMB[12][11] ), .Z(n1665) );
  ND2 U2503 ( .A(\CARRYB[12][10] ), .B(n596), .Z(n1666) );
  ND2 U2504 ( .A(\SUMB[12][11] ), .B(n596), .Z(n1667) );
  ND3 U2505 ( .A(n1665), .B(n1666), .C(n1667), .Z(\CARRYB[13][10] ) );
  ND3 U2506 ( .A(n2090), .B(n2091), .C(n2092), .Z(\CARRYB[9][14] ) );
  ND2 U2507 ( .A(\SUMB[40][25] ), .B(\CARRYB[40][24] ), .Z(n1668) );
  ND2 U2508 ( .A(\SUMB[40][25] ), .B(\ab[41][24] ), .Z(n1669) );
  ND2 U2509 ( .A(\CARRYB[40][24] ), .B(\ab[41][24] ), .Z(n1670) );
  ND3 U2510 ( .A(n1668), .B(n1669), .C(n1670), .Z(\CARRYB[41][24] ) );
  EOP U2511 ( .A(\CARRYB[19][32] ), .B(\ab[32][20] ), .Z(n1671) );
  EOP U2512 ( .A(\SUMB[19][33] ), .B(n1671), .Z(\SUMB[20][32] ) );
  ND2 U2513 ( .A(\SUMB[19][33] ), .B(\CARRYB[19][32] ), .Z(n1672) );
  ND2 U2514 ( .A(\SUMB[19][33] ), .B(\ab[32][20] ), .Z(n1673) );
  ND2 U2515 ( .A(\CARRYB[19][32] ), .B(\ab[32][20] ), .Z(n1674) );
  AN2 U2516 ( .A(n2180), .B(n2183), .Z(\CARRYB[1][11] ) );
  ND2P U2517 ( .A(n1675), .B(n1676), .Z(\SUMB[14][13] ) );
  EOP U2518 ( .A(\CARRYB[20][11] ), .B(n619), .Z(n1677) );
  EOP U2519 ( .A(\SUMB[20][12] ), .B(n1677), .Z(\SUMB[21][11] ) );
  ND2 U2520 ( .A(\CARRYB[20][11] ), .B(n619), .Z(n1680) );
  EO U2521 ( .A(\CARRYB[13][15] ), .B(n707), .Z(n1681) );
  AN2 U2522 ( .A(n2241), .B(n333), .Z(\CARRYB[1][14] ) );
  ND2 U2523 ( .A(\SUMB[28][31] ), .B(\CARRYB[28][30] ), .Z(n1683) );
  ND2 U2524 ( .A(\SUMB[28][31] ), .B(\ab[30][29] ), .Z(n1684) );
  ND2 U2525 ( .A(\CARRYB[28][30] ), .B(\ab[30][29] ), .Z(n1685) );
  EO3 U2526 ( .A(\CARRYB[26][23] ), .B(\ab[27][23] ), .C(\SUMB[26][24] ), .Z(
        \SUMB[27][23] ) );
  ND2P U2527 ( .A(\CARRYB[26][23] ), .B(\ab[27][23] ), .Z(n1687) );
  ND2 U2528 ( .A(\SUMB[26][24] ), .B(\ab[27][23] ), .Z(n1688) );
  ND3P U2529 ( .A(n1686), .B(n1687), .C(n1688), .Z(\CARRYB[27][23] ) );
  AN2 U2530 ( .A(\ab[13][13] ), .B(n2117), .Z(n2191) );
  ND2 U2531 ( .A(\SUMB[21][18] ), .B(\CARRYB[21][17] ), .Z(n1690) );
  ND2 U2532 ( .A(\SUMB[21][18] ), .B(\ab[22][17] ), .Z(n1691) );
  ND2 U2533 ( .A(\CARRYB[21][17] ), .B(\ab[22][17] ), .Z(n1692) );
  ND3P U2534 ( .A(n1690), .B(n1691), .C(n1692), .Z(\CARRYB[22][17] ) );
  ND2 U2535 ( .A(\CARRYB[13][13] ), .B(\SUMB[13][14] ), .Z(n1694) );
  ND2 U2536 ( .A(\CARRYB[13][13] ), .B(n675), .Z(n1695) );
  ND2 U2537 ( .A(\SUMB[13][14] ), .B(n675), .Z(n1696) );
  AN2 U2538 ( .A(n2164), .B(n2169), .Z(\CARRYB[1][29] ) );
  ND2P U2539 ( .A(\CARRYB[9][13] ), .B(\SUMB[9][14] ), .Z(n1994) );
  ND2P U2540 ( .A(n596), .B(\SUMB[9][14] ), .Z(n1993) );
  EOP U2541 ( .A(\SUMB[9][14] ), .B(n1831), .Z(\SUMB[10][13] ) );
  ND2 U2542 ( .A(\SUMB[24][30] ), .B(\CARRYB[24][29] ), .Z(n1697) );
  ND2 U2543 ( .A(\SUMB[24][30] ), .B(\ab[29][25] ), .Z(n1698) );
  ND2 U2544 ( .A(\CARRYB[24][29] ), .B(\ab[29][25] ), .Z(n1699) );
  EO3 U2545 ( .A(\CARRYB[26][28] ), .B(\ab[28][27] ), .C(\SUMB[26][29] ), .Z(
        \SUMB[27][28] ) );
  ND2P U2546 ( .A(\CARRYB[26][28] ), .B(\SUMB[26][29] ), .Z(n1700) );
  ND2P U2547 ( .A(\CARRYB[26][28] ), .B(\ab[28][27] ), .Z(n1701) );
  EOP U2548 ( .A(\CARRYB[44][3] ), .B(n2290), .Z(n1703) );
  ND2 U2549 ( .A(\SUMB[44][4] ), .B(\CARRYB[44][3] ), .Z(n1704) );
  ND2 U2550 ( .A(\SUMB[44][4] ), .B(n2290), .Z(n1705) );
  ND2 U2551 ( .A(\CARRYB[44][3] ), .B(n2290), .Z(n1706) );
  ND2 U2552 ( .A(\SUMB[23][11] ), .B(\CARRYB[23][10] ), .Z(n1708) );
  ND2 U2553 ( .A(\SUMB[23][11] ), .B(n597), .Z(n1709) );
  ND2 U2554 ( .A(\CARRYB[23][10] ), .B(n597), .Z(n1710) );
  EOP U2555 ( .A(\CARRYB[18][12] ), .B(n658), .Z(n1711) );
  EOP U2556 ( .A(\SUMB[18][13] ), .B(n1711), .Z(\SUMB[19][12] ) );
  ND2 U2557 ( .A(\SUMB[18][13] ), .B(\CARRYB[18][12] ), .Z(n1712) );
  ND2 U2558 ( .A(\SUMB[18][13] ), .B(n658), .Z(n1713) );
  ND2 U2559 ( .A(\CARRYB[18][12] ), .B(n658), .Z(n1714) );
  ND3 U2560 ( .A(n1712), .B(n1713), .C(n1714), .Z(\CARRYB[19][12] ) );
  EOP U2561 ( .A(n2203), .B(n2201), .Z(\SUMB[1][45] ) );
  ND2 U2562 ( .A(\SUMB[26][22] ), .B(\CARRYB[26][21] ), .Z(n1715) );
  ND2 U2563 ( .A(\SUMB[26][22] ), .B(\ab[27][21] ), .Z(n1716) );
  ND2 U2564 ( .A(\CARRYB[26][21] ), .B(\ab[27][21] ), .Z(n1717) );
  ND3 U2565 ( .A(n1715), .B(n1716), .C(n1717), .Z(\CARRYB[27][21] ) );
  ND3 U2566 ( .A(n1775), .B(n1776), .C(n1777), .Z(\CARRYB[5][16] ) );
  EO3P U2567 ( .A(\CARRYB[6][32] ), .B(n476), .C(\SUMB[6][33] ), .Z(
        \SUMB[7][32] ) );
  ND2 U2568 ( .A(\CARRYB[6][32] ), .B(\SUMB[6][33] ), .Z(n1718) );
  ND2 U2569 ( .A(\CARRYB[6][32] ), .B(n476), .Z(n1719) );
  ND2 U2570 ( .A(\SUMB[6][33] ), .B(n476), .Z(n1720) );
  ND3 U2571 ( .A(n1718), .B(n1719), .C(n1720), .Z(\CARRYB[7][32] ) );
  ND2 U2572 ( .A(\CARRYB[15][29] ), .B(\SUMB[15][30] ), .Z(n1871) );
  ND2 U2573 ( .A(\SUMB[15][30] ), .B(\ab[29][16] ), .Z(n1873) );
  EO3P U2574 ( .A(\CARRYB[18][16] ), .B(\ab[19][16] ), .C(\SUMB[18][17] ), .Z(
        \SUMB[19][16] ) );
  ND2 U2575 ( .A(\CARRYB[18][16] ), .B(\SUMB[18][17] ), .Z(n1721) );
  ND2 U2576 ( .A(\CARRYB[18][16] ), .B(\ab[19][16] ), .Z(n1722) );
  ND2 U2577 ( .A(\SUMB[18][17] ), .B(\ab[19][16] ), .Z(n1723) );
  ND3 U2578 ( .A(n1721), .B(n1722), .C(n1723), .Z(\CARRYB[19][16] ) );
  EOP U2579 ( .A(n1724), .B(\SUMB[42][10] ), .Z(\SUMB[43][9] ) );
  ND2P U2580 ( .A(\SUMB[42][10] ), .B(\CARRYB[42][9] ), .Z(n1725) );
  ND2P U2581 ( .A(\SUMB[42][10] ), .B(n586), .Z(n1726) );
  ND2 U2582 ( .A(\CARRYB[42][9] ), .B(n586), .Z(n1727) );
  ND3P U2583 ( .A(n1725), .B(n1726), .C(n1727), .Z(\CARRYB[43][9] ) );
  EO3 U2584 ( .A(\CARRYB[7][17] ), .B(n517), .C(\SUMB[7][18] ), .Z(
        \SUMB[8][17] ) );
  ND2 U2585 ( .A(\CARRYB[7][17] ), .B(\SUMB[7][18] ), .Z(n1728) );
  ND2 U2586 ( .A(\CARRYB[7][17] ), .B(n517), .Z(n1729) );
  ND2 U2587 ( .A(\SUMB[7][18] ), .B(n517), .Z(n1730) );
  ND3 U2588 ( .A(n1728), .B(n1729), .C(n1730), .Z(\CARRYB[8][17] ) );
  EOP U2589 ( .A(\CARRYB[25][8] ), .B(n523), .Z(n1732) );
  ND2 U2590 ( .A(\SUMB[25][9] ), .B(\CARRYB[25][8] ), .Z(n1733) );
  ND2 U2591 ( .A(\SUMB[25][9] ), .B(n523), .Z(n1734) );
  ND2 U2592 ( .A(\CARRYB[25][8] ), .B(n523), .Z(n1735) );
  EO U2593 ( .A(\ab[44][15] ), .B(\SUMB[43][16] ), .Z(n1908) );
  ND2 U2594 ( .A(n715), .B(\CARRYB[25][15] ), .Z(n1786) );
  EOP U2595 ( .A(\CARRYB[39][15] ), .B(\ab[40][15] ), .Z(n1736) );
  ND2 U2596 ( .A(\SUMB[39][16] ), .B(\CARRYB[39][15] ), .Z(n1737) );
  ND2 U2597 ( .A(\SUMB[39][16] ), .B(\ab[40][15] ), .Z(n1738) );
  ND2 U2598 ( .A(\CARRYB[39][15] ), .B(\ab[40][15] ), .Z(n1739) );
  ND2 U2599 ( .A(\CARRYB[2][22] ), .B(\SUMB[2][23] ), .Z(n1742) );
  ND2 U2600 ( .A(\CARRYB[2][22] ), .B(n2292), .Z(n1743) );
  ND2 U2601 ( .A(\SUMB[2][23] ), .B(n2292), .Z(n1744) );
  ND3 U2602 ( .A(n1742), .B(n1743), .C(n1744), .Z(n1745) );
  IVAP U2603 ( .A(n2053), .Z(n2054) );
  IVP U2604 ( .A(\SUMB[8][15] ), .Z(n2053) );
  EO3P U2605 ( .A(\CARRYB[11][14] ), .B(n659), .C(\SUMB[11][15] ), .Z(
        \SUMB[12][14] ) );
  ND2 U2606 ( .A(\CARRYB[11][14] ), .B(\SUMB[11][15] ), .Z(n1746) );
  ND2 U2607 ( .A(\CARRYB[11][14] ), .B(n659), .Z(n1747) );
  ND2 U2608 ( .A(\SUMB[11][15] ), .B(n659), .Z(n1748) );
  EOP U2609 ( .A(\CARRYB[1][22] ), .B(n2263), .Z(n1749) );
  ND2 U2610 ( .A(\SUMB[1][23] ), .B(\CARRYB[1][22] ), .Z(n1750) );
  ND2 U2611 ( .A(\SUMB[1][23] ), .B(n2263), .Z(n1751) );
  ND2 U2612 ( .A(\CARRYB[1][22] ), .B(n2263), .Z(n1752) );
  ND3P U2613 ( .A(n1750), .B(n1751), .C(n1752), .Z(\CARRYB[2][22] ) );
  EOP U2614 ( .A(\SUMB[5][21] ), .B(n1753), .Z(\SUMB[6][20] ) );
  ND2P U2615 ( .A(\SUMB[5][21] ), .B(\CARRYB[5][20] ), .Z(n1754) );
  ND2P U2616 ( .A(\SUMB[5][21] ), .B(n429), .Z(n1755) );
  ND2 U2617 ( .A(\CARRYB[5][20] ), .B(n429), .Z(n1756) );
  ND3P U2618 ( .A(n1754), .B(n1755), .C(n1756), .Z(\CARRYB[6][20] ) );
  ND2P U2619 ( .A(\CARRYB[6][20] ), .B(n470), .Z(n1769) );
  EOP U2620 ( .A(\CARRYB[10][21] ), .B(n619), .Z(n1757) );
  EOP U2621 ( .A(\SUMB[10][22] ), .B(n1757), .Z(\SUMB[11][21] ) );
  ND2 U2622 ( .A(\SUMB[10][22] ), .B(\CARRYB[10][21] ), .Z(n1758) );
  ND2 U2623 ( .A(\SUMB[10][22] ), .B(n619), .Z(n1759) );
  ND2 U2624 ( .A(\CARRYB[10][21] ), .B(n619), .Z(n1760) );
  ND3 U2625 ( .A(n1758), .B(n1759), .C(n1760), .Z(\CARRYB[11][21] ) );
  EOP U2626 ( .A(n1761), .B(\SUMB[30][14] ), .Z(\SUMB[31][13] ) );
  EOP U2627 ( .A(\CARRYB[24][16] ), .B(\ab[25][16] ), .Z(n1762) );
  EOP U2628 ( .A(\SUMB[24][17] ), .B(n1762), .Z(\SUMB[25][16] ) );
  IVDA U2629 ( .A(\CARRYB[42][15] ), .Z(n1763) );
  B4IP U2630 ( .A(n2324), .Z(n2322) );
  ND2 U2631 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Z(n1765) );
  ND2 U2632 ( .A(\SUMB[7][21] ), .B(n515), .Z(n1766) );
  ND2 U2633 ( .A(\CARRYB[7][20] ), .B(n515), .Z(n1767) );
  ND3P U2634 ( .A(n1765), .B(n1766), .C(n1767), .Z(\CARRYB[8][20] ) );
  EOP U2635 ( .A(n1839), .B(\SUMB[42][16] ), .Z(\SUMB[43][15] ) );
  EOP U2636 ( .A(\CARRYB[42][15] ), .B(\ab[43][15] ), .Z(n1839) );
  AN2P U2637 ( .A(A[7]), .B(A[0]), .Z(n2255) );
  AN2 U2638 ( .A(n2319), .B(n243), .Z(n2428) );
  EO3P U2639 ( .A(\CARRYB[6][20] ), .B(n470), .C(\SUMB[6][21] ), .Z(
        \SUMB[7][20] ) );
  ND2 U2640 ( .A(\CARRYB[6][20] ), .B(\SUMB[6][21] ), .Z(n1768) );
  ND2 U2641 ( .A(\SUMB[6][21] ), .B(n470), .Z(n1770) );
  ND3P U2642 ( .A(n1768), .B(n1769), .C(n1770), .Z(\CARRYB[7][20] ) );
  EO3 U2643 ( .A(\CARRYB[3][16] ), .B(n359), .C(\SUMB[3][17] ), .Z(
        \SUMB[4][16] ) );
  ND2 U2644 ( .A(\SUMB[3][17] ), .B(n359), .Z(n1773) );
  ND3P U2645 ( .A(n1771), .B(n1772), .C(n1773), .Z(\CARRYB[4][16] ) );
  ND2 U2646 ( .A(\SUMB[4][17] ), .B(\CARRYB[4][16] ), .Z(n1775) );
  ND2 U2647 ( .A(\SUMB[4][17] ), .B(n400), .Z(n1776) );
  ND2 U2648 ( .A(\CARRYB[4][16] ), .B(n400), .Z(n1777) );
  EOP U2649 ( .A(\SUMB[9][21] ), .B(n1778), .Z(\SUMB[10][20] ) );
  ND2 U2650 ( .A(\SUMB[9][21] ), .B(n1741), .Z(n1779) );
  ND2 U2651 ( .A(\SUMB[9][21] ), .B(n581), .Z(n1780) );
  ND2 U2652 ( .A(n1741), .B(n581), .Z(n1781) );
  ND3 U2653 ( .A(n1779), .B(n1780), .C(n1781), .Z(\CARRYB[10][20] ) );
  EOP U2654 ( .A(n715), .B(\CARRYB[25][15] ), .Z(n1782) );
  ND2 U2655 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .Z(n1783) );
  ND2 U2656 ( .A(\ab[25][16] ), .B(\SUMB[24][17] ), .Z(n1784) );
  ND2 U2657 ( .A(\CARRYB[24][16] ), .B(\SUMB[24][17] ), .Z(n1785) );
  ND2 U2658 ( .A(\CARRYB[30][13] ), .B(\SUMB[30][14] ), .Z(n1789) );
  ND2 U2659 ( .A(\CARRYB[30][13] ), .B(n685), .Z(n1790) );
  ND2 U2660 ( .A(\SUMB[30][14] ), .B(n685), .Z(n1791) );
  ND3 U2661 ( .A(n1789), .B(n1790), .C(n1791), .Z(\CARRYB[31][13] ) );
  EOP U2662 ( .A(\SUMB[3][16] ), .B(n1792), .Z(\SUMB[4][15] ) );
  ND2 U2663 ( .A(\SUMB[3][16] ), .B(\CARRYB[3][15] ), .Z(n1793) );
  ND2 U2664 ( .A(\SUMB[3][16] ), .B(n367), .Z(n1794) );
  ND2 U2665 ( .A(\CARRYB[3][15] ), .B(n367), .Z(n1795) );
  AN2 U2666 ( .A(n347), .B(n2117), .Z(n2424) );
  ND2 U2667 ( .A(\SUMB[45][25] ), .B(\ab[46][24] ), .Z(n1961) );
  ND3 U2668 ( .A(n1960), .B(n1961), .C(n1962), .Z(\CARRYB[46][24] ) );
  EOP U2669 ( .A(\CARRYB[39][10] ), .B(n637), .Z(n1796) );
  EOP U2670 ( .A(\SUMB[39][11] ), .B(n1796), .Z(\SUMB[40][10] ) );
  ND2 U2671 ( .A(\CARRYB[39][10] ), .B(n637), .Z(n1799) );
  ND2 U2672 ( .A(\CARRYB[15][14] ), .B(\SUMB[15][15] ), .Z(n1800) );
  ND2 U2673 ( .A(\CARRYB[15][14] ), .B(n701), .Z(n1801) );
  ND2 U2674 ( .A(\SUMB[15][15] ), .B(n701), .Z(n1802) );
  ND3 U2675 ( .A(n1800), .B(n1801), .C(n1802), .Z(\CARRYB[16][14] ) );
  ND2 U2676 ( .A(\SUMB[3][37] ), .B(n2300), .Z(n1880) );
  ND2 U2677 ( .A(\SUMB[3][37] ), .B(n1071), .Z(n1879) );
  EOP U2678 ( .A(\SUMB[5][19] ), .B(n464), .Z(n1803) );
  ND2 U2679 ( .A(\CARRYB[5][18] ), .B(\SUMB[5][19] ), .Z(n1804) );
  ND2 U2680 ( .A(\CARRYB[5][18] ), .B(n464), .Z(n1805) );
  ND2 U2681 ( .A(\SUMB[5][19] ), .B(n464), .Z(n1806) );
  ND2 U2682 ( .A(\CARRYB[2][18] ), .B(\SUMB[2][19] ), .Z(n1807) );
  ND2 U2683 ( .A(\CARRYB[2][18] ), .B(n2278), .Z(n1808) );
  ND2 U2684 ( .A(\SUMB[2][19] ), .B(n2278), .Z(n1809) );
  EOP U2685 ( .A(\CARRYB[4][21] ), .B(n395), .Z(n1810) );
  EOP U2686 ( .A(\SUMB[4][22] ), .B(n1810), .Z(\SUMB[5][21] ) );
  ND2P U2687 ( .A(\SUMB[4][22] ), .B(\CARRYB[4][21] ), .Z(n1811) );
  ND2P U2688 ( .A(\SUMB[4][22] ), .B(n395), .Z(n1812) );
  ND3P U2689 ( .A(n1811), .B(n1812), .C(n1813), .Z(\CARRYB[5][21] ) );
  EOP U2690 ( .A(\CARRYB[41][4] ), .B(n384), .Z(n1814) );
  ND2 U2691 ( .A(\CARRYB[41][4] ), .B(n384), .Z(n1817) );
  ND2 U2692 ( .A(\CARRYB[27][8] ), .B(\SUMB[27][9] ), .Z(n1818) );
  ND2 U2693 ( .A(\CARRYB[27][8] ), .B(n530), .Z(n1819) );
  ND2 U2694 ( .A(\SUMB[27][9] ), .B(n530), .Z(n1820) );
  ND3 U2695 ( .A(n1818), .B(n1819), .C(n1820), .Z(\CARRYB[28][8] ) );
  AN2P U2696 ( .A(n2166), .B(n2174), .Z(\CARRYB[1][27] ) );
  EO3P U2697 ( .A(\SUMB[17][29] ), .B(\ab[28][18] ), .C(\CARRYB[17][28] ), .Z(
        \SUMB[18][28] ) );
  B3IP U2698 ( .A(\ab[1][1] ), .Z1(n2039), .Z2(n2070) );
  B3I U2699 ( .A(n2324), .Z1(n2319) );
  ND2 U2700 ( .A(\CARRYB[20][15] ), .B(\SUMB[20][16] ), .Z(n1821) );
  ND2 U2701 ( .A(\CARRYB[20][15] ), .B(n719), .Z(n1822) );
  ND2 U2702 ( .A(\SUMB[20][16] ), .B(n719), .Z(n1823) );
  ND2 U2703 ( .A(\SUMB[13][16] ), .B(\CARRYB[13][15] ), .Z(n1824) );
  ND2 U2704 ( .A(\SUMB[13][16] ), .B(n707), .Z(n1825) );
  ND2 U2705 ( .A(\CARRYB[13][15] ), .B(n707), .Z(n1826) );
  ND2P U2706 ( .A(\SUMB[11][20] ), .B(n658), .Z(n1829) );
  ND2 U2707 ( .A(\CARRYB[11][19] ), .B(n658), .Z(n1830) );
  B4IP U2708 ( .A(n2324), .Z(n2321) );
  EOP U2709 ( .A(\SUMB[3][23] ), .B(n1958), .Z(\SUMB[4][22] ) );
  EOP U2710 ( .A(\CARRYB[3][22] ), .B(n356), .Z(n1958) );
  EOP U2711 ( .A(n2235), .B(n2240), .Z(\SUMB[1][24] ) );
  ND2 U2712 ( .A(\SUMB[45][25] ), .B(\CARRYB[45][24] ), .Z(n1960) );
  EO U2713 ( .A(\CARRYB[9][13] ), .B(n596), .Z(n1831) );
  EOP U2714 ( .A(n2089), .B(\CARRYB[8][14] ), .Z(\SUMB[9][14] ) );
  ND2P U2715 ( .A(\CARRYB[27][37] ), .B(\SUMB[27][38] ), .Z(n1833) );
  ND2 U2716 ( .A(\SUMB[27][38] ), .B(\ab[37][28] ), .Z(n1835) );
  EO3P U2717 ( .A(\CARRYB[20][29] ), .B(\ab[29][21] ), .C(\SUMB[20][30] ), .Z(
        \SUMB[21][29] ) );
  ND2 U2718 ( .A(\CARRYB[20][29] ), .B(\SUMB[20][30] ), .Z(n1836) );
  ND2 U2719 ( .A(\CARRYB[20][29] ), .B(\ab[29][21] ), .Z(n1837) );
  ND2 U2720 ( .A(\SUMB[20][30] ), .B(\ab[29][21] ), .Z(n1838) );
  ND3P U2721 ( .A(n1836), .B(n1837), .C(n1838), .Z(\CARRYB[21][29] ) );
  EO3P U2722 ( .A(\CARRYB[28][38] ), .B(\ab[38][29] ), .C(\SUMB[28][39] ), .Z(
        \SUMB[29][38] ) );
  ND2 U2723 ( .A(\CARRYB[28][38] ), .B(\SUMB[28][39] ), .Z(n1840) );
  ND2 U2724 ( .A(\CARRYB[28][38] ), .B(\ab[38][29] ), .Z(n1841) );
  ND2 U2725 ( .A(\SUMB[28][39] ), .B(\ab[38][29] ), .Z(n1842) );
  ND2 U2726 ( .A(\CARRYB[14][43] ), .B(\SUMB[14][44] ), .Z(n1844) );
  ND2 U2727 ( .A(\SUMB[14][44] ), .B(\ab[43][15] ), .Z(n1846) );
  ND2P U2728 ( .A(\CARRYB[36][33] ), .B(\ab[37][33] ), .Z(n1848) );
  ND2 U2729 ( .A(\SUMB[36][34] ), .B(\ab[37][33] ), .Z(n1849) );
  ND2 U2730 ( .A(\CARRYB[45][21] ), .B(\SUMB[45][22] ), .Z(n1850) );
  ND2 U2731 ( .A(\CARRYB[45][21] ), .B(\ab[46][21] ), .Z(n1851) );
  ND2 U2732 ( .A(\SUMB[45][22] ), .B(\ab[46][21] ), .Z(n1852) );
  ND2P U2733 ( .A(\CARRYB[40][36] ), .B(\ab[41][36] ), .Z(n1855) );
  ND2 U2734 ( .A(\SUMB[40][37] ), .B(\ab[41][36] ), .Z(n1856) );
  EOP U2735 ( .A(\SUMB[38][5] ), .B(n383), .Z(n1857) );
  EOP U2736 ( .A(\CARRYB[38][4] ), .B(n1857), .Z(\SUMB[39][4] ) );
  ND2 U2737 ( .A(\CARRYB[38][4] ), .B(\SUMB[38][5] ), .Z(n1858) );
  ND2 U2738 ( .A(\CARRYB[38][4] ), .B(n383), .Z(n1859) );
  ND2 U2739 ( .A(\SUMB[38][5] ), .B(n383), .Z(n1860) );
  EO3P U2740 ( .A(n1063), .B(\CARRYB[34][0] ), .C(\SUMB[34][1] ), .Z(\A1[33] )
         );
  ND2 U2741 ( .A(n1063), .B(\SUMB[34][1] ), .Z(n1862) );
  EO U2742 ( .A(n2172), .B(\SUMB[35][1] ), .Z(n1864) );
  EO U2743 ( .A(n1864), .B(\CARRYB[35][0] ), .Z(\A1[34] ) );
  ND2 U2744 ( .A(n2172), .B(\SUMB[35][1] ), .Z(n1865) );
  ND2 U2745 ( .A(n2172), .B(\CARRYB[35][0] ), .Z(n1866) );
  ND2 U2746 ( .A(\SUMB[35][1] ), .B(\CARRYB[35][0] ), .Z(n1867) );
  ND2 U2747 ( .A(\CARRYB[15][37] ), .B(\SUMB[15][38] ), .Z(n1868) );
  ND2 U2748 ( .A(\CARRYB[15][37] ), .B(\ab[37][16] ), .Z(n1869) );
  ND2 U2749 ( .A(\SUMB[15][38] ), .B(\ab[37][16] ), .Z(n1870) );
  ND3P U2750 ( .A(n1868), .B(n1869), .C(n1870), .Z(\CARRYB[16][37] ) );
  ND2 U2751 ( .A(\CARRYB[15][29] ), .B(\ab[29][16] ), .Z(n1872) );
  ND3P U2752 ( .A(n1871), .B(n1872), .C(n1873), .Z(\CARRYB[16][29] ) );
  EOP U2753 ( .A(\SUMB[22][9] ), .B(n1874), .Z(\SUMB[23][8] ) );
  ND2 U2754 ( .A(\CARRYB[22][8] ), .B(n533), .Z(n1877) );
  EOP U2755 ( .A(\CARRYB[3][36] ), .B(n2300), .Z(n1878) );
  EOP U2756 ( .A(\SUMB[3][37] ), .B(n1878), .Z(\SUMB[4][36] ) );
  ND2 U2757 ( .A(n1071), .B(n2300), .Z(n1881) );
  ND3P U2758 ( .A(n1879), .B(n1880), .C(n1881), .Z(\CARRYB[4][36] ) );
  EO3P U2759 ( .A(\SUMB[46][26] ), .B(\ab[47][25] ), .C(\CARRYB[46][25] ), .Z(
        \SUMB[47][25] ) );
  ND2 U2760 ( .A(\CARRYB[46][25] ), .B(\SUMB[46][26] ), .Z(n1882) );
  ND2 U2761 ( .A(\CARRYB[46][25] ), .B(\ab[47][25] ), .Z(n1883) );
  ND2 U2762 ( .A(\SUMB[46][26] ), .B(\ab[47][25] ), .Z(n1884) );
  ND2 U2763 ( .A(\CARRYB[36][29] ), .B(\SUMB[36][30] ), .Z(n1885) );
  ND2 U2764 ( .A(\CARRYB[36][29] ), .B(\ab[37][29] ), .Z(n1886) );
  ND2 U2765 ( .A(\SUMB[36][30] ), .B(\ab[37][29] ), .Z(n1887) );
  ND3P U2766 ( .A(n1885), .B(n1886), .C(n1887), .Z(\CARRYB[37][29] ) );
  EO3 U2767 ( .A(\CARRYB[17][36] ), .B(\ab[36][18] ), .C(\SUMB[17][37] ), .Z(
        \SUMB[18][36] ) );
  ND2 U2768 ( .A(\CARRYB[17][36] ), .B(\SUMB[17][37] ), .Z(n1888) );
  ND2 U2769 ( .A(\CARRYB[17][36] ), .B(\ab[36][18] ), .Z(n1889) );
  ND2 U2770 ( .A(\SUMB[17][37] ), .B(\ab[36][18] ), .Z(n1890) );
  ND2 U2771 ( .A(n2181), .B(\SUMB[32][2] ), .Z(n1892) );
  ND3P U2772 ( .A(n1891), .B(n1892), .C(n1893), .Z(\CARRYB[33][1] ) );
  EO U2773 ( .A(n2178), .B(\SUMB[33][2] ), .Z(n1894) );
  EOP U2774 ( .A(n1894), .B(\CARRYB[33][1] ), .Z(\SUMB[34][1] ) );
  ND2 U2775 ( .A(n2178), .B(\SUMB[33][2] ), .Z(n1895) );
  ND2 U2776 ( .A(n2178), .B(\CARRYB[33][1] ), .Z(n1896) );
  ND2 U2777 ( .A(\SUMB[33][2] ), .B(\CARRYB[33][1] ), .Z(n1897) );
  EOP U2778 ( .A(\CARRYB[32][8] ), .B(n537), .Z(n1898) );
  EOP U2779 ( .A(\SUMB[44][31] ), .B(\ab[45][30] ), .Z(n1899) );
  EOP U2780 ( .A(\CARRYB[44][30] ), .B(n1899), .Z(\SUMB[45][30] ) );
  ND2 U2781 ( .A(\CARRYB[44][30] ), .B(\SUMB[44][31] ), .Z(n1900) );
  ND2 U2782 ( .A(\CARRYB[44][30] ), .B(\ab[45][30] ), .Z(n1901) );
  ND2 U2783 ( .A(\SUMB[44][31] ), .B(\ab[45][30] ), .Z(n1902) );
  ND3P U2784 ( .A(n1900), .B(n1901), .C(n1902), .Z(\CARRYB[45][30] ) );
  EOP U2785 ( .A(\CARRYB[41][16] ), .B(\ab[42][16] ), .Z(n1903) );
  EOP U2786 ( .A(\SUMB[41][17] ), .B(n1903), .Z(\SUMB[42][16] ) );
  ND2 U2787 ( .A(\ab[43][15] ), .B(n1763), .Z(n1905) );
  ND2 U2788 ( .A(\ab[43][15] ), .B(\SUMB[42][16] ), .Z(n1906) );
  ND2 U2789 ( .A(n1763), .B(\SUMB[42][16] ), .Z(n1907) );
  ND2 U2790 ( .A(\ab[44][15] ), .B(\SUMB[43][16] ), .Z(n1909) );
  ND2 U2791 ( .A(\ab[44][15] ), .B(\CARRYB[43][15] ), .Z(n1910) );
  ND2 U2792 ( .A(\SUMB[43][16] ), .B(\CARRYB[43][15] ), .Z(n1911) );
  ND3 U2793 ( .A(n1909), .B(n1910), .C(n1911), .Z(\CARRYB[44][15] ) );
  ND2 U2794 ( .A(n584), .B(\CARRYB[22][9] ), .Z(n1913) );
  ND2 U2795 ( .A(n584), .B(\SUMB[22][10] ), .Z(n1914) );
  ND2 U2796 ( .A(\CARRYB[22][9] ), .B(\SUMB[22][10] ), .Z(n1915) );
  ND3 U2797 ( .A(n1913), .B(n1914), .C(n1915), .Z(\CARRYB[23][9] ) );
  ND2 U2798 ( .A(n534), .B(\CARRYB[23][8] ), .Z(n1916) );
  ND2P U2799 ( .A(n534), .B(\SUMB[23][9] ), .Z(n1917) );
  ND3P U2800 ( .A(n1916), .B(n1917), .C(n1918), .Z(\CARRYB[24][8] ) );
  EOP U2801 ( .A(\SUMB[18][8] ), .B(n497), .Z(n1919) );
  EOP U2802 ( .A(\CARRYB[18][7] ), .B(n1919), .Z(\SUMB[19][7] ) );
  ND2 U2803 ( .A(\CARRYB[18][7] ), .B(n497), .Z(n1921) );
  EOP U2804 ( .A(\SUMB[17][9] ), .B(n1926), .Z(\SUMB[18][8] ) );
  ND2 U2805 ( .A(\CARRYB[41][16] ), .B(\SUMB[41][17] ), .Z(n1923) );
  ND2 U2806 ( .A(\CARRYB[41][16] ), .B(\ab[42][16] ), .Z(n1924) );
  ND2 U2807 ( .A(\SUMB[41][17] ), .B(\ab[42][16] ), .Z(n1925) );
  ND2 U2808 ( .A(\CARRYB[17][28] ), .B(\SUMB[17][29] ), .Z(n1927) );
  ND2 U2809 ( .A(\CARRYB[17][28] ), .B(\ab[28][18] ), .Z(n1928) );
  ND2 U2810 ( .A(\SUMB[17][29] ), .B(\ab[28][18] ), .Z(n1929) );
  EO3P U2811 ( .A(n434), .B(\CARRYB[20][6] ), .C(\SUMB[20][7] ), .Z(
        \SUMB[21][6] ) );
  ND2 U2812 ( .A(n434), .B(\CARRYB[20][6] ), .Z(n1931) );
  ND2 U2813 ( .A(n434), .B(\SUMB[20][7] ), .Z(n1932) );
  ND2 U2814 ( .A(\CARRYB[20][6] ), .B(\SUMB[20][7] ), .Z(n1933) );
  ND2 U2815 ( .A(n380), .B(\CARRYB[21][5] ), .Z(n1934) );
  ND2P U2816 ( .A(\CARRYB[21][5] ), .B(\SUMB[21][6] ), .Z(n1936) );
  EOP U2817 ( .A(\SUMB[37][35] ), .B(\ab[38][34] ), .Z(n1937) );
  EOP U2818 ( .A(\CARRYB[37][34] ), .B(n1937), .Z(\SUMB[38][34] ) );
  ND2 U2819 ( .A(\CARRYB[37][34] ), .B(\SUMB[37][35] ), .Z(n1938) );
  ND2 U2820 ( .A(\CARRYB[37][34] ), .B(\ab[38][34] ), .Z(n1939) );
  ND2 U2821 ( .A(\SUMB[37][35] ), .B(\ab[38][34] ), .Z(n1940) );
  EO3 U2822 ( .A(n338), .B(\SUMB[1][8] ), .C(\CARRYB[1][7] ), .Z(\SUMB[2][7] )
         );
  ND2 U2823 ( .A(n338), .B(\CARRYB[1][7] ), .Z(n1941) );
  EOP U2824 ( .A(n2229), .B(n2232), .Z(\SUMB[1][8] ) );
  EOP U2825 ( .A(n1048), .B(\ab[46][16] ), .Z(n1944) );
  ND2 U2826 ( .A(\CARRYB[45][16] ), .B(\SUMB[45][17] ), .Z(n1945) );
  ND2 U2827 ( .A(\CARRYB[45][16] ), .B(\ab[46][16] ), .Z(n1946) );
  ND2 U2828 ( .A(\SUMB[45][17] ), .B(\ab[46][16] ), .Z(n1947) );
  ND3 U2829 ( .A(n1945), .B(n1946), .C(n1947), .Z(\CARRYB[46][16] ) );
  ND2 U2830 ( .A(\CARRYB[1][42] ), .B(\SUMB[1][43] ), .Z(n1948) );
  ND2 U2831 ( .A(\CARRYB[1][42] ), .B(n2265), .Z(n1949) );
  ND2 U2832 ( .A(\SUMB[1][43] ), .B(n2265), .Z(n1950) );
  ND3P U2833 ( .A(n1948), .B(n1949), .C(n1950), .Z(\CARRYB[2][42] ) );
  EOP U2834 ( .A(n2204), .B(n2202), .Z(\SUMB[1][43] ) );
  ND2P U2835 ( .A(\CARRYB[19][43] ), .B(\ab[43][20] ), .Z(n1953) );
  ND2 U2836 ( .A(\SUMB[19][44] ), .B(\ab[43][20] ), .Z(n1954) );
  EO3P U2837 ( .A(\CARRYB[19][10] ), .B(n581), .C(\SUMB[19][11] ), .Z(
        \SUMB[20][10] ) );
  ND2 U2838 ( .A(\CARRYB[19][10] ), .B(\SUMB[19][11] ), .Z(n1955) );
  ND2 U2839 ( .A(\SUMB[19][11] ), .B(n581), .Z(n1957) );
  ND3 U2840 ( .A(n1955), .B(n1956), .C(n1957), .Z(\CARRYB[20][10] ) );
  ND2 U2841 ( .A(\CARRYB[45][24] ), .B(\ab[46][24] ), .Z(n1962) );
  EO3P U2842 ( .A(\ab[42][14] ), .B(\CARRYB[13][42] ), .C(\SUMB[13][43] ), .Z(
        \SUMB[14][42] ) );
  EOP U2843 ( .A(n1963), .B(\SUMB[14][42] ), .Z(\SUMB[15][41] ) );
  ND2 U2844 ( .A(\ab[42][14] ), .B(\CARRYB[13][42] ), .Z(n1964) );
  ND2 U2845 ( .A(\ab[42][14] ), .B(\SUMB[13][43] ), .Z(n1965) );
  ND2 U2846 ( .A(\CARRYB[13][42] ), .B(\SUMB[13][43] ), .Z(n1966) );
  ND2 U2847 ( .A(\ab[41][15] ), .B(\CARRYB[14][41] ), .Z(n1967) );
  EOP U2848 ( .A(\SUMB[17][10] ), .B(n560), .Z(n1970) );
  EOP U2849 ( .A(\CARRYB[17][9] ), .B(n1970), .Z(\SUMB[18][9] ) );
  ND2 U2850 ( .A(\CARRYB[13][6] ), .B(\SUMB[13][7] ), .Z(n1972) );
  ND2 U2851 ( .A(\CARRYB[13][6] ), .B(n452), .Z(n1973) );
  ND2 U2852 ( .A(\SUMB[13][7] ), .B(n452), .Z(n1974) );
  EO3 U2853 ( .A(\CARRYB[1][13] ), .B(\SUMB[1][14] ), .C(n2266), .Z(
        \SUMB[2][13] ) );
  ND2 U2854 ( .A(\CARRYB[1][13] ), .B(n2266), .Z(n1975) );
  EO3 U2855 ( .A(\CARRYB[29][2] ), .B(n2208), .C(\SUMB[29][3] ), .Z(
        \SUMB[30][2] ) );
  ND2 U2856 ( .A(\CARRYB[29][2] ), .B(\SUMB[29][3] ), .Z(n1978) );
  ND2 U2857 ( .A(\CARRYB[29][2] ), .B(n2208), .Z(n1979) );
  ND2 U2858 ( .A(\SUMB[29][3] ), .B(n2208), .Z(n1980) );
  EO3 U2859 ( .A(\CARRYB[39][27] ), .B(\ab[40][27] ), .C(\SUMB[39][28] ), .Z(
        \SUMB[40][27] ) );
  ND2 U2860 ( .A(\CARRYB[39][27] ), .B(\SUMB[39][28] ), .Z(n1981) );
  ND2 U2861 ( .A(\CARRYB[39][27] ), .B(\ab[40][27] ), .Z(n1982) );
  ND2 U2862 ( .A(\SUMB[39][28] ), .B(\ab[40][27] ), .Z(n1983) );
  ND3P U2863 ( .A(n1981), .B(n1982), .C(n1983), .Z(\CARRYB[40][27] ) );
  ND2 U2864 ( .A(\CARRYB[45][32] ), .B(\SUMB[45][33] ), .Z(n1985) );
  ND2 U2865 ( .A(\CARRYB[45][32] ), .B(\ab[46][32] ), .Z(n1986) );
  ND2 U2866 ( .A(\SUMB[45][33] ), .B(\ab[46][32] ), .Z(n1987) );
  ND3P U2867 ( .A(n1985), .B(n1986), .C(n1987), .Z(\CARRYB[46][32] ) );
  EOP U2868 ( .A(\SUMB[22][26] ), .B(\ab[25][23] ), .Z(n1988) );
  EOP U2869 ( .A(n1988), .B(\CARRYB[22][25] ), .Z(\SUMB[23][25] ) );
  ND2 U2870 ( .A(\CARRYB[22][25] ), .B(\SUMB[22][26] ), .Z(n1989) );
  ND2 U2871 ( .A(\CARRYB[22][25] ), .B(\ab[25][23] ), .Z(n1990) );
  ND2 U2872 ( .A(\SUMB[22][26] ), .B(\ab[25][23] ), .Z(n1991) );
  ND2 U2873 ( .A(n596), .B(\CARRYB[9][13] ), .Z(n1992) );
  ND3P U2874 ( .A(n1992), .B(n1993), .C(n1994), .Z(\CARRYB[10][13] ) );
  EOP U2875 ( .A(n635), .B(\SUMB[10][14] ), .Z(n1995) );
  EOP U2876 ( .A(\CARRYB[10][13] ), .B(n1995), .Z(\SUMB[11][13] ) );
  ND2 U2877 ( .A(n635), .B(\SUMB[10][14] ), .Z(n1996) );
  ND2 U2878 ( .A(n635), .B(\CARRYB[10][13] ), .Z(n1997) );
  ND2 U2879 ( .A(\SUMB[10][14] ), .B(\CARRYB[10][13] ), .Z(n1998) );
  EO3P U2880 ( .A(\CARRYB[25][7] ), .B(n468), .C(\SUMB[25][8] ), .Z(
        \SUMB[26][7] ) );
  ND2 U2881 ( .A(\CARRYB[25][7] ), .B(\SUMB[25][8] ), .Z(n1999) );
  ND2 U2882 ( .A(\CARRYB[25][7] ), .B(n468), .Z(n2000) );
  ND2 U2883 ( .A(\SUMB[25][8] ), .B(n468), .Z(n2001) );
  ND2 U2884 ( .A(\CARRYB[17][9] ), .B(\SUMB[17][10] ), .Z(n2002) );
  ND2 U2885 ( .A(\CARRYB[17][9] ), .B(n560), .Z(n2003) );
  ND2 U2886 ( .A(\SUMB[17][10] ), .B(n560), .Z(n2004) );
  ND3P U2887 ( .A(n2002), .B(n2003), .C(n2004), .Z(\CARRYB[18][9] ) );
  ND2 U2888 ( .A(n1745), .B(\SUMB[3][23] ), .Z(n2005) );
  ND2 U2889 ( .A(n1745), .B(n356), .Z(n2006) );
  ND2 U2890 ( .A(\SUMB[3][23] ), .B(n356), .Z(n2007) );
  ND3P U2891 ( .A(n2005), .B(n2006), .C(n2007), .Z(\CARRYB[4][22] ) );
  ND2 U2892 ( .A(\CARRYB[37][1] ), .B(n2233), .Z(n2047) );
  EOP U2893 ( .A(\CARRYB[47][2] ), .B(\SUMB[47][3] ), .Z(\A1[48] ) );
  EO3P U2894 ( .A(n536), .B(\CARRYB[7][14] ), .C(\SUMB[7][15] ), .Z(
        \SUMB[8][14] ) );
  EOP U2895 ( .A(\CARRYB[47][22] ), .B(\SUMB[47][23] ), .Z(\A1[68] ) );
  AN2P U2896 ( .A(n2326), .B(n1350), .Z(n2429) );
  AN2P U2897 ( .A(n2319), .B(n1350), .Z(n2430) );
  AN2 U2898 ( .A(n2325), .B(PRODUCT[0]), .Z(n2425) );
  EOP U2899 ( .A(n2164), .B(n2169), .Z(\SUMB[1][29] ) );
  AN2 U2900 ( .A(n2323), .B(A[0]), .Z(n2427) );
  ND2 U2901 ( .A(\CARRYB[2][28] ), .B(\SUMB[2][29] ), .Z(n2008) );
  ND2 U2902 ( .A(\CARRYB[2][28] ), .B(n2284), .Z(n2009) );
  ND2 U2903 ( .A(\SUMB[2][29] ), .B(n2284), .Z(n2010) );
  ND2 U2904 ( .A(\CARRYB[9][27] ), .B(\SUMB[9][28] ), .Z(n2011) );
  ND2 U2905 ( .A(\CARRYB[9][27] ), .B(n611), .Z(n2012) );
  ND2 U2906 ( .A(\SUMB[9][28] ), .B(n611), .Z(n2013) );
  IVP U2907 ( .A(n377), .Z(n2336) );
  EO U2908 ( .A(\SUMB[35][3] ), .B(n2260), .Z(n2015) );
  EOP U2909 ( .A(\CARRYB[35][2] ), .B(n2015), .Z(\SUMB[36][2] ) );
  ND2P U2910 ( .A(\CARRYB[35][2] ), .B(n2260), .Z(n2017) );
  ND2 U2911 ( .A(\SUMB[35][3] ), .B(n2260), .Z(n2018) );
  ND3P U2912 ( .A(n2016), .B(n2017), .C(n2018), .Z(\CARRYB[36][2] ) );
  EOP U2913 ( .A(\SUMB[30][4] ), .B(n2268), .Z(n2019) );
  EOP U2914 ( .A(\CARRYB[30][3] ), .B(n2019), .Z(\SUMB[31][3] ) );
  ND2 U2915 ( .A(\SUMB[30][4] ), .B(n2268), .Z(n2022) );
  ND2P U2916 ( .A(\CARRYB[9][11] ), .B(n2024), .Z(n2025) );
  ND2 U2917 ( .A(n2023), .B(n2118), .Z(n2026) );
  ND2P U2918 ( .A(n2025), .B(n2026), .Z(\SUMB[10][11] ) );
  IVDA U2919 ( .A(\CARRYB[9][11] ), .Y(n2023) );
  IV U2920 ( .A(n2118), .Z(n2024) );
  EOP U2921 ( .A(\SUMB[9][12] ), .B(n606), .Z(n2118) );
  EOP U2922 ( .A(\SUMB[2][14] ), .B(n2287), .Z(n2027) );
  EOP U2923 ( .A(\CARRYB[2][13] ), .B(n2027), .Z(\SUMB[3][13] ) );
  ND2 U2924 ( .A(\CARRYB[2][13] ), .B(\SUMB[2][14] ), .Z(n2028) );
  ND2 U2925 ( .A(\CARRYB[2][13] ), .B(n2287), .Z(n2029) );
  ND2 U2926 ( .A(\SUMB[2][14] ), .B(n2287), .Z(n2030) );
  ND3 U2927 ( .A(n2028), .B(n2029), .C(n2030), .Z(\CARRYB[3][13] ) );
  ND2 U2928 ( .A(\SUMB[13][33] ), .B(\ab[32][14] ), .Z(n2034) );
  EOP U2929 ( .A(\SUMB[5][30] ), .B(n455), .Z(n2035) );
  EOP U2930 ( .A(\CARRYB[5][29] ), .B(n2035), .Z(\SUMB[6][29] ) );
  ND2 U2931 ( .A(\SUMB[5][30] ), .B(n455), .Z(n2038) );
  B4IP U2932 ( .A(n2039), .Z(n2040) );
  EOP U2933 ( .A(\SUMB[11][46] ), .B(\ab[45][12] ), .Z(n2041) );
  EOP U2934 ( .A(\CARRYB[11][45] ), .B(n2041), .Z(\SUMB[12][45] ) );
  ND2 U2935 ( .A(\SUMB[11][46] ), .B(\ab[45][12] ), .Z(n2044) );
  ND2 U2936 ( .A(\SUMB[37][2] ), .B(n2233), .Z(n2048) );
  ND2 U2937 ( .A(\CARRYB[24][1] ), .B(\SUMB[24][2] ), .Z(n2050) );
  ND2 U2938 ( .A(\CARRYB[24][1] ), .B(n2177), .Z(n2051) );
  ND2 U2939 ( .A(\SUMB[24][2] ), .B(n2177), .Z(n2052) );
  EO3P U2940 ( .A(\CARRYB[16][43] ), .B(\ab[43][17] ), .C(\SUMB[16][44] ), .Z(
        \SUMB[17][43] ) );
  ND2 U2941 ( .A(\CARRYB[16][43] ), .B(\SUMB[16][44] ), .Z(n2055) );
  ND2 U2942 ( .A(\CARRYB[16][43] ), .B(\ab[43][17] ), .Z(n2056) );
  ND2 U2943 ( .A(\SUMB[16][44] ), .B(\ab[43][17] ), .Z(n2057) );
  EOP U2944 ( .A(\SUMB[36][4] ), .B(n342), .Z(n2059) );
  EOP U2945 ( .A(\CARRYB[36][3] ), .B(n2059), .Z(\SUMB[37][3] ) );
  ND2P U2946 ( .A(\CARRYB[36][3] ), .B(\SUMB[36][4] ), .Z(n2060) );
  ND2P U2947 ( .A(\CARRYB[36][3] ), .B(n342), .Z(n2061) );
  ND2 U2948 ( .A(\SUMB[36][4] ), .B(n342), .Z(n2062) );
  EO3 U2949 ( .A(\CARRYB[2][30] ), .B(n2273), .C(\SUMB[2][31] ), .Z(
        \SUMB[3][30] ) );
  ND2 U2950 ( .A(n2273), .B(\CARRYB[2][30] ), .Z(n2063) );
  ND2 U2951 ( .A(n2273), .B(\SUMB[2][31] ), .Z(n2064) );
  ND2 U2952 ( .A(\CARRYB[2][30] ), .B(\SUMB[2][31] ), .Z(n2065) );
  EOP U2953 ( .A(n2281), .B(\SUMB[3][31] ), .Z(n2066) );
  EO U2954 ( .A(\SUMB[40][4] ), .B(n2286), .Z(n2078) );
  EO U2955 ( .A(\CARRYB[40][3] ), .B(n2078), .Z(\SUMB[41][3] ) );
  ND3 U2956 ( .A(n2079), .B(n2080), .C(n2081), .Z(\CARRYB[41][3] ) );
  ND3 U2957 ( .A(n2075), .B(n2076), .C(n2077), .Z(\CARRYB[3][7] ) );
  EO3 U2958 ( .A(\CARRYB[28][10] ), .B(n605), .C(\SUMB[28][11] ), .Z(
        \SUMB[29][10] ) );
  ND2 U2959 ( .A(\CARRYB[28][10] ), .B(\SUMB[28][11] ), .Z(n2071) );
  ND2 U2960 ( .A(\CARRYB[28][10] ), .B(n605), .Z(n2072) );
  ND2 U2961 ( .A(\SUMB[28][11] ), .B(n605), .Z(n2073) );
  ND3P U2962 ( .A(n2071), .B(n2072), .C(n2073), .Z(\CARRYB[29][10] ) );
  EOP U2963 ( .A(\SUMB[2][8] ), .B(n352), .Z(n2074) );
  EOP U2964 ( .A(\CARRYB[2][7] ), .B(n2074), .Z(\SUMB[3][7] ) );
  ND2 U2965 ( .A(\CARRYB[2][7] ), .B(\SUMB[2][8] ), .Z(n2075) );
  ND2 U2966 ( .A(\CARRYB[2][7] ), .B(n352), .Z(n2076) );
  ND2 U2967 ( .A(\SUMB[2][8] ), .B(n352), .Z(n2077) );
  ND2 U2968 ( .A(\CARRYB[40][3] ), .B(\SUMB[40][4] ), .Z(n2079) );
  ND2 U2969 ( .A(\CARRYB[40][3] ), .B(n2286), .Z(n2080) );
  ND2 U2970 ( .A(\SUMB[40][4] ), .B(n2286), .Z(n2081) );
  EOP U2971 ( .A(\SUMB[34][11] ), .B(n582), .Z(n2082) );
  EOP U2972 ( .A(\CARRYB[34][10] ), .B(n2082), .Z(\SUMB[35][10] ) );
  ND2 U2973 ( .A(\CARRYB[34][10] ), .B(\SUMB[34][11] ), .Z(n2083) );
  ND2 U2974 ( .A(\CARRYB[34][10] ), .B(n582), .Z(n2084) );
  ND2 U2975 ( .A(\SUMB[34][11] ), .B(n582), .Z(n2085) );
  ND3 U2976 ( .A(n2083), .B(n2084), .C(n2085), .Z(\CARRYB[35][10] ) );
  ND2 U2977 ( .A(n536), .B(\CARRYB[7][14] ), .Z(n2086) );
  ND2 U2978 ( .A(n536), .B(\SUMB[7][15] ), .Z(n2087) );
  ND2 U2979 ( .A(\CARRYB[7][14] ), .B(\SUMB[7][15] ), .Z(n2088) );
  ND2 U2980 ( .A(n576), .B(\SUMB[8][15] ), .Z(n2090) );
  ND2 U2981 ( .A(n576), .B(\CARRYB[8][14] ), .Z(n2091) );
  ND2 U2982 ( .A(\SUMB[8][15] ), .B(\CARRYB[8][14] ), .Z(n2092) );
  ND2 U2983 ( .A(\CARRYB[13][8] ), .B(\SUMB[13][9] ), .Z(n2094) );
  ND2 U2984 ( .A(\CARRYB[13][8] ), .B(n536), .Z(n2095) );
  ND3 U2985 ( .A(n2094), .B(n2095), .C(n2096), .Z(\CARRYB[14][8] ) );
  ND3 U2986 ( .A(n2097), .B(n2098), .C(n2099), .Z(\CARRYB[7][8] ) );
  ND2 U2987 ( .A(\SUMB[13][9] ), .B(n536), .Z(n2096) );
  EO3 U2988 ( .A(\CARRYB[6][8] ), .B(n518), .C(\SUMB[6][9] ), .Z(\SUMB[7][8] )
         );
  ND2 U2989 ( .A(\CARRYB[6][8] ), .B(\SUMB[6][9] ), .Z(n2097) );
  ND2 U2990 ( .A(\CARRYB[6][8] ), .B(n518), .Z(n2098) );
  ND2 U2991 ( .A(\SUMB[6][9] ), .B(n518), .Z(n2099) );
  EO3P U2992 ( .A(n2304), .B(\CARRYB[30][4] ), .C(\SUMB[30][5] ), .Z(
        \SUMB[31][4] ) );
  ND2 U2993 ( .A(n2304), .B(\SUMB[30][5] ), .Z(n2101) );
  ND2P U2994 ( .A(\CARRYB[30][4] ), .B(\SUMB[30][5] ), .Z(n2102) );
  ND3P U2995 ( .A(n2100), .B(n2101), .C(n2102), .Z(\CARRYB[31][4] ) );
  EOP U2996 ( .A(n358), .B(\SUMB[31][5] ), .Z(n2103) );
  EOP U2997 ( .A(n2103), .B(\CARRYB[31][4] ), .Z(\SUMB[32][4] ) );
  ND2 U2998 ( .A(n358), .B(\SUMB[31][5] ), .Z(n2104) );
  ND2 U2999 ( .A(\CARRYB[17][8] ), .B(\SUMB[17][9] ), .Z(n2107) );
  ND2 U3000 ( .A(\CARRYB[17][8] ), .B(n519), .Z(n2108) );
  ND2 U3001 ( .A(\SUMB[17][9] ), .B(n519), .Z(n2109) );
  EO U3002 ( .A(\SUMB[11][10] ), .B(n566), .Z(n2110) );
  EO U3003 ( .A(\CARRYB[11][9] ), .B(n2110), .Z(\SUMB[12][9] ) );
  ND2 U3004 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(n2111) );
  ND2 U3005 ( .A(\CARRYB[11][9] ), .B(n566), .Z(n2112) );
  ND2 U3006 ( .A(\SUMB[11][10] ), .B(n566), .Z(n2113) );
  ND2 U3007 ( .A(\CARRYB[32][8] ), .B(\SUMB[32][9] ), .Z(n2114) );
  ND2 U3008 ( .A(\CARRYB[32][8] ), .B(n537), .Z(n2115) );
  ND2 U3009 ( .A(\SUMB[32][9] ), .B(n537), .Z(n2116) );
  ND3P U3010 ( .A(n2114), .B(n2115), .C(n2116), .Z(\CARRYB[33][8] ) );
  ND3 U3011 ( .A(n2119), .B(n2120), .C(n2121), .Z(\CARRYB[10][11] ) );
  ND2 U3012 ( .A(\CARRYB[9][11] ), .B(\SUMB[9][12] ), .Z(n2119) );
  ND2 U3013 ( .A(\CARRYB[9][11] ), .B(n606), .Z(n2120) );
  ND2 U3014 ( .A(\SUMB[9][12] ), .B(n606), .Z(n2121) );
  ND2 U3015 ( .A(\CARRYB[34][5] ), .B(\SUMB[34][6] ), .Z(n2122) );
  ND2 U3016 ( .A(\CARRYB[34][5] ), .B(n374), .Z(n2123) );
  ND2 U3017 ( .A(\SUMB[34][6] ), .B(n374), .Z(n2124) );
  EO3 U3018 ( .A(\CARRYB[45][0] ), .B(n887), .C(n2125), .Z(\A1[44] ) );
  EO U3019 ( .A(n2146), .B(\CARRYB[44][1] ), .Z(n2125) );
  ND2 U3020 ( .A(\CARRYB[34][2] ), .B(\SUMB[34][3] ), .Z(n2128) );
  ND2 U3021 ( .A(\CARRYB[34][2] ), .B(n2214), .Z(n2129) );
  EOP U3022 ( .A(n2201), .B(\SUMB[44][2] ), .Z(n2146) );
  EOP U3023 ( .A(n2146), .B(\CARRYB[44][1] ), .Z(\SUMB[45][1] ) );
  EOP U3024 ( .A(\SUMB[34][3] ), .B(n2214), .Z(n2127) );
  EOP U3025 ( .A(\CARRYB[34][2] ), .B(n2127), .Z(\SUMB[35][2] ) );
  ND2 U3026 ( .A(\SUMB[34][3] ), .B(n2214), .Z(n2130) );
  EO U3027 ( .A(n2256), .B(n2253), .Z(\SUMB[1][4] ) );
  EO U3028 ( .A(\CARRYB[5][1] ), .B(n2139), .Z(\SUMB[6][1] ) );
  ND2 U3029 ( .A(\CARRYB[5][1] ), .B(\SUMB[5][2] ), .Z(n2140) );
  ND2 U3030 ( .A(\CARRYB[5][1] ), .B(n2242), .Z(n2141) );
  EO U3031 ( .A(\SUMB[9][2] ), .B(n2234), .Z(n2135) );
  ND2 U3032 ( .A(\SUMB[45][1] ), .B(n887), .Z(n2133) );
  ND2 U3033 ( .A(\CARRYB[9][1] ), .B(\SUMB[9][2] ), .Z(n2136) );
  ND2 U3034 ( .A(\CARRYB[9][1] ), .B(n2234), .Z(n2137) );
  ND2 U3035 ( .A(\SUMB[9][2] ), .B(n2234), .Z(n2138) );
  EO U3036 ( .A(\SUMB[5][2] ), .B(n2242), .Z(n2139) );
  ND2 U3037 ( .A(\SUMB[5][2] ), .B(n2242), .Z(n2142) );
  EOP U3038 ( .A(\CARRYB[47][31] ), .B(\SUMB[47][32] ), .Z(\A1[77] ) );
  EOP U3039 ( .A(n2193), .B(n2187), .Z(\SUMB[1][16] ) );
  EO U3040 ( .A(n289), .B(n2234), .Z(\SUMB[1][10] ) );
  EO U3041 ( .A(n2239), .B(n2195), .Z(\SUMB[1][40] ) );
  EO3 U3042 ( .A(n2237), .B(\CARRYB[43][1] ), .C(\SUMB[43][2] ), .Z(
        \SUMB[44][1] ) );
  ND2 U3043 ( .A(n2237), .B(\CARRYB[43][1] ), .Z(n2143) );
  ND2 U3044 ( .A(n2237), .B(\SUMB[43][2] ), .Z(n2144) );
  ND2 U3045 ( .A(\CARRYB[43][1] ), .B(\SUMB[43][2] ), .Z(n2145) );
  ND3P U3046 ( .A(n2143), .B(n2144), .C(n2145), .Z(\CARRYB[44][1] ) );
  ND2P U3047 ( .A(\SUMB[44][2] ), .B(\CARRYB[44][1] ), .Z(n2149) );
  EO3 U3048 ( .A(\CARRYB[2][2] ), .B(n301), .C(\SUMB[2][3] ), .Z(\SUMB[3][2] )
         );
  ND2 U3049 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Z(n2150) );
  ND2 U3050 ( .A(\CARRYB[2][2] ), .B(n301), .Z(n2151) );
  ND2 U3051 ( .A(\SUMB[2][3] ), .B(n301), .Z(n2152) );
  ND3 U3052 ( .A(n2150), .B(n2151), .C(n2152), .Z(\CARRYB[3][2] ) );
  EOP U3053 ( .A(n2190), .B(n2168), .Z(\SUMB[1][18] ) );
  ND3 U3054 ( .A(n2157), .B(n2158), .C(n2159), .Z(\CARRYB[13][2] ) );
  AN2P U3055 ( .A(A[30]), .B(n2321), .Z(n2208) );
  AN2P U3056 ( .A(A[34]), .B(n2321), .Z(n2213) );
  AN2P U3057 ( .A(A[32]), .B(n2321), .Z(n2211) );
  AN2P U3058 ( .A(n554), .B(n2325), .Z(n2298) );
  AN2P U3059 ( .A(A[33]), .B(n2321), .Z(n2212) );
  AN2P U3060 ( .A(A[35]), .B(n2322), .Z(n2214) );
  AN2P U3061 ( .A(A[40]), .B(n2322), .Z(n2250) );
  AN2P U3062 ( .A(A[38]), .B(n2322), .Z(n2249) );
  AN2P U3063 ( .A(A[22]), .B(n2320), .Z(n2263) );
  AN2P U3064 ( .A(A[20]), .B(n2320), .Z(n2176) );
  AN2P U3065 ( .A(n2384), .B(n2328), .Z(n2273) );
  AN2P U3066 ( .A(A[24]), .B(n2321), .Z(n2259) );
  AN2P U3067 ( .A(A[21]), .B(n2320), .Z(n2264) );
  AN2P U3068 ( .A(A[26]), .B(n2321), .Z(n2258) );
  AN2P U3069 ( .A(A[41]), .B(n2322), .Z(n2251) );
  AN2P U3070 ( .A(n2368), .B(n2328), .Z(n2289) );
  AN2P U3071 ( .A(n2376), .B(n2330), .Z(n2307) );
  ND2 U3072 ( .A(\CARRYB[41][2] ), .B(\SUMB[41][3] ), .Z(n2154) );
  ND2 U3073 ( .A(\CARRYB[41][2] ), .B(n2265), .Z(n2155) );
  ND2 U3074 ( .A(\SUMB[41][3] ), .B(n2265), .Z(n2156) );
  ND3P U3075 ( .A(n2154), .B(n2155), .C(n2156), .Z(\CARRYB[42][2] ) );
  AN2P U3076 ( .A(A[42]), .B(n2322), .Z(n2265) );
  ND2 U3077 ( .A(\CARRYB[12][2] ), .B(\SUMB[12][3] ), .Z(n2157) );
  ND2 U3078 ( .A(\CARRYB[12][2] ), .B(n2266), .Z(n2158) );
  ND2 U3079 ( .A(\SUMB[12][3] ), .B(n2266), .Z(n2159) );
  EOP U3080 ( .A(\CARRYB[47][3] ), .B(\SUMB[47][4] ), .Z(\A1[49] ) );
  EOP U3081 ( .A(\CARRYB[47][42] ), .B(\SUMB[47][43] ), .Z(\A1[88] ) );
  EOP U3082 ( .A(\CARRYB[47][23] ), .B(\SUMB[47][24] ), .Z(\A1[69] ) );
  EOP U3083 ( .A(\CARRYB[47][18] ), .B(\SUMB[47][19] ), .Z(\A1[64] ) );
  EOP U3084 ( .A(\CARRYB[47][15] ), .B(\SUMB[47][16] ), .Z(\A1[61] ) );
  EOP U3085 ( .A(\SUMB[47][29] ), .B(\CARRYB[47][28] ), .Z(\A1[74] ) );
  EOP U3086 ( .A(\CARRYB[47][29] ), .B(\SUMB[47][30] ), .Z(\A1[75] ) );
  EOP U3087 ( .A(\CARRYB[47][8] ), .B(\SUMB[47][9] ), .Z(\A1[54] ) );
  EOP U3088 ( .A(n333), .B(n2241), .Z(\SUMB[1][14] ) );
  EOP U3089 ( .A(n2236), .B(n2315), .Z(\SUMB[1][23] ) );
  EOP U3090 ( .A(n2173), .B(n2165), .Z(\SUMB[1][19] ) );
  EOP U3091 ( .A(n2205), .B(n2221), .Z(\SUMB[1][39] ) );
  AN2 U3092 ( .A(A[28]), .B(n2321), .Z(n2210) );
  AN2 U3093 ( .A(A[27]), .B(n2321), .Z(n2209) );
  IV U3094 ( .A(n346), .Z(n2327) );
  IV U3095 ( .A(n375), .Z(n2331) );
  IV U3096 ( .A(n425), .Z(n2333) );
  IV U3097 ( .A(n427), .Z(n2335) );
  IV U3098 ( .A(n425), .Z(n2334) );
  IV U3099 ( .A(n553), .Z(n2337) );
  IVDA U3100 ( .A(n578), .Y(n2339) );
  IVDA U3101 ( .A(n578), .Y(n2340) );
  IVDA U3102 ( .A(n2344), .Y(n2341) );
  IVDA U3103 ( .A(n2344), .Y(n2343) );
  IVDA U3104 ( .A(n2344), .Y(n2342) );
  IVDA U3105 ( .A(n260), .Y(n2348) );
  IVDA U3106 ( .A(n260), .Y(n2347) );
  IVDA U3107 ( .A(n2351), .Y(n2349) );
  IVDA U3108 ( .A(n2351), .Y(n2350) );
  ND2 U3109 ( .A(\CARRYB[4][6] ), .B(\SUMB[4][7] ), .Z(n2161) );
  ND2 U3110 ( .A(\CARRYB[4][6] ), .B(n448), .Z(n2162) );
  ND2 U3111 ( .A(\SUMB[4][7] ), .B(n448), .Z(n2163) );
  ND3 U3112 ( .A(n2161), .B(n2162), .C(n2163), .Z(\CARRYB[5][6] ) );
  EO U3113 ( .A(\CARRYB[47][1] ), .B(\SUMB[47][2] ), .Z(\A1[47] ) );
  EO U3114 ( .A(\CARRYB[47][33] ), .B(\SUMB[47][34] ), .Z(\A1[79] ) );
  EO U3115 ( .A(\CARRYB[47][41] ), .B(\SUMB[47][42] ), .Z(\A1[87] ) );
  EO U3116 ( .A(\CARRYB[47][40] ), .B(\SUMB[47][41] ), .Z(\A1[86] ) );
  EO U3117 ( .A(\CARRYB[47][0] ), .B(\SUMB[47][1] ), .Z(\A1[46] ) );
  EO U3118 ( .A(n331), .B(n270), .Z(\SUMB[1][20] ) );
  EO U3119 ( .A(n2191), .B(n2192), .Z(\SUMB[1][12] ) );
  EO U3120 ( .A(n2228), .B(n2231), .Z(\SUMB[1][17] ) );
  EO U3121 ( .A(n286), .B(n2194), .Z(\SUMB[1][13] ) );
  EO U3122 ( .A(n269), .B(n2218), .Z(\SUMB[1][15] ) );
  EO U3123 ( .A(n2230), .B(n2217), .Z(\SUMB[1][9] ) );
  EO U3124 ( .A(n2255), .B(n2242), .Z(\SUMB[1][6] ) );
  EO U3125 ( .A(\CARRYB[47][45] ), .B(\CARRYB[46][46] ), .Z(\A1[91] ) );
  AN2P U3126 ( .A(\ab[29][29] ), .B(n2070), .Z(n2164) );
  AN2P U3127 ( .A(\ab[19][19] ), .B(n2040), .Z(n2165) );
  AN2P U3128 ( .A(A[27]), .B(n2040), .Z(n2166) );
  AN2P U3129 ( .A(A[30]), .B(n2070), .Z(n2167) );
  AN2P U3130 ( .A(\ab[18][18] ), .B(n2040), .Z(n2168) );
  AN2P U3131 ( .A(A[31]), .B(n2117), .Z(n2170) );
  AN2P U3132 ( .A(A[29]), .B(PRODUCT[0]), .Z(n2171) );
  AN2P U3133 ( .A(\ab[36][36] ), .B(n243), .Z(n2172) );
  AN2P U3134 ( .A(A[28]), .B(A[0]), .Z(n2174) );
  AN2P U3135 ( .A(\ab[37][37] ), .B(n2070), .Z(n2175) );
  AN2P U3136 ( .A(A[25]), .B(n2040), .Z(n2177) );
  AN2P U3137 ( .A(\ab[34][34] ), .B(n2070), .Z(n2178) );
  AN2P U3138 ( .A(\ab[21][21] ), .B(n2040), .Z(n2179) );
  AN2P U3139 ( .A(\ab[11][11] ), .B(A[1]), .Z(n2180) );
  AN2P U3140 ( .A(A[33]), .B(n2040), .Z(n2181) );
  AN2P U3141 ( .A(A[26]), .B(n2117), .Z(n2182) );
  AN2P U3142 ( .A(\ab[12][12] ), .B(n2117), .Z(n2183) );
  AN2P U3143 ( .A(\ab[31][31] ), .B(n2070), .Z(n2185) );
  AN2P U3144 ( .A(\ab[28][28] ), .B(n2070), .Z(n2186) );
  AN2P U3145 ( .A(\ab[16][16] ), .B(n2070), .Z(n2187) );
  AN2P U3146 ( .A(\ab[35][35] ), .B(n2070), .Z(n2188) );
  AN2P U3147 ( .A(A[34]), .B(A[0]), .Z(n2189) );
  AN2P U3148 ( .A(A[19]), .B(PRODUCT[0]), .Z(n2190) );
  AN2P U3149 ( .A(A[12]), .B(A[1]), .Z(n2192) );
  AN2P U3150 ( .A(A[13]), .B(n2040), .Z(n2194) );
  AN2P U3151 ( .A(A[40]), .B(n2040), .Z(n2195) );
  AN2P U3152 ( .A(\ab[46][46] ), .B(n2070), .Z(n2196) );
  AN2P U3153 ( .A(A[36]), .B(n2040), .Z(n2197) );
  AN2P U3154 ( .A(A[31]), .B(n2321), .Z(n2198) );
  AN2P U3155 ( .A(A[23]), .B(n2321), .Z(n2199) );
  AN2P U3156 ( .A(\ab[45][45] ), .B(n2070), .Z(n2201) );
  AN2P U3157 ( .A(A[43]), .B(n2040), .Z(n2202) );
  AN2P U3158 ( .A(A[46]), .B(n243), .Z(n2203) );
  AN2P U3159 ( .A(A[44]), .B(A[0]), .Z(n2204) );
  AN2P U3160 ( .A(\ab[40][40] ), .B(n49), .Z(n2205) );
  AN2P U3161 ( .A(\ab[42][42] ), .B(n2040), .Z(n2206) );
  AN2P U3162 ( .A(A[25]), .B(n2321), .Z(n2207) );
  AN2P U3163 ( .A(A[19]), .B(n2320), .Z(n2215) );
  AN2P U3164 ( .A(A[18]), .B(n2320), .Z(n2216) );
  AN2P U3165 ( .A(A[9]), .B(A[1]), .Z(n2217) );
  AN2P U3166 ( .A(A[15]), .B(n2070), .Z(n2218) );
  AN2P U3167 ( .A(\ab[5][5] ), .B(A[1]), .Z(n2219) );
  AN2P U3168 ( .A(\ab[26][26] ), .B(n2040), .Z(n2220) );
  AN2P U3169 ( .A(\ab[39][39] ), .B(n2040), .Z(n2221) );
  AN2P U3170 ( .A(\ab[41][41] ), .B(n2040), .Z(n2222) );
  AN2P U3171 ( .A(\ab[22][22] ), .B(n2040), .Z(n2223) );
  AN2P U3172 ( .A(\ab[27][27] ), .B(n243), .Z(n2224) );
  AN2P U3173 ( .A(A[42]), .B(PRODUCT[0]), .Z(n2225) );
  AN2P U3174 ( .A(\ab[38][38] ), .B(n243), .Z(n2226) );
  AN2P U3175 ( .A(A[18]), .B(PRODUCT[0]), .Z(n2228) );
  AN2P U3176 ( .A(\ab[9][9] ), .B(A[0]), .Z(n2229) );
  AN2P U3177 ( .A(\ab[10][10] ), .B(A[0]), .Z(n2230) );
  AN2P U3178 ( .A(\ab[17][17] ), .B(A[1]), .Z(n2231) );
  AN2P U3179 ( .A(A[8]), .B(A[1]), .Z(n2232) );
  AN2P U3180 ( .A(A[10]), .B(n2040), .Z(n2234) );
  AN2P U3181 ( .A(A[24]), .B(n2117), .Z(n2236) );
  AN2P U3182 ( .A(\ab[44][44] ), .B(n2070), .Z(n2237) );
  EO U3183 ( .A(n2189), .B(n2181), .Z(\SUMB[1][33] ) );
  AN2P U3184 ( .A(A[29]), .B(n2321), .Z(n2238) );
  AN2P U3185 ( .A(A[41]), .B(A[0]), .Z(n2239) );
  AN2P U3186 ( .A(\ab[24][24] ), .B(n2070), .Z(n2240) );
  AN2P U3187 ( .A(\ab[14][14] ), .B(n2070), .Z(n2241) );
  AN2P U3188 ( .A(A[6]), .B(A[1]), .Z(n2242) );
  AN2P U3189 ( .A(\ab[45][45] ), .B(n49), .Z(n2243) );
  AN2P U3190 ( .A(\ab[7][7] ), .B(A[1]), .Z(n2244) );
  AN2P U3191 ( .A(n2040), .B(A[47]), .Z(n2245) );
  AN2P U3192 ( .A(n49), .B(A[47]), .Z(n2246) );
  AN2P U3193 ( .A(A[45]), .B(n2322), .Z(n2247) );
  AN2P U3194 ( .A(A[44]), .B(n2322), .Z(n2248) );
  AN2P U3195 ( .A(A[43]), .B(n2322), .Z(n2252) );
  AN2P U3196 ( .A(\ab[4][4] ), .B(A[1]), .Z(n2253) );
  AN2P U3197 ( .A(A[9]), .B(n2319), .Z(n2254) );
  AN2P U3198 ( .A(A[5]), .B(A[0]), .Z(n2256) );
  AN2P U3199 ( .A(A[46]), .B(n2322), .Z(n2257) );
  AN2P U3200 ( .A(A[36]), .B(n2322), .Z(n2260) );
  AN2P U3201 ( .A(A[39]), .B(n2322), .Z(n2261) );
  AN2P U3202 ( .A(A[17]), .B(n2320), .Z(n2262) );
  AN2P U3203 ( .A(A[13]), .B(n2320), .Z(n2266) );
  AN2P U3204 ( .A(n376), .B(n2319), .Z(n2267) );
  EO U3205 ( .A(n326), .B(n2423), .Z(\SUMB[1][3] ) );
  AN2P U3206 ( .A(A[31]), .B(n2327), .Z(n2268) );
  AN2P U3207 ( .A(n247), .B(n2325), .Z(n2269) );
  AN2P U3208 ( .A(A[29]), .B(n2326), .Z(n2270) );
  AN2P U3209 ( .A(A[23]), .B(n2326), .Z(n2271) );
  AN2P U3210 ( .A(n250), .B(n2326), .Z(n2272) );
  AN2P U3211 ( .A(n2373), .B(n2327), .Z(n2274) );
  AN2P U3212 ( .A(n2394), .B(n2328), .Z(n2275) );
  AN2P U3213 ( .A(n735), .B(n2327), .Z(n2276) );
  AN2P U3214 ( .A(A[36]), .B(n2327), .Z(n2277) );
  AN2P U3215 ( .A(n259), .B(n2328), .Z(n2278) );
  AN2P U3216 ( .A(n728), .B(n2327), .Z(n2279) );
  AN2P U3217 ( .A(n245), .B(n2325), .Z(n2280) );
  AN2P U3218 ( .A(n2383), .B(n2330), .Z(n2281) );
  AN2P U3219 ( .A(A[46]), .B(n2327), .Z(n2282) );
  AN2P U3220 ( .A(n2390), .B(n2325), .Z(n2283) );
  AN2P U3221 ( .A(A[44]), .B(n2326), .Z(n2285) );
  AN2P U3222 ( .A(A[41]), .B(n2328), .Z(n2286) );
  AN2P U3223 ( .A(n646), .B(n2326), .Z(n2287) );
  AN2P U3224 ( .A(A[26]), .B(n2328), .Z(n2288) );
  AN2P U3225 ( .A(A[45]), .B(n2327), .Z(n2290) );
  AN2P U3226 ( .A(n300), .B(n2326), .Z(n2291) );
  AN2P U3227 ( .A(n732), .B(n2326), .Z(n2292) );
  AN2P U3228 ( .A(n730), .B(n2326), .Z(n2293) );
  AN2P U3229 ( .A(n2406), .B(n2328), .Z(n2294) );
  AN2P U3230 ( .A(n652), .B(n2327), .Z(n2295) );
  AN2P U3231 ( .A(n650), .B(n2325), .Z(n2296) );
  AN2P U3232 ( .A(n737), .B(n2325), .Z(n2297) );
  AN2P U3233 ( .A(n2380), .B(n2330), .Z(n2299) );
  AN2P U3234 ( .A(n254), .B(n2330), .Z(n2300) );
  AN2P U3235 ( .A(n2359), .B(n349), .Z(n2301) );
  AN2P U3236 ( .A(n2361), .B(n349), .Z(n2302) );
  AN2P U3237 ( .A(n2397), .B(n2330), .Z(n2303) );
  AN2P U3238 ( .A(n2387), .B(n2330), .Z(n2304) );
  AN2P U3239 ( .A(A[39]), .B(n2328), .Z(n2305) );
  AN2P U3240 ( .A(n2393), .B(n2330), .Z(n2306) );
  AN2P U3241 ( .A(n2357), .B(n349), .Z(n2308) );
  AN2P U3242 ( .A(n2372), .B(n2330), .Z(n2309) );
  AN2P U3243 ( .A(n2332), .B(n2325), .Z(n2310) );
  EO U3244 ( .A(\CARRYB[47][46] ), .B(n2421), .Z(\A1[92] ) );
  EO U3245 ( .A(n2424), .B(n2426), .Z(\SUMB[1][2] ) );
  IV U3246 ( .A(n346), .Z(n2328) );
  IV U3247 ( .A(n346), .Z(n2326) );
  IV U3248 ( .A(n346), .Z(n2325) );
  IV U3249 ( .A(n348), .Z(n2330) );
  IV U3250 ( .A(n348), .Z(n2329) );
  IV U3251 ( .A(n375), .Z(n2332) );
  IVDA U3252 ( .A(n553), .Y(n2338) );
  IVDA U3253 ( .A(n2388), .Y(n2387) );
  IVDA U3254 ( .A(n2391), .Y(n2390) );
  IVDA U3255 ( .A(n264), .Y(n2345) );
  IVDA U3256 ( .A(n645), .Y(n2346) );
  IVDA U3257 ( .A(n729), .Y(n2363) );
  IVDA U3258 ( .A(n731), .Y(n2365) );
  IVDA U3259 ( .A(n2381), .Y(n2380) );
  IVDA U3260 ( .A(n734), .Y(n2397) );
  IVDA U3261 ( .A(n2385), .Y(n2384) );
  IVDA U3262 ( .A(n2395), .Y(n2394) );
  IVDA U3263 ( .A(n2403), .Y(n2402) );
  IVDA U3264 ( .A(n255), .Y(n2420) );
  IVDA U3265 ( .A(n2407), .Y(n2406) );
  IVDA U3266 ( .A(n279), .Y(n2417) );
  IVP U3267 ( .A(n2354), .Z(n2352) );
  IVDA U3268 ( .A(n727), .Y(n2355) );
  IVP U3269 ( .A(n2354), .Z(n2353) );
  IVDA U3270 ( .A(n258), .Y(n2356) );
  IVDA U3271 ( .A(n244), .Y(n2360) );
  IVDA U3272 ( .A(n258), .Y(n2357) );
  IVDA U3273 ( .A(n249), .Y(n2359) );
  IVDA U3274 ( .A(n729), .Y(n2362) );
  IVDA U3275 ( .A(n244), .Y(n2361) );
  IVDA U3276 ( .A(n731), .Y(n2364) );
  IVDA U3277 ( .A(n277), .Y(n2366) );
  IVDA U3278 ( .A(n266), .Y(n2368) );
  IVDA U3279 ( .A(n277), .Y(n2367) );
  IVDA U3280 ( .A(n2385), .Y(n2383) );
  IVDA U3281 ( .A(n2381), .Y(n2379) );
  IVDA U3282 ( .A(n2377), .Y(n2376) );
  IVDA U3283 ( .A(n2374), .Y(n2373) );
  IVDA U3284 ( .A(n651), .Y(n2412) );
  IVDA U3285 ( .A(n2410), .Y(n2409) );
  IVDA U3286 ( .A(n2395), .Y(n2393) );
  IVDA U3287 ( .A(n246), .Y(n2369) );
  IVDA U3288 ( .A(n649), .Y(n2414) );
  IVDA U3289 ( .A(n736), .Y(n2415) );
  IVDA U3290 ( .A(n262), .Y(n2418) );
  IVDA U3291 ( .A(n255), .Y(n2419) );
  IVDA U3292 ( .A(n2407), .Y(n2405) );
  IVDA U3293 ( .A(n2403), .Y(n2401) );
  IVDA U3294 ( .A(n299), .Y(n2398) );
  IVDA U3295 ( .A(n734), .Y(n2396) );
  IVDA U3296 ( .A(n2371), .Y(n2370) );
  IVDA U3297 ( .A(n279), .Y(n2416) );
  IVDA U3298 ( .A(n2374), .Y(n2372) );
  IVDA U3299 ( .A(n2377), .Y(n2375) );
  IVDA U3300 ( .A(n2381), .Y(n2378) );
  IVDA U3301 ( .A(n2385), .Y(n2382) );
  IVDA U3302 ( .A(n2388), .Y(n2386) );
  IVDA U3303 ( .A(n2391), .Y(n2389) );
  IVDA U3304 ( .A(n2395), .Y(n2392) );
  IVDA U3305 ( .A(n2410), .Y(n2408) );
  IVDA U3306 ( .A(n253), .Y(n2399) );
  IVDA U3307 ( .A(n651), .Y(n2411) );
  IVDA U3308 ( .A(n2407), .Y(n2404) );
  IVDA U3309 ( .A(n649), .Y(n2413) );
  IVDA U3310 ( .A(n2403), .Y(n2400) );
  AN2P U3311 ( .A(\CARRYB[47][14] ), .B(\SUMB[47][15] ), .Z(\A2[61] ) );
  AN2P U3312 ( .A(\CARRYB[47][16] ), .B(\SUMB[47][17] ), .Z(\A2[63] ) );
  EOP U3313 ( .A(\CARRYB[47][16] ), .B(\SUMB[47][17] ), .Z(\A1[62] ) );
  AN2P U3314 ( .A(\CARRYB[47][19] ), .B(\SUMB[47][20] ), .Z(\A2[66] ) );
  EOP U3315 ( .A(\CARRYB[47][19] ), .B(\SUMB[47][20] ), .Z(\A1[65] ) );
  AN2P U3316 ( .A(\CARRYB[47][20] ), .B(\SUMB[47][21] ), .Z(\A2[67] ) );
  EOP U3317 ( .A(\SUMB[47][21] ), .B(\CARRYB[47][20] ), .Z(\A1[66] ) );
  AN2P U3318 ( .A(\CARRYB[47][21] ), .B(\SUMB[47][22] ), .Z(\A2[68] ) );
  AN2P U3319 ( .A(\CARRYB[47][22] ), .B(\SUMB[47][23] ), .Z(\A2[69] ) );
  AN2P U3320 ( .A(\CARRYB[47][23] ), .B(\SUMB[47][24] ), .Z(\A2[70] ) );
  EOP U3321 ( .A(\CARRYB[47][24] ), .B(\SUMB[47][25] ), .Z(\A1[70] ) );
  AN2P U3322 ( .A(\CARRYB[47][26] ), .B(\SUMB[47][27] ), .Z(\A2[73] ) );
  EOP U3323 ( .A(\CARRYB[47][26] ), .B(\SUMB[47][27] ), .Z(\A1[72] ) );
  AN2P U3324 ( .A(\CARRYB[47][28] ), .B(\SUMB[47][29] ), .Z(\A2[75] ) );
  AN2P U3325 ( .A(\CARRYB[47][30] ), .B(\SUMB[47][31] ), .Z(\A2[77] ) );
  AN2P U3326 ( .A(\CARRYB[47][34] ), .B(\SUMB[47][35] ), .Z(\A2[81] ) );
  EOP U3327 ( .A(\CARRYB[47][34] ), .B(\SUMB[47][35] ), .Z(\A1[80] ) );
  AN2P U3328 ( .A(\CARRYB[47][36] ), .B(\SUMB[47][37] ), .Z(\A2[83] ) );
  EOP U3329 ( .A(\CARRYB[47][36] ), .B(\SUMB[47][37] ), .Z(\A1[82] ) );
  AN2P U3330 ( .A(\CARRYB[47][37] ), .B(\SUMB[47][38] ), .Z(\A2[84] ) );
  EOP U3331 ( .A(\CARRYB[47][37] ), .B(\SUMB[47][38] ), .Z(\A1[83] ) );
  AN2P U3332 ( .A(\CARRYB[47][38] ), .B(\SUMB[47][39] ), .Z(\A2[85] ) );
  EOP U3333 ( .A(\CARRYB[47][38] ), .B(\SUMB[47][39] ), .Z(\A1[84] ) );
  AN2P U3334 ( .A(\CARRYB[47][39] ), .B(\SUMB[47][40] ), .Z(\A2[86] ) );
  EOP U3335 ( .A(\CARRYB[47][39] ), .B(\SUMB[47][40] ), .Z(\A1[85] ) );
  AN2P U3336 ( .A(\CARRYB[47][42] ), .B(\SUMB[47][43] ), .Z(\A2[89] ) );
  AN2P U3337 ( .A(\CARRYB[47][43] ), .B(\SUMB[47][44] ), .Z(\A2[90] ) );
  AN2P U3338 ( .A(\CARRYB[47][44] ), .B(\SUMB[47][45] ), .Z(\A2[91] ) );
  AN2P U3339 ( .A(\CARRYB[47][45] ), .B(\CARRYB[46][46] ), .Z(\A2[92] ) );
  AN2P U3340 ( .A(n2426), .B(n2424), .Z(\CARRYB[1][2] ) );
  AN2P U3341 ( .A(n2423), .B(n326), .Z(\CARRYB[1][3] ) );
  AN2P U3342 ( .A(n2253), .B(n2256), .Z(\CARRYB[1][4] ) );
  AN2P U3343 ( .A(n2219), .B(n285), .Z(\CARRYB[1][5] ) );
  AN2P U3344 ( .A(n2242), .B(n2255), .Z(\CARRYB[1][6] ) );
  AN2P U3345 ( .A(n2244), .B(n327), .Z(\CARRYB[1][7] ) );
  AN2P U3346 ( .A(n2217), .B(n2230), .Z(\CARRYB[1][9] ) );
  AN2P U3347 ( .A(n2194), .B(n286), .Z(\CARRYB[1][13] ) );
  EOP U3348 ( .A(n334), .B(n2233), .Z(\SUMB[1][38] ) );
  AN2P U3349 ( .A(n2192), .B(n2191), .Z(\CARRYB[1][12] ) );
  AN2P U3350 ( .A(\CARRYB[47][11] ), .B(\SUMB[47][12] ), .Z(\A2[58] ) );
  EOP U3351 ( .A(\SUMB[47][12] ), .B(\CARRYB[47][11] ), .Z(\A1[57] ) );
  AN2P U3352 ( .A(n2232), .B(n2229), .Z(\CARRYB[1][8] ) );
  AN2P U3353 ( .A(\CARRYB[47][18] ), .B(\SUMB[47][19] ), .Z(\A2[65] ) );
  AN2P U3354 ( .A(\CARRYB[47][31] ), .B(\SUMB[47][32] ), .Z(\A2[78] ) );
  AN2P U3355 ( .A(n2186), .B(n2171), .Z(\CARRYB[1][28] ) );
  AN2P U3356 ( .A(\CARRYB[47][40] ), .B(\SUMB[47][41] ), .Z(\A2[87] ) );
  EOP U3357 ( .A(\SUMB[47][11] ), .B(\CARRYB[47][10] ), .Z(\A1[56] ) );
  AN2P U3358 ( .A(\CARRYB[47][46] ), .B(n2421), .Z(\A2[93] ) );
  AN2P U3359 ( .A(n270), .B(n331), .Z(\CARRYB[1][20] ) );
  AN2P U3360 ( .A(n2197), .B(n320), .Z(\CARRYB[1][36] ) );
  AN2P U3361 ( .A(\CARRYB[47][29] ), .B(\SUMB[47][30] ), .Z(\A2[76] ) );
  AN2P U3362 ( .A(\CARRYB[47][4] ), .B(\SUMB[47][5] ), .Z(\A2[51] ) );
  EOP U3363 ( .A(\SUMB[47][5] ), .B(\CARRYB[47][4] ), .Z(\A1[50] ) );
  AN2P U3364 ( .A(\CARRYB[47][9] ), .B(\SUMB[47][10] ), .Z(\A2[56] ) );
  EOP U3365 ( .A(\CARRYB[47][9] ), .B(\SUMB[47][10] ), .Z(\A1[55] ) );
  AN2P U3366 ( .A(\CARRYB[47][33] ), .B(\SUMB[47][34] ), .Z(\A2[80] ) );
  AN2P U3367 ( .A(\CARRYB[47][6] ), .B(\SUMB[47][7] ), .Z(\A2[53] ) );
  EOP U3368 ( .A(\CARRYB[47][6] ), .B(\SUMB[47][7] ), .Z(\A1[52] ) );
  AN2P U3369 ( .A(n2195), .B(n2239), .Z(\CARRYB[1][40] ) );
  AN2P U3370 ( .A(\CARRYB[47][7] ), .B(\SUMB[47][8] ), .Z(\A2[54] ) );
  EOP U3371 ( .A(\CARRYB[47][7] ), .B(\SUMB[47][8] ), .Z(\A1[53] ) );
  AN2P U3372 ( .A(\CARRYB[47][5] ), .B(\SUMB[47][6] ), .Z(\A2[52] ) );
  EOP U3373 ( .A(\CARRYB[47][5] ), .B(\SUMB[47][6] ), .Z(\A1[51] ) );
  AN2P U3374 ( .A(\CARRYB[47][25] ), .B(\SUMB[47][26] ), .Z(\A2[72] ) );
  EOP U3375 ( .A(\CARRYB[47][25] ), .B(\SUMB[47][26] ), .Z(\A1[71] ) );
  AN2P U3376 ( .A(\CARRYB[47][17] ), .B(\SUMB[47][18] ), .Z(\A2[64] ) );
  EOP U3377 ( .A(\SUMB[47][18] ), .B(\CARRYB[47][17] ), .Z(\A1[63] ) );
  AN2P U3378 ( .A(\CARRYB[47][3] ), .B(\SUMB[47][4] ), .Z(\A2[50] ) );
  AN2P U3379 ( .A(n2177), .B(n2182), .Z(\CARRYB[1][25] ) );
  AN2P U3380 ( .A(\CARRYB[47][32] ), .B(\SUMB[47][33] ), .Z(\A2[79] ) );
  AN2P U3381 ( .A(\CARRYB[47][8] ), .B(\SUMB[47][9] ), .Z(\A2[55] ) );
  AN2P U3382 ( .A(\CARRYB[47][13] ), .B(\SUMB[47][14] ), .Z(\A2[60] ) );
  EOP U3383 ( .A(\CARRYB[47][13] ), .B(\SUMB[47][14] ), .Z(\A1[59] ) );
  AN2P U3384 ( .A(\CARRYB[47][12] ), .B(\SUMB[47][13] ), .Z(\A2[59] ) );
  EOP U3385 ( .A(\CARRYB[47][12] ), .B(\SUMB[47][13] ), .Z(\A1[58] ) );
  AN2P U3386 ( .A(\CARRYB[47][2] ), .B(\SUMB[47][3] ), .Z(\A2[49] ) );
  AN2P U3387 ( .A(\CARRYB[47][27] ), .B(\SUMB[47][28] ), .Z(\A2[74] ) );
  EOP U3388 ( .A(\CARRYB[47][27] ), .B(\SUMB[47][28] ), .Z(\A1[73] ) );
  AN2P U3389 ( .A(n2218), .B(n269), .Z(\CARRYB[1][15] ) );
  AN2P U3390 ( .A(n2315), .B(n2236), .Z(\CARRYB[1][23] ) );
  AN2P U3391 ( .A(n2181), .B(n2189), .Z(\CARRYB[1][33] ) );
  AN2P U3392 ( .A(n2178), .B(n2184), .Z(\CARRYB[1][34] ) );
  AN2P U3393 ( .A(n2223), .B(n2227), .Z(\CARRYB[1][22] ) );
  AN2P U3394 ( .A(n2231), .B(n2228), .Z(\CARRYB[1][17] ) );
  AN2P U3395 ( .A(n2234), .B(n289), .Z(\CARRYB[1][10] ) );
  AN2P U3396 ( .A(n2185), .B(n332), .Z(\CARRYB[1][31] ) );
  AN2P U3397 ( .A(\CARRYB[47][35] ), .B(\SUMB[47][36] ), .Z(\A2[82] ) );
  EOP U3398 ( .A(\CARRYB[47][35] ), .B(\SUMB[47][36] ), .Z(\A1[81] ) );
  AN2P U3399 ( .A(n2201), .B(n2203), .Z(\CARRYB[1][45] ) );
  AN2P U3400 ( .A(\CARRYB[47][15] ), .B(\SUMB[47][16] ), .Z(\A2[62] ) );
  NR2 U3401 ( .A(n2391), .B(n257), .Z(n2311) );
  AN2P U3402 ( .A(n2392), .B(n2117), .Z(n2313) );
  AN2P U3403 ( .A(\ab[23][23] ), .B(n2040), .Z(n2315) );
  IVDA U3404 ( .A(n249), .Y(n2358) );
  AN2 U3405 ( .A(n1350), .B(A[0]), .Z(\ab[1][0] ) );
  AN2 U3406 ( .A(n2323), .B(n2040), .Z(n2426) );
  IVP U3407 ( .A(n2324), .Z(n2323) );
  AN2 U3409 ( .A(n2421), .B(n2337), .Z(\ab[9][47] ) );
  AN2 U3410 ( .A(n2421), .B(n2336), .Z(\ab[8][47] ) );
  AN2 U3411 ( .A(n256), .B(n2337), .Z(\ab[9][46] ) );
  AN2 U3412 ( .A(n256), .B(\ab[47][47] ), .Z(\CARRYB[47][46] ) );
  AN2 U3413 ( .A(n263), .B(n2337), .Z(\ab[9][45] ) );
  AN2 U3414 ( .A(n263), .B(n2421), .Z(\ab[47][45] ) );
  AN2 U3415 ( .A(n263), .B(n256), .Z(\ab[46][45] ) );
  AN2 U3416 ( .A(n280), .B(n2337), .Z(\ab[9][44] ) );
  AN2 U3417 ( .A(n280), .B(n2421), .Z(\ab[47][44] ) );
  AN2 U3418 ( .A(n280), .B(n256), .Z(\ab[46][44] ) );
  AN2 U3419 ( .A(n280), .B(n263), .Z(\ab[45][44] ) );
  AN2 U3420 ( .A(n737), .B(\ab[47][47] ), .Z(\ab[47][43] ) );
  AN2 U3421 ( .A(n737), .B(n256), .Z(\ab[46][43] ) );
  AN2 U3422 ( .A(n737), .B(n263), .Z(\ab[45][43] ) );
  AN2 U3423 ( .A(n737), .B(n280), .Z(\ab[44][43] ) );
  AN2 U3424 ( .A(n2413), .B(n2421), .Z(\ab[47][42] ) );
  AN2 U3425 ( .A(n2413), .B(n256), .Z(\ab[46][42] ) );
  AN2 U3426 ( .A(n2413), .B(n263), .Z(\ab[45][42] ) );
  AN2 U3427 ( .A(n2413), .B(n280), .Z(\ab[44][42] ) );
  AN2 U3428 ( .A(n2413), .B(n737), .Z(\ab[43][42] ) );
  AN2 U3429 ( .A(n316), .B(n2421), .Z(\ab[47][41] ) );
  AN2 U3430 ( .A(n316), .B(n256), .Z(\ab[46][41] ) );
  AN2 U3431 ( .A(n316), .B(n263), .Z(\ab[45][41] ) );
  AN2 U3432 ( .A(n316), .B(n280), .Z(\ab[44][41] ) );
  AN2 U3433 ( .A(n316), .B(n737), .Z(\ab[43][41] ) );
  AN2 U3434 ( .A(n316), .B(n2413), .Z(\ab[42][41] ) );
  AN2 U3435 ( .A(n2411), .B(\ab[47][47] ), .Z(\ab[47][40] ) );
  AN2 U3436 ( .A(n2411), .B(n256), .Z(\ab[46][40] ) );
  AN2 U3437 ( .A(n2411), .B(n263), .Z(\ab[45][40] ) );
  AN2 U3438 ( .A(n2411), .B(n280), .Z(\ab[44][40] ) );
  AN2 U3439 ( .A(n2411), .B(n737), .Z(\ab[43][40] ) );
  AN2 U3440 ( .A(n2411), .B(n2413), .Z(\ab[42][40] ) );
  AN2 U3441 ( .A(n2411), .B(n316), .Z(\ab[41][40] ) );
  AN2 U3442 ( .A(n2408), .B(n2421), .Z(\ab[47][39] ) );
  AN2 U3443 ( .A(n2408), .B(n256), .Z(\ab[46][39] ) );
  AN2 U3444 ( .A(n2408), .B(n263), .Z(\ab[45][39] ) );
  AN2 U3445 ( .A(n2408), .B(n280), .Z(\ab[44][39] ) );
  AN2 U3446 ( .A(n2408), .B(n737), .Z(\ab[43][39] ) );
  AN2 U3447 ( .A(n2408), .B(n2413), .Z(\ab[42][39] ) );
  AN2 U3448 ( .A(n2408), .B(n316), .Z(\ab[41][39] ) );
  AN2 U3449 ( .A(n2408), .B(n2411), .Z(\ab[40][39] ) );
  AN2 U3450 ( .A(n2404), .B(n2421), .Z(\ab[47][38] ) );
  AN2 U3451 ( .A(n2404), .B(n256), .Z(\ab[46][38] ) );
  AN2 U3452 ( .A(n2404), .B(n263), .Z(\ab[45][38] ) );
  AN2 U3453 ( .A(n2404), .B(n280), .Z(\ab[44][38] ) );
  AN2 U3454 ( .A(n2404), .B(n737), .Z(\ab[43][38] ) );
  AN2 U3455 ( .A(n2404), .B(n2413), .Z(\ab[42][38] ) );
  AN2 U3456 ( .A(n2404), .B(n316), .Z(\ab[41][38] ) );
  AN2 U3457 ( .A(n2404), .B(n2411), .Z(\ab[40][38] ) );
  AN2 U3458 ( .A(n2404), .B(n2408), .Z(\ab[39][38] ) );
  AN2 U3459 ( .A(n2400), .B(\ab[47][47] ), .Z(\ab[47][37] ) );
  AN2 U3460 ( .A(n2400), .B(n256), .Z(\ab[46][37] ) );
  AN2 U3461 ( .A(n2400), .B(n263), .Z(\ab[45][37] ) );
  AN2 U3462 ( .A(n2400), .B(n280), .Z(\ab[44][37] ) );
  AN2 U3463 ( .A(n2400), .B(n737), .Z(\ab[43][37] ) );
  AN2 U3464 ( .A(n2400), .B(n2413), .Z(\ab[42][37] ) );
  AN2 U3465 ( .A(n2400), .B(n316), .Z(\ab[41][37] ) );
  AN2 U3466 ( .A(n2400), .B(n2411), .Z(\ab[40][37] ) );
  AN2 U3467 ( .A(n2400), .B(n2408), .Z(\ab[39][37] ) );
  AN2 U3468 ( .A(n2400), .B(n2404), .Z(\ab[38][37] ) );
  AN2 U3469 ( .A(n2399), .B(n2421), .Z(\ab[47][36] ) );
  AN2 U3470 ( .A(n2399), .B(n2419), .Z(\ab[46][36] ) );
  AN2 U3471 ( .A(n2399), .B(n2418), .Z(\ab[45][36] ) );
  AN2 U3472 ( .A(n2399), .B(n2416), .Z(\ab[44][36] ) );
  AN2 U3473 ( .A(n2399), .B(n737), .Z(\ab[43][36] ) );
  AN2 U3474 ( .A(n2399), .B(n2413), .Z(\ab[42][36] ) );
  AN2 U3475 ( .A(n2399), .B(n316), .Z(\ab[41][36] ) );
  AN2 U3476 ( .A(n2399), .B(n2411), .Z(\ab[40][36] ) );
  AN2 U3477 ( .A(n2399), .B(n2408), .Z(\ab[39][36] ) );
  AN2 U3478 ( .A(n2399), .B(n2404), .Z(\ab[38][36] ) );
  AN2 U3479 ( .A(n2399), .B(n2400), .Z(\ab[37][36] ) );
  AN2 U3480 ( .A(n2398), .B(n2421), .Z(\ab[47][35] ) );
  AN2 U3481 ( .A(n300), .B(n2419), .Z(\ab[46][35] ) );
  AN2 U3482 ( .A(n300), .B(n2418), .Z(\ab[45][35] ) );
  AN2 U3483 ( .A(n2398), .B(n2416), .Z(\ab[44][35] ) );
  AN2 U3484 ( .A(n300), .B(n2415), .Z(\ab[43][35] ) );
  AN2 U3485 ( .A(n300), .B(n2414), .Z(\ab[42][35] ) );
  AN2 U3486 ( .A(n2398), .B(n316), .Z(\ab[41][35] ) );
  AN2 U3487 ( .A(n2398), .B(n2412), .Z(\ab[40][35] ) );
  AN2 U3488 ( .A(n2398), .B(n2409), .Z(\ab[39][35] ) );
  AN2 U3489 ( .A(n2398), .B(n2405), .Z(\ab[38][35] ) );
  AN2 U3490 ( .A(n2398), .B(n2401), .Z(\ab[37][35] ) );
  AN2 U3491 ( .A(n2398), .B(n254), .Z(\ab[36][35] ) );
  AN2 U3492 ( .A(n735), .B(\ab[47][47] ), .Z(\ab[47][34] ) );
  AN2 U3493 ( .A(n735), .B(n2419), .Z(\ab[46][34] ) );
  AN2 U3494 ( .A(n735), .B(n2418), .Z(\ab[45][34] ) );
  AN2 U3495 ( .A(n735), .B(n2416), .Z(\ab[44][34] ) );
  AN2 U3496 ( .A(n735), .B(n2415), .Z(\ab[43][34] ) );
  AN2 U3497 ( .A(n735), .B(n2414), .Z(\ab[42][34] ) );
  AN2 U3498 ( .A(n735), .B(n316), .Z(\ab[41][34] ) );
  AN2 U3499 ( .A(n735), .B(n2412), .Z(\ab[40][34] ) );
  AN2 U3500 ( .A(n735), .B(n2409), .Z(\ab[39][34] ) );
  AN2 U3501 ( .A(n735), .B(n2405), .Z(\ab[38][34] ) );
  AN2 U3502 ( .A(n735), .B(n2401), .Z(\ab[37][34] ) );
  AN2 U3503 ( .A(n2396), .B(n254), .Z(\ab[36][34] ) );
  AN2 U3504 ( .A(n2396), .B(n2398), .Z(\ab[35][34] ) );
  AN2 U3505 ( .A(n2392), .B(n2421), .Z(\ab[47][33] ) );
  AN2 U3506 ( .A(n2392), .B(n2419), .Z(\ab[46][33] ) );
  AN2 U3507 ( .A(n2392), .B(n2418), .Z(\ab[45][33] ) );
  AN2 U3508 ( .A(n2392), .B(n2416), .Z(\ab[44][33] ) );
  AN2 U3509 ( .A(n2392), .B(n2415), .Z(\ab[43][33] ) );
  AN2 U3510 ( .A(n2392), .B(n2414), .Z(\ab[42][33] ) );
  AN2 U3511 ( .A(n2392), .B(n316), .Z(\ab[41][33] ) );
  AN2 U3512 ( .A(n2392), .B(n2412), .Z(\ab[40][33] ) );
  AN2 U3513 ( .A(n2392), .B(n2409), .Z(\ab[39][33] ) );
  AN2 U3514 ( .A(n2392), .B(n2405), .Z(\ab[38][33] ) );
  AN2 U3515 ( .A(n2392), .B(n2401), .Z(\ab[37][33] ) );
  AN2 U3516 ( .A(n2393), .B(n254), .Z(\ab[36][33] ) );
  AN2 U3517 ( .A(n2393), .B(n2398), .Z(\ab[35][33] ) );
  AN2 U3518 ( .A(n2393), .B(n2396), .Z(\ab[34][33] ) );
  AN2 U3519 ( .A(n2389), .B(n2421), .Z(\ab[47][32] ) );
  AN2 U3520 ( .A(n2389), .B(n2419), .Z(\ab[46][32] ) );
  AN2 U3521 ( .A(n2389), .B(n2418), .Z(\ab[45][32] ) );
  AN2 U3522 ( .A(n2389), .B(n2416), .Z(\ab[44][32] ) );
  AN2 U3523 ( .A(n2389), .B(n2415), .Z(\ab[43][32] ) );
  AN2 U3524 ( .A(n2389), .B(n2414), .Z(\ab[42][32] ) );
  AN2 U3525 ( .A(n2389), .B(n316), .Z(\ab[41][32] ) );
  AN2 U3526 ( .A(n2389), .B(n2412), .Z(\ab[40][32] ) );
  AN2 U3527 ( .A(n2389), .B(n2409), .Z(\ab[39][32] ) );
  AN2 U3528 ( .A(n2389), .B(n2405), .Z(\ab[38][32] ) );
  AN2 U3529 ( .A(n2389), .B(n2401), .Z(\ab[37][32] ) );
  AN2 U3530 ( .A(n2389), .B(n254), .Z(\ab[36][32] ) );
  AN2 U3531 ( .A(A[32]), .B(n2398), .Z(\ab[35][32] ) );
  AN2 U3532 ( .A(A[32]), .B(n2396), .Z(\ab[34][32] ) );
  AN2 U3533 ( .A(n2389), .B(n2393), .Z(\ab[33][32] ) );
  AN2 U3534 ( .A(n2386), .B(\ab[47][47] ), .Z(\ab[47][31] ) );
  AN2 U3535 ( .A(n2386), .B(n2419), .Z(\ab[46][31] ) );
  AN2 U3536 ( .A(n2386), .B(n2418), .Z(\ab[45][31] ) );
  AN2 U3537 ( .A(n2386), .B(n2416), .Z(\ab[44][31] ) );
  AN2 U3538 ( .A(n2386), .B(n2415), .Z(\ab[43][31] ) );
  AN2 U3539 ( .A(n2386), .B(n2414), .Z(\ab[42][31] ) );
  AN2 U3540 ( .A(n2386), .B(n316), .Z(\ab[41][31] ) );
  AN2 U3541 ( .A(n2386), .B(n2412), .Z(\ab[40][31] ) );
  AN2 U3542 ( .A(n2386), .B(n2409), .Z(\ab[39][31] ) );
  AN2 U3543 ( .A(n2386), .B(n2405), .Z(\ab[38][31] ) );
  AN2 U3544 ( .A(n2386), .B(n2401), .Z(\ab[37][31] ) );
  AN2 U3545 ( .A(A[31]), .B(n254), .Z(\ab[36][31] ) );
  AN2 U3546 ( .A(A[31]), .B(n2398), .Z(\ab[35][31] ) );
  AN2 U3547 ( .A(A[31]), .B(n2396), .Z(\ab[34][31] ) );
  AN2 U3548 ( .A(n2386), .B(n2393), .Z(\ab[33][31] ) );
  AN2 U3549 ( .A(n2386), .B(n2389), .Z(\ab[32][31] ) );
  AN2 U3550 ( .A(n2382), .B(n2421), .Z(\ab[47][30] ) );
  AN2 U3551 ( .A(n2382), .B(n2419), .Z(\ab[46][30] ) );
  AN2 U3552 ( .A(n2382), .B(n2418), .Z(\ab[45][30] ) );
  AN2 U3553 ( .A(n2382), .B(n2416), .Z(\ab[44][30] ) );
  AN2 U3554 ( .A(n2382), .B(n2415), .Z(\ab[43][30] ) );
  AN2 U3555 ( .A(n2382), .B(n2414), .Z(\ab[42][30] ) );
  AN2 U3556 ( .A(n2382), .B(n316), .Z(\ab[41][30] ) );
  AN2 U3557 ( .A(n2382), .B(n2412), .Z(\ab[40][30] ) );
  AN2 U3558 ( .A(n2382), .B(n2409), .Z(\ab[39][30] ) );
  AN2 U3559 ( .A(n2382), .B(n2405), .Z(\ab[38][30] ) );
  AN2 U3560 ( .A(n2382), .B(n2401), .Z(\ab[37][30] ) );
  AN2 U3561 ( .A(n2383), .B(n254), .Z(\ab[36][30] ) );
  AN2 U3562 ( .A(n2383), .B(n2398), .Z(\ab[35][30] ) );
  AN2 U3563 ( .A(n2383), .B(n2396), .Z(\ab[34][30] ) );
  AN2 U3564 ( .A(n2383), .B(n2393), .Z(\ab[33][30] ) );
  AN2 U3565 ( .A(n2383), .B(n2389), .Z(\ab[32][30] ) );
  AN2 U3566 ( .A(n2383), .B(n2386), .Z(\ab[31][30] ) );
  AN2 U3567 ( .A(n2378), .B(n2421), .Z(\ab[47][29] ) );
  AN2 U3568 ( .A(n2378), .B(n2419), .Z(\ab[46][29] ) );
  AN2 U3569 ( .A(n2378), .B(n2418), .Z(\ab[45][29] ) );
  AN2 U3570 ( .A(n2378), .B(n2416), .Z(\ab[44][29] ) );
  AN2 U3571 ( .A(n2378), .B(n2415), .Z(\ab[43][29] ) );
  AN2 U3572 ( .A(n2378), .B(n2414), .Z(\ab[42][29] ) );
  AN2 U3573 ( .A(n2378), .B(n316), .Z(\ab[41][29] ) );
  AN2 U3574 ( .A(n2378), .B(n2412), .Z(\ab[40][29] ) );
  AN2 U3575 ( .A(n2378), .B(n2409), .Z(\ab[39][29] ) );
  AN2 U3576 ( .A(n2378), .B(n2405), .Z(\ab[38][29] ) );
  AN2 U3577 ( .A(n2378), .B(n2401), .Z(\ab[37][29] ) );
  AN2 U3578 ( .A(n2379), .B(n254), .Z(\ab[36][29] ) );
  AN2 U3579 ( .A(n2379), .B(n2398), .Z(\ab[35][29] ) );
  AN2 U3580 ( .A(n2379), .B(n2396), .Z(\ab[34][29] ) );
  AN2 U3581 ( .A(n2379), .B(n2393), .Z(\ab[33][29] ) );
  AN2 U3582 ( .A(n2379), .B(n2389), .Z(\ab[32][29] ) );
  AN2 U3583 ( .A(n2379), .B(n2386), .Z(\ab[31][29] ) );
  AN2 U3584 ( .A(n2379), .B(n2383), .Z(\ab[30][29] ) );
  AN2 U3585 ( .A(n2375), .B(\ab[47][47] ), .Z(\ab[47][28] ) );
  AN2 U3586 ( .A(n2375), .B(n2419), .Z(\ab[46][28] ) );
  AN2 U3587 ( .A(n2375), .B(n2418), .Z(\ab[45][28] ) );
  AN2 U3588 ( .A(n2375), .B(n2416), .Z(\ab[44][28] ) );
  AN2 U3589 ( .A(n2375), .B(n2415), .Z(\ab[43][28] ) );
  AN2 U3590 ( .A(n2375), .B(n2414), .Z(\ab[42][28] ) );
  AN2 U3591 ( .A(n2375), .B(n316), .Z(\ab[41][28] ) );
  AN2 U3592 ( .A(n2375), .B(n2412), .Z(\ab[40][28] ) );
  AN2 U3593 ( .A(n2375), .B(n2409), .Z(\ab[39][28] ) );
  AN2 U3594 ( .A(n2375), .B(n2405), .Z(\ab[38][28] ) );
  AN2 U3595 ( .A(n2375), .B(n2401), .Z(\ab[37][28] ) );
  AN2 U3596 ( .A(n2376), .B(n254), .Z(\ab[36][28] ) );
  AN2 U3597 ( .A(n2376), .B(n2398), .Z(\ab[35][28] ) );
  AN2 U3598 ( .A(n2376), .B(n2396), .Z(\ab[34][28] ) );
  AN2 U3599 ( .A(n2376), .B(n2393), .Z(\ab[33][28] ) );
  AN2 U3600 ( .A(n2376), .B(n2389), .Z(\ab[32][28] ) );
  AN2 U3601 ( .A(n2376), .B(n2386), .Z(\ab[31][28] ) );
  AN2 U3602 ( .A(n2376), .B(n2383), .Z(\ab[30][28] ) );
  AN2 U3603 ( .A(n2376), .B(n2379), .Z(\ab[29][28] ) );
  AN2 U3604 ( .A(n2372), .B(n2421), .Z(\ab[47][27] ) );
  AN2 U3605 ( .A(n2372), .B(n2419), .Z(\ab[46][27] ) );
  AN2 U3606 ( .A(n2372), .B(n2418), .Z(\ab[45][27] ) );
  AN2 U3607 ( .A(n2372), .B(n2416), .Z(\ab[44][27] ) );
  AN2 U3608 ( .A(n2372), .B(n2415), .Z(\ab[43][27] ) );
  AN2 U3609 ( .A(n2372), .B(n2414), .Z(\ab[42][27] ) );
  AN2 U3610 ( .A(n2372), .B(n316), .Z(\ab[41][27] ) );
  AN2 U3611 ( .A(n2372), .B(n2412), .Z(\ab[40][27] ) );
  AN2 U3612 ( .A(n2372), .B(n2409), .Z(\ab[39][27] ) );
  AN2 U3613 ( .A(n2372), .B(n2405), .Z(\ab[38][27] ) );
  AN2 U3614 ( .A(n2372), .B(n2401), .Z(\ab[37][27] ) );
  AN2 U3615 ( .A(n2373), .B(n254), .Z(\ab[36][27] ) );
  AN2 U3616 ( .A(n2373), .B(n2398), .Z(\ab[35][27] ) );
  AN2 U3617 ( .A(n2373), .B(n2396), .Z(\ab[34][27] ) );
  AN2 U3618 ( .A(n2373), .B(n2393), .Z(\ab[33][27] ) );
  AN2 U3619 ( .A(n2373), .B(n2389), .Z(\ab[32][27] ) );
  AN2 U3620 ( .A(n2373), .B(n2386), .Z(\ab[31][27] ) );
  AN2 U3621 ( .A(n2373), .B(n2383), .Z(\ab[30][27] ) );
  AN2 U3622 ( .A(n2373), .B(n2379), .Z(\ab[29][27] ) );
  AN2 U3623 ( .A(n2373), .B(n2376), .Z(\ab[28][27] ) );
  AN2 U3624 ( .A(n2370), .B(n2421), .Z(\ab[47][26] ) );
  AN2 U3625 ( .A(n2370), .B(n2419), .Z(\ab[46][26] ) );
  AN2 U3626 ( .A(n2370), .B(n2418), .Z(\ab[45][26] ) );
  AN2 U3627 ( .A(n2370), .B(n2416), .Z(\ab[44][26] ) );
  AN2 U3628 ( .A(n2370), .B(n2415), .Z(\ab[43][26] ) );
  AN2 U3629 ( .A(n2370), .B(n2414), .Z(\ab[42][26] ) );
  AN2 U3630 ( .A(n2370), .B(n316), .Z(\ab[41][26] ) );
  AN2 U3631 ( .A(n2370), .B(n2412), .Z(\ab[40][26] ) );
  AN2 U3632 ( .A(n2370), .B(n2409), .Z(\ab[39][26] ) );
  AN2 U3633 ( .A(n2370), .B(n2405), .Z(\ab[38][26] ) );
  AN2 U3634 ( .A(n2370), .B(n2401), .Z(\ab[37][26] ) );
  AN2 U3635 ( .A(n2370), .B(n254), .Z(\ab[36][26] ) );
  AN2 U3636 ( .A(n2370), .B(n2398), .Z(\ab[35][26] ) );
  AN2 U3637 ( .A(A[26]), .B(n2396), .Z(\ab[34][26] ) );
  AN2 U3638 ( .A(A[26]), .B(n2393), .Z(\ab[33][26] ) );
  AN2 U3639 ( .A(n2370), .B(n2389), .Z(\ab[32][26] ) );
  AN2 U3640 ( .A(A[26]), .B(n2386), .Z(\ab[31][26] ) );
  AN2 U3641 ( .A(n2370), .B(n2383), .Z(\ab[30][26] ) );
  AN2 U3642 ( .A(n2370), .B(n2379), .Z(\ab[29][26] ) );
  AN2 U3643 ( .A(n2370), .B(n2376), .Z(\ab[28][26] ) );
  AN2 U3644 ( .A(n2370), .B(n2373), .Z(\ab[27][26] ) );
  AN2 U3645 ( .A(n2369), .B(\ab[47][47] ), .Z(\ab[47][25] ) );
  AN2 U3646 ( .A(n2369), .B(n2419), .Z(\ab[46][25] ) );
  AN2 U3647 ( .A(n2369), .B(n2418), .Z(\ab[45][25] ) );
  AN2 U3648 ( .A(n2369), .B(n2416), .Z(\ab[44][25] ) );
  AN2 U3649 ( .A(n2369), .B(n2415), .Z(\ab[43][25] ) );
  AN2 U3650 ( .A(n2369), .B(n2414), .Z(\ab[42][25] ) );
  AN2 U3651 ( .A(n2369), .B(n316), .Z(\ab[41][25] ) );
  AN2 U3652 ( .A(n2369), .B(n2412), .Z(\ab[40][25] ) );
  AN2 U3653 ( .A(n2369), .B(n2409), .Z(\ab[39][25] ) );
  AN2 U3654 ( .A(n2369), .B(n2405), .Z(\ab[38][25] ) );
  AN2 U3655 ( .A(n2369), .B(n2401), .Z(\ab[37][25] ) );
  AN2 U3656 ( .A(n247), .B(n254), .Z(\ab[36][25] ) );
  AN2 U3657 ( .A(n247), .B(n2398), .Z(\ab[35][25] ) );
  AN2 U3658 ( .A(n247), .B(n2396), .Z(\ab[34][25] ) );
  AN2 U3659 ( .A(n247), .B(n2393), .Z(\ab[33][25] ) );
  AN2 U3660 ( .A(n247), .B(A[32]), .Z(\ab[32][25] ) );
  AN2 U3661 ( .A(n247), .B(A[31]), .Z(\ab[31][25] ) );
  AN2 U3662 ( .A(n247), .B(n2383), .Z(\ab[30][25] ) );
  AN2 U3663 ( .A(n247), .B(n2379), .Z(\ab[29][25] ) );
  AN2 U3664 ( .A(n247), .B(n2376), .Z(\ab[28][25] ) );
  AN2 U3665 ( .A(n247), .B(n2373), .Z(\ab[27][25] ) );
  AN2 U3666 ( .A(n247), .B(n2370), .Z(\ab[26][25] ) );
  AN2 U3667 ( .A(n2368), .B(n2421), .Z(\ab[47][24] ) );
  AN2 U3668 ( .A(n2368), .B(n2420), .Z(\ab[46][24] ) );
  AN2 U3669 ( .A(n2368), .B(n2418), .Z(\ab[45][24] ) );
  AN2 U3670 ( .A(n2368), .B(n2417), .Z(\ab[44][24] ) );
  AN2 U3671 ( .A(n2368), .B(n2415), .Z(\ab[43][24] ) );
  AN2 U3672 ( .A(n2368), .B(n2414), .Z(\ab[42][24] ) );
  AN2 U3673 ( .A(n2368), .B(n316), .Z(\ab[41][24] ) );
  AN2 U3674 ( .A(n2368), .B(n2412), .Z(\ab[40][24] ) );
  AN2 U3675 ( .A(n2368), .B(n2409), .Z(\ab[39][24] ) );
  AN2 U3676 ( .A(n2368), .B(n2405), .Z(\ab[38][24] ) );
  AN2 U3677 ( .A(n2368), .B(n2401), .Z(\ab[37][24] ) );
  AN2 U3678 ( .A(n267), .B(n254), .Z(\ab[36][24] ) );
  AN2 U3679 ( .A(n267), .B(n2398), .Z(\ab[35][24] ) );
  AN2 U3680 ( .A(n267), .B(n2396), .Z(\ab[34][24] ) );
  AN2 U3681 ( .A(n267), .B(n2393), .Z(\ab[33][24] ) );
  AN2 U3682 ( .A(n267), .B(A[32]), .Z(\ab[32][24] ) );
  AN2 U3683 ( .A(n267), .B(A[31]), .Z(\ab[31][24] ) );
  AN2 U3684 ( .A(n267), .B(n2383), .Z(\ab[30][24] ) );
  AN2 U3685 ( .A(n267), .B(n2379), .Z(\ab[29][24] ) );
  AN2 U3686 ( .A(n267), .B(n2376), .Z(\ab[28][24] ) );
  AN2 U3687 ( .A(n267), .B(n2373), .Z(\ab[27][24] ) );
  AN2 U3688 ( .A(n267), .B(n2370), .Z(\ab[26][24] ) );
  AN2 U3689 ( .A(n267), .B(n247), .Z(\ab[25][24] ) );
  AN2 U3690 ( .A(n2366), .B(n2421), .Z(\ab[47][23] ) );
  AN2 U3691 ( .A(n2366), .B(n2420), .Z(\ab[46][23] ) );
  AN2 U3692 ( .A(n2366), .B(n2418), .Z(\ab[45][23] ) );
  AN2 U3693 ( .A(n2366), .B(n2417), .Z(\ab[44][23] ) );
  AN2 U3694 ( .A(n2366), .B(n737), .Z(\ab[43][23] ) );
  AN2 U3695 ( .A(n2366), .B(n650), .Z(\ab[42][23] ) );
  AN2 U3696 ( .A(n2366), .B(n316), .Z(\ab[41][23] ) );
  AN2 U3697 ( .A(n2366), .B(n652), .Z(\ab[40][23] ) );
  AN2 U3698 ( .A(n2366), .B(n2408), .Z(\ab[39][23] ) );
  AN2 U3699 ( .A(n2366), .B(n2406), .Z(\ab[38][23] ) );
  AN2 U3700 ( .A(n2366), .B(n2402), .Z(\ab[37][23] ) );
  AN2 U3701 ( .A(n2367), .B(n2399), .Z(\ab[36][23] ) );
  AN2 U3702 ( .A(n2367), .B(n300), .Z(\ab[35][23] ) );
  AN2 U3703 ( .A(n2367), .B(n2397), .Z(\ab[34][23] ) );
  AN2 U3704 ( .A(n2367), .B(n2394), .Z(\ab[33][23] ) );
  AN2 U3705 ( .A(n2367), .B(n2390), .Z(\ab[32][23] ) );
  AN2 U3706 ( .A(n2367), .B(n2387), .Z(\ab[31][23] ) );
  AN2 U3707 ( .A(n2367), .B(n2384), .Z(\ab[30][23] ) );
  AN2 U3708 ( .A(n2367), .B(n2380), .Z(\ab[29][23] ) );
  AN2 U3709 ( .A(n2367), .B(n2375), .Z(\ab[28][23] ) );
  AN2 U3710 ( .A(n2367), .B(n2372), .Z(\ab[27][23] ) );
  AN2 U3711 ( .A(n2367), .B(n2370), .Z(\ab[26][23] ) );
  AN2 U3712 ( .A(n2367), .B(n2369), .Z(\ab[25][23] ) );
  AN2 U3713 ( .A(n278), .B(n267), .Z(\ab[24][23] ) );
  AN2 U3714 ( .A(n2364), .B(A[47]), .Z(\ab[47][22] ) );
  AN2 U3715 ( .A(n2364), .B(n2420), .Z(\ab[46][22] ) );
  AN2 U3716 ( .A(n2364), .B(n2418), .Z(\ab[45][22] ) );
  AN2 U3717 ( .A(n2364), .B(n2417), .Z(\ab[44][22] ) );
  AN2 U3718 ( .A(n2364), .B(n2415), .Z(\ab[43][22] ) );
  AN2 U3719 ( .A(n2364), .B(n650), .Z(\ab[42][22] ) );
  AN2 U3720 ( .A(n2364), .B(n316), .Z(\ab[41][22] ) );
  AN2 U3721 ( .A(n2364), .B(n652), .Z(\ab[40][22] ) );
  AN2 U3722 ( .A(n2364), .B(n2408), .Z(\ab[39][22] ) );
  AN2 U3723 ( .A(n2364), .B(n2406), .Z(\ab[38][22] ) );
  AN2 U3724 ( .A(n2364), .B(n2402), .Z(\ab[37][22] ) );
  AN2 U3725 ( .A(n732), .B(n2399), .Z(\ab[36][22] ) );
  AN2 U3726 ( .A(n732), .B(n300), .Z(\ab[35][22] ) );
  AN2 U3727 ( .A(n732), .B(n2397), .Z(\ab[34][22] ) );
  AN2 U3728 ( .A(n732), .B(n2394), .Z(\ab[33][22] ) );
  AN2 U3729 ( .A(n732), .B(n2390), .Z(\ab[32][22] ) );
  AN2 U3730 ( .A(n732), .B(n2387), .Z(\ab[31][22] ) );
  AN2 U3731 ( .A(n732), .B(n2384), .Z(\ab[30][22] ) );
  AN2 U3732 ( .A(n732), .B(n2380), .Z(\ab[29][22] ) );
  AN2 U3733 ( .A(n732), .B(n2375), .Z(\ab[28][22] ) );
  AN2 U3734 ( .A(n732), .B(n2372), .Z(\ab[27][22] ) );
  AN2 U3735 ( .A(n732), .B(n2370), .Z(\ab[26][22] ) );
  AN2 U3736 ( .A(n732), .B(n2369), .Z(\ab[25][22] ) );
  AN2 U3737 ( .A(n2365), .B(n267), .Z(\ab[24][22] ) );
  AN2 U3738 ( .A(n2365), .B(n278), .Z(\ab[23][22] ) );
  AN2 U3739 ( .A(n2362), .B(n2421), .Z(\ab[47][21] ) );
  AN2 U3740 ( .A(n2362), .B(n2420), .Z(\ab[46][21] ) );
  AN2 U3741 ( .A(n2362), .B(n2418), .Z(\ab[45][21] ) );
  AN2 U3742 ( .A(n2362), .B(n2417), .Z(\ab[44][21] ) );
  AN2 U3743 ( .A(n2362), .B(n737), .Z(\ab[43][21] ) );
  AN2 U3744 ( .A(n2362), .B(n650), .Z(\ab[42][21] ) );
  AN2 U3745 ( .A(n2362), .B(n316), .Z(\ab[41][21] ) );
  AN2 U3746 ( .A(n2362), .B(n652), .Z(\ab[40][21] ) );
  AN2 U3747 ( .A(n2362), .B(n2408), .Z(\ab[39][21] ) );
  AN2 U3748 ( .A(n2362), .B(n2406), .Z(\ab[38][21] ) );
  AN2 U3749 ( .A(n2362), .B(n2402), .Z(\ab[37][21] ) );
  AN2 U3750 ( .A(n730), .B(n2399), .Z(\ab[36][21] ) );
  AN2 U3751 ( .A(n730), .B(n300), .Z(\ab[35][21] ) );
  AN2 U3752 ( .A(n730), .B(n2397), .Z(\ab[34][21] ) );
  AN2 U3753 ( .A(n730), .B(n2394), .Z(\ab[33][21] ) );
  AN2 U3754 ( .A(n730), .B(n2390), .Z(\ab[32][21] ) );
  AN2 U3755 ( .A(n730), .B(n2387), .Z(\ab[31][21] ) );
  AN2 U3756 ( .A(n730), .B(n2384), .Z(\ab[30][21] ) );
  AN2 U3757 ( .A(n730), .B(n2380), .Z(\ab[29][21] ) );
  AN2 U3758 ( .A(n730), .B(n2375), .Z(\ab[28][21] ) );
  AN2 U3759 ( .A(n730), .B(n2372), .Z(\ab[27][21] ) );
  AN2 U3760 ( .A(n730), .B(n2370), .Z(\ab[26][21] ) );
  AN2 U3761 ( .A(n730), .B(n2369), .Z(\ab[25][21] ) );
  AN2 U3762 ( .A(n2363), .B(n267), .Z(\ab[24][21] ) );
  AN2 U3763 ( .A(n2363), .B(n278), .Z(\ab[23][21] ) );
  AN2 U3764 ( .A(n2363), .B(n2365), .Z(\ab[22][21] ) );
  AN2 U3765 ( .A(n2360), .B(n2421), .Z(\ab[47][20] ) );
  AN2 U3766 ( .A(n2360), .B(n2420), .Z(\ab[46][20] ) );
  AN2 U3767 ( .A(n2360), .B(n2418), .Z(\ab[45][20] ) );
  AN2 U3768 ( .A(n2360), .B(n2417), .Z(\ab[44][20] ) );
  AN2 U3769 ( .A(n2360), .B(n737), .Z(\ab[43][20] ) );
  AN2 U3770 ( .A(n2360), .B(n650), .Z(\ab[42][20] ) );
  AN2 U3771 ( .A(n2360), .B(n316), .Z(\ab[41][20] ) );
  AN2 U3772 ( .A(n2360), .B(n652), .Z(\ab[40][20] ) );
  AN2 U3773 ( .A(n2360), .B(n2408), .Z(\ab[39][20] ) );
  AN2 U3774 ( .A(n2360), .B(n2406), .Z(\ab[38][20] ) );
  AN2 U3775 ( .A(n2360), .B(n2402), .Z(\ab[37][20] ) );
  AN2 U3776 ( .A(n2361), .B(n2399), .Z(\ab[36][20] ) );
  AN2 U3777 ( .A(n2361), .B(n300), .Z(\ab[35][20] ) );
  AN2 U3778 ( .A(n2361), .B(n2397), .Z(\ab[34][20] ) );
  AN2 U3779 ( .A(n2361), .B(n2394), .Z(\ab[33][20] ) );
  AN2 U3780 ( .A(n2361), .B(n2390), .Z(\ab[32][20] ) );
  AN2 U3781 ( .A(n2361), .B(n2387), .Z(\ab[31][20] ) );
  AN2 U3782 ( .A(n2361), .B(n2384), .Z(\ab[30][20] ) );
  AN2 U3783 ( .A(n2361), .B(n2380), .Z(\ab[29][20] ) );
  AN2 U3784 ( .A(n2361), .B(n2375), .Z(\ab[28][20] ) );
  AN2 U3785 ( .A(n2361), .B(n2372), .Z(\ab[27][20] ) );
  AN2 U3786 ( .A(n2361), .B(n2370), .Z(\ab[26][20] ) );
  AN2 U3787 ( .A(n2361), .B(n2369), .Z(\ab[25][20] ) );
  AN2 U3788 ( .A(n245), .B(n267), .Z(\ab[24][20] ) );
  AN2 U3789 ( .A(n245), .B(n278), .Z(\ab[23][20] ) );
  AN2 U3790 ( .A(n245), .B(n2365), .Z(\ab[22][20] ) );
  AN2 U3791 ( .A(n245), .B(n2363), .Z(\ab[21][20] ) );
  AN2 U3792 ( .A(n2358), .B(A[47]), .Z(\ab[47][19] ) );
  AN2 U3793 ( .A(n2358), .B(n2420), .Z(\ab[46][19] ) );
  AN2 U3794 ( .A(n2358), .B(n2418), .Z(\ab[45][19] ) );
  AN2 U3795 ( .A(n2358), .B(n2417), .Z(\ab[44][19] ) );
  AN2 U3796 ( .A(n2358), .B(n2415), .Z(\ab[43][19] ) );
  AN2 U3797 ( .A(n2358), .B(n650), .Z(\ab[42][19] ) );
  AN2 U3798 ( .A(n2358), .B(n316), .Z(\ab[41][19] ) );
  AN2 U3799 ( .A(n2358), .B(n652), .Z(\ab[40][19] ) );
  AN2 U3800 ( .A(n2358), .B(n2408), .Z(\ab[39][19] ) );
  AN2 U3801 ( .A(n2358), .B(n2406), .Z(\ab[38][19] ) );
  AN2 U3802 ( .A(n2358), .B(n2402), .Z(\ab[37][19] ) );
  AN2 U3803 ( .A(n2359), .B(n2399), .Z(\ab[36][19] ) );
  AN2 U3804 ( .A(n2359), .B(n300), .Z(\ab[35][19] ) );
  AN2 U3805 ( .A(n2359), .B(n2397), .Z(\ab[34][19] ) );
  AN2 U3806 ( .A(n2359), .B(n2394), .Z(\ab[33][19] ) );
  AN2 U3807 ( .A(n2359), .B(n2390), .Z(\ab[32][19] ) );
  AN2 U3808 ( .A(n2359), .B(n2387), .Z(\ab[31][19] ) );
  AN2 U3809 ( .A(n2359), .B(n2384), .Z(\ab[30][19] ) );
  AN2 U3810 ( .A(n2359), .B(n2380), .Z(\ab[29][19] ) );
  AN2 U3811 ( .A(n2359), .B(n2375), .Z(\ab[28][19] ) );
  AN2 U3812 ( .A(n2359), .B(n2372), .Z(\ab[27][19] ) );
  AN2 U3813 ( .A(n2359), .B(n2370), .Z(\ab[26][19] ) );
  AN2 U3814 ( .A(n2359), .B(n2369), .Z(\ab[25][19] ) );
  AN2 U3815 ( .A(n250), .B(n267), .Z(\ab[24][19] ) );
  AN2 U3816 ( .A(n250), .B(n278), .Z(\ab[23][19] ) );
  AN2 U3817 ( .A(n250), .B(n2365), .Z(\ab[22][19] ) );
  AN2 U3818 ( .A(n250), .B(n2363), .Z(\ab[21][19] ) );
  AN2 U3819 ( .A(n250), .B(n245), .Z(\ab[20][19] ) );
  AN2 U3820 ( .A(n2356), .B(n2421), .Z(\ab[47][18] ) );
  AN2 U3821 ( .A(n2356), .B(n2420), .Z(\ab[46][18] ) );
  AN2 U3822 ( .A(n2356), .B(n2418), .Z(\ab[45][18] ) );
  AN2 U3823 ( .A(n2356), .B(n2417), .Z(\ab[44][18] ) );
  AN2 U3824 ( .A(n2356), .B(n737), .Z(\ab[43][18] ) );
  AN2 U3825 ( .A(n2356), .B(n650), .Z(\ab[42][18] ) );
  AN2 U3826 ( .A(n2356), .B(n316), .Z(\ab[41][18] ) );
  AN2 U3827 ( .A(n2356), .B(n652), .Z(\ab[40][18] ) );
  AN2 U3828 ( .A(n2356), .B(n2408), .Z(\ab[39][18] ) );
  AN2 U3829 ( .A(n2356), .B(n2406), .Z(\ab[38][18] ) );
  AN2 U3830 ( .A(n2356), .B(n2402), .Z(\ab[37][18] ) );
  AN2 U3831 ( .A(n2357), .B(n2399), .Z(\ab[36][18] ) );
  AN2 U3832 ( .A(n2357), .B(n300), .Z(\ab[35][18] ) );
  AN2 U3833 ( .A(n2357), .B(n2397), .Z(\ab[34][18] ) );
  AN2 U3834 ( .A(n2357), .B(n2394), .Z(\ab[33][18] ) );
  AN2 U3835 ( .A(n2357), .B(n2390), .Z(\ab[32][18] ) );
  AN2 U3836 ( .A(n2357), .B(n2387), .Z(\ab[31][18] ) );
  AN2 U3837 ( .A(n2357), .B(n2384), .Z(\ab[30][18] ) );
  AN2 U3838 ( .A(n2357), .B(n2380), .Z(\ab[29][18] ) );
  AN2 U3839 ( .A(n2357), .B(n2375), .Z(\ab[28][18] ) );
  AN2 U3840 ( .A(n2357), .B(n2372), .Z(\ab[27][18] ) );
  AN2 U3841 ( .A(n2357), .B(n2370), .Z(\ab[26][18] ) );
  AN2 U3842 ( .A(n2357), .B(n2369), .Z(\ab[25][18] ) );
  AN2 U3843 ( .A(n259), .B(n267), .Z(\ab[24][18] ) );
  AN2 U3844 ( .A(n259), .B(n278), .Z(\ab[23][18] ) );
  AN2 U3845 ( .A(n259), .B(n2365), .Z(\ab[22][18] ) );
  AN2 U3846 ( .A(n259), .B(n2363), .Z(\ab[21][18] ) );
  AN2 U3847 ( .A(n259), .B(n245), .Z(\ab[20][18] ) );
  AN2 U3848 ( .A(n259), .B(n250), .Z(\ab[19][18] ) );
  AN2 U3849 ( .A(n2355), .B(n2421), .Z(\ab[47][17] ) );
  AN2 U3850 ( .A(n2355), .B(n2420), .Z(\ab[46][17] ) );
  AN2 U3851 ( .A(n2355), .B(n2418), .Z(\ab[45][17] ) );
  AN2 U3852 ( .A(n2355), .B(n2417), .Z(\ab[44][17] ) );
  AN2 U3853 ( .A(n2355), .B(n737), .Z(\ab[43][17] ) );
  AN2 U3854 ( .A(n2355), .B(n650), .Z(\ab[42][17] ) );
  AN2 U3855 ( .A(n2355), .B(n316), .Z(\ab[41][17] ) );
  AN2 U3856 ( .A(n2355), .B(n652), .Z(\ab[40][17] ) );
  AN2 U3857 ( .A(n2355), .B(n2408), .Z(\ab[39][17] ) );
  AN2 U3858 ( .A(n2355), .B(n2406), .Z(\ab[38][17] ) );
  AN2 U3859 ( .A(n2355), .B(n2402), .Z(\ab[37][17] ) );
  AN2 U3860 ( .A(n728), .B(n2399), .Z(\ab[36][17] ) );
  AN2 U3861 ( .A(n728), .B(n300), .Z(\ab[35][17] ) );
  AN2 U3862 ( .A(n728), .B(n2397), .Z(\ab[34][17] ) );
  AN2 U3863 ( .A(n728), .B(n2394), .Z(\ab[33][17] ) );
  AN2 U3864 ( .A(n728), .B(n2390), .Z(\ab[32][17] ) );
  AN2 U3865 ( .A(n728), .B(n2387), .Z(\ab[31][17] ) );
  AN2 U3866 ( .A(n728), .B(n2384), .Z(\ab[30][17] ) );
  AN2 U3867 ( .A(n728), .B(n2380), .Z(\ab[29][17] ) );
  AN2 U3868 ( .A(n728), .B(n2375), .Z(\ab[28][17] ) );
  AN2 U3869 ( .A(n728), .B(n2372), .Z(\ab[27][17] ) );
  AN2 U3870 ( .A(n728), .B(n2370), .Z(\ab[26][17] ) );
  AN2 U3871 ( .A(n728), .B(n2369), .Z(\ab[25][17] ) );
  AN2 U3872 ( .A(n2355), .B(n267), .Z(\ab[24][17] ) );
  AN2 U3873 ( .A(n2355), .B(n278), .Z(\ab[23][17] ) );
  AN2 U3874 ( .A(n2355), .B(n2365), .Z(\ab[22][17] ) );
  AN2 U3875 ( .A(n2355), .B(n2363), .Z(\ab[21][17] ) );
  AN2 U3876 ( .A(n728), .B(n245), .Z(\ab[20][17] ) );
  AN2 U3877 ( .A(n2355), .B(n250), .Z(\ab[19][17] ) );
  AN2 U3878 ( .A(n2355), .B(n259), .Z(\ab[18][17] ) );
  AN2 U3879 ( .A(n2352), .B(A[47]), .Z(\ab[47][16] ) );
  AN2 U3880 ( .A(n2352), .B(n2420), .Z(\ab[46][16] ) );
  AN2 U3881 ( .A(n2352), .B(n2418), .Z(\ab[45][16] ) );
  AN2 U3882 ( .A(n2352), .B(n2417), .Z(\ab[44][16] ) );
  AN2 U3883 ( .A(n2352), .B(n2415), .Z(\ab[43][16] ) );
  AN2 U3884 ( .A(n2352), .B(n650), .Z(\ab[42][16] ) );
  AN2 U3885 ( .A(n2352), .B(n316), .Z(\ab[41][16] ) );
  AN2 U3886 ( .A(n2352), .B(n652), .Z(\ab[40][16] ) );
  AN2 U3887 ( .A(n2352), .B(n2408), .Z(\ab[39][16] ) );
  AN2 U3888 ( .A(n2352), .B(n2406), .Z(\ab[38][16] ) );
  AN2 U3889 ( .A(n2352), .B(n2402), .Z(\ab[37][16] ) );
  AN2 U3890 ( .A(n2353), .B(n2399), .Z(\ab[36][16] ) );
  AN2 U3891 ( .A(n2353), .B(n300), .Z(\ab[35][16] ) );
  AN2 U3892 ( .A(n2353), .B(n2397), .Z(\ab[34][16] ) );
  AN2 U3893 ( .A(n2353), .B(n2394), .Z(\ab[33][16] ) );
  AN2 U3894 ( .A(n2353), .B(n2390), .Z(\ab[32][16] ) );
  AN2 U3895 ( .A(n2353), .B(n2387), .Z(\ab[31][16] ) );
  AN2 U3896 ( .A(n2353), .B(n2384), .Z(\ab[30][16] ) );
  AN2 U3897 ( .A(n2353), .B(n2380), .Z(\ab[29][16] ) );
  AN2 U3898 ( .A(n2353), .B(n2375), .Z(\ab[28][16] ) );
  AN2 U3899 ( .A(n2353), .B(n2372), .Z(\ab[27][16] ) );
  AN2 U3900 ( .A(n2353), .B(n2370), .Z(\ab[26][16] ) );
  AN2 U3901 ( .A(n2353), .B(n2369), .Z(\ab[25][16] ) );
  AN2 U3902 ( .A(n2352), .B(n267), .Z(\ab[24][16] ) );
  AN2 U3903 ( .A(n2352), .B(n278), .Z(\ab[23][16] ) );
  AN2 U3904 ( .A(n2352), .B(n2365), .Z(\ab[22][16] ) );
  AN2 U3905 ( .A(n2352), .B(n2363), .Z(\ab[21][16] ) );
  AN2 U3906 ( .A(n2352), .B(n245), .Z(\ab[20][16] ) );
  AN2 U3907 ( .A(n2352), .B(n250), .Z(\ab[19][16] ) );
  AN2 U3908 ( .A(n2352), .B(n259), .Z(\ab[18][16] ) );
  AN2 U3909 ( .A(n2352), .B(n2355), .Z(\ab[17][16] ) );
  AN2 U3910 ( .A(n2349), .B(n2421), .Z(\ab[47][15] ) );
  AN2 U3911 ( .A(n2349), .B(n2420), .Z(\ab[46][15] ) );
  AN2 U3912 ( .A(n2349), .B(n2418), .Z(\ab[45][15] ) );
  AN2 U3913 ( .A(n2349), .B(n2417), .Z(\ab[44][15] ) );
  AN2 U3914 ( .A(n2349), .B(n737), .Z(\ab[43][15] ) );
  AN2 U3915 ( .A(n2349), .B(n650), .Z(\ab[42][15] ) );
  AN2 U3916 ( .A(n2349), .B(n316), .Z(\ab[41][15] ) );
  AN2 U3917 ( .A(n2349), .B(n652), .Z(\ab[40][15] ) );
  AN2 U3918 ( .A(n2349), .B(n2408), .Z(\ab[39][15] ) );
  AN2 U3919 ( .A(n2349), .B(n2406), .Z(\ab[38][15] ) );
  AN2 U3920 ( .A(n2349), .B(n2402), .Z(\ab[37][15] ) );
  AN2 U3921 ( .A(n2350), .B(n2399), .Z(\ab[36][15] ) );
  AN2 U3922 ( .A(n2350), .B(n300), .Z(\ab[35][15] ) );
  AN2 U3923 ( .A(n2350), .B(n2397), .Z(\ab[34][15] ) );
  AN2 U3924 ( .A(n2350), .B(n2394), .Z(\ab[33][15] ) );
  AN2 U3925 ( .A(n2350), .B(n2390), .Z(\ab[32][15] ) );
  AN2 U3926 ( .A(n2350), .B(n2387), .Z(\ab[31][15] ) );
  AN2 U3927 ( .A(n2350), .B(n2384), .Z(\ab[30][15] ) );
  AN2 U3928 ( .A(n261), .B(n2421), .Z(\ab[47][14] ) );
  AN2 U3929 ( .A(n261), .B(n2420), .Z(\ab[46][14] ) );
  AN2 U3930 ( .A(n261), .B(A[45]), .Z(\ab[45][14] ) );
  AN2 U3931 ( .A(n261), .B(n2417), .Z(\ab[44][14] ) );
  AN2 U3932 ( .A(n261), .B(n2415), .Z(\ab[43][14] ) );
  AN2 U3933 ( .A(n261), .B(n650), .Z(\ab[42][14] ) );
  AN2 U3934 ( .A(n261), .B(n316), .Z(\ab[41][14] ) );
  AN2 U3935 ( .A(n261), .B(n652), .Z(\ab[40][14] ) );
  AN2 U3936 ( .A(n261), .B(n2409), .Z(\ab[39][14] ) );
  AN2 U3937 ( .A(n261), .B(n2406), .Z(\ab[38][14] ) );
  AN2 U3938 ( .A(n261), .B(n2402), .Z(\ab[37][14] ) );
  AN2 U3939 ( .A(n2347), .B(n254), .Z(\ab[36][14] ) );
  AN2 U3940 ( .A(n2347), .B(n300), .Z(\ab[35][14] ) );
  AN2 U3941 ( .A(n2347), .B(n2397), .Z(\ab[34][14] ) );
  AN2 U3942 ( .A(n2347), .B(n2394), .Z(\ab[33][14] ) );
  AN2 U3943 ( .A(n2347), .B(n2390), .Z(\ab[32][14] ) );
  AN2 U3944 ( .A(n2347), .B(n2387), .Z(\ab[31][14] ) );
  AN2 U3945 ( .A(n2346), .B(A[47]), .Z(\ab[47][13] ) );
  AN2 U3946 ( .A(n2346), .B(n2420), .Z(\ab[46][13] ) );
  AN2 U3947 ( .A(n2346), .B(A[45]), .Z(\ab[45][13] ) );
  AN2 U3948 ( .A(n2346), .B(n2417), .Z(\ab[44][13] ) );
  AN2 U3949 ( .A(n2346), .B(n737), .Z(\ab[43][13] ) );
  AN2 U3950 ( .A(n2346), .B(n650), .Z(\ab[42][13] ) );
  AN2 U3951 ( .A(n2346), .B(A[41]), .Z(\ab[41][13] ) );
  AN2 U3952 ( .A(n2346), .B(n652), .Z(\ab[40][13] ) );
  AN2 U3953 ( .A(n2346), .B(A[39]), .Z(\ab[39][13] ) );
  AN2 U3954 ( .A(n2346), .B(n2406), .Z(\ab[38][13] ) );
  AN2 U3955 ( .A(n2346), .B(n2402), .Z(\ab[37][13] ) );
  AN2 U3956 ( .A(n2346), .B(A[36]), .Z(\ab[36][13] ) );
  AN2 U3957 ( .A(n2346), .B(n300), .Z(\ab[35][13] ) );
  AN2 U3958 ( .A(n2346), .B(n2397), .Z(\ab[34][13] ) );
  AN2 U3959 ( .A(n2346), .B(n2394), .Z(\ab[33][13] ) );
  AN2 U3960 ( .A(n265), .B(n2421), .Z(\ab[47][12] ) );
  AN2 U3961 ( .A(n265), .B(n2419), .Z(\ab[46][12] ) );
  AN2 U3962 ( .A(n265), .B(n2418), .Z(\ab[45][12] ) );
  AN2 U3963 ( .A(n265), .B(n280), .Z(\ab[44][12] ) );
  AN2 U3964 ( .A(n265), .B(A[43]), .Z(\ab[43][12] ) );
  AN2 U3965 ( .A(n265), .B(n650), .Z(\ab[42][12] ) );
  AN2 U3966 ( .A(n265), .B(A[41]), .Z(\ab[41][12] ) );
  AN2 U3967 ( .A(n265), .B(n652), .Z(\ab[40][12] ) );
  AN2 U3968 ( .A(n265), .B(A[39]), .Z(\ab[39][12] ) );
  AN2 U3969 ( .A(n265), .B(n2406), .Z(\ab[38][12] ) );
  AN2 U3970 ( .A(n265), .B(n2402), .Z(\ab[37][12] ) );
  AN2 U3971 ( .A(n265), .B(A[36]), .Z(\ab[36][12] ) );
  AN2 U3972 ( .A(n2341), .B(n2421), .Z(\ab[47][11] ) );
  AN2 U3973 ( .A(n2341), .B(n2419), .Z(\ab[46][11] ) );
  AN2 U3974 ( .A(n2341), .B(n2418), .Z(\ab[45][11] ) );
  AN2 U3975 ( .A(n2341), .B(n280), .Z(\ab[44][11] ) );
  AN2 U3976 ( .A(n2341), .B(n2415), .Z(\ab[43][11] ) );
  AN2 U3977 ( .A(n2341), .B(n2413), .Z(\ab[42][11] ) );
  AN2 U3978 ( .A(n2341), .B(n316), .Z(\ab[41][11] ) );
  AN2 U3979 ( .A(n2341), .B(n2411), .Z(\ab[40][11] ) );
  AN2 U3980 ( .A(n2341), .B(n2409), .Z(\ab[39][11] ) );
  AN2 U3981 ( .A(n2341), .B(n2404), .Z(\ab[38][11] ) );
  AN2 U3982 ( .A(n2339), .B(A[47]), .Z(\ab[47][10] ) );
  AN2 U3983 ( .A(n2339), .B(n2419), .Z(\ab[46][10] ) );
  AN2 U3984 ( .A(n2339), .B(n2418), .Z(\ab[45][10] ) );
  AN2 U3985 ( .A(n2339), .B(n280), .Z(\ab[44][10] ) );
  AN2 U3986 ( .A(n2339), .B(n2415), .Z(\ab[43][10] ) );
  AN2 U3987 ( .A(n2339), .B(n2413), .Z(\ab[42][10] ) );
  AN2 U3988 ( .A(n2339), .B(n316), .Z(\ab[41][10] ) );
endmodule


module LOG_POLY ( clk, reset, LogIn, LogOut );
  input [47:0] LogIn;
  output [30:0] LogOut;
  input clk, reset;
  wire   N9, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N254, N255, N256, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, N277, N292, N293,
         N294, N295, N296, N297, N298, N284, N283, N282, N281, N280, N279,
         N278, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243,
         N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232,
         N231, N230, \add_1_root_sub_1_root_add_225_2/carry[6] ,
         \add_1_root_sub_1_root_add_225_2/carry[5] ,
         \add_1_root_sub_1_root_add_225_2/carry[4] ,
         \add_1_root_sub_1_root_add_225_2/carry[3] ,
         \add_1_root_sub_1_root_add_225_2/carry[2] ,
         \add_1_root_sub_1_root_add_225_2/carry[1] , n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071;
  wire   [95:0] LogInSquare;
  wire   [47:0] LogIn2;
  wire   [118:89] Term1;
  wire   [67:38] Term2;
  wire   [26:1] Term3;
  wire   [118:112] Term11;
  wire   [67:61] Term21;
  wire   [26:24] Term31;
  wire   [23:0] FractionBit;
  wire   [6:0] IntegerBits;
  wire   [22:0] LogPipe;
  wire   [29:0] Log;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136;
  assign LogOut[0] = 1'b0;

  LOG_POLY_DW02_mult_2 mult_214 ( .A({n29, n28, n27, n70, n64, n63, N171, N172, 
        N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, 
        N185, N186}), .B(LogIn2), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, N216, N215, N214, N213, N212, N211, N210, 
        N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, 
        N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39}) );
  LOG_POLY_DW02_mult_1 mult_213 ( .A({n34, n33, n32, n31, n30, n81, n80, n444, 
        n72, n69, n67, N116, N117, N118, N119, N120, N121, N122, N123, N124, 
        N125, N126, N127, N128, N129, N130, N131, N132, N133, N134}), .B(
        LogInSquare), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N164, N163, N162, 
        N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, 
        N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137, N136, N135, SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135}) );
  LOG_POLY_DW01_sub_0 sub_0_root_sub_1_root_add_225_2 ( .A({N284, N283, N282, 
        N281, N280, N279, N278}), .B(Term21), .CI(1'b0), .DIFF({N298, N297, 
        N296, N295, N294, N293, N292}) );
  LOG_POLY_DW01_sub_1 sub_0_root_sub_0_root_add_222 ( .A({n445, N252, N251, 
        N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, 
        N238, N237, N236, N235, N234, N233, N232, N231, N230}), .B({1'b0, 
        Term2[60:38]}), .CI(1'b0), .DIFF({N277, N276, N275, N274, N273, N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254}) );
  LOG_POLY_DW02_mult_0 mult_209 ( .A({LogIn[47:8], n22, LogIn[6:2], n405, n35}), .B({LogIn[47:8], n22, LogIn[6:0]}), .TC(1'b0), .PRODUCT({N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, SYNOPSYS_UNCONNECTED__136, N9}) );
  FDS2L \LogIn2_reg[0]  ( .CR(1'b1), .D(n35), .LD(n5040), .CP(clk), .Q(
        LogIn2[0]) );
  FDS2L \LogIn2_reg[1]  ( .CR(1'b1), .D(n405), .LD(n5041), .CP(clk), .Q(
        LogIn2[1]) );
  FDS2L \LogIn2_reg[12]  ( .CR(1'b1), .D(LogIn[12]), .LD(n5041), .CP(clk), .Q(
        LogIn2[12]) );
  FDS2L \LogInSquare_reg[33]  ( .CR(1'b1), .D(N42), .LD(n5027), .CP(clk), .Q(
        LogInSquare[33]) );
  FD1 \LogInSquare_reg[68]  ( .D(n36), .CP(clk), .Q(LogInSquare[68]) );
  FD1 \LogInSquare_reg[73]  ( .D(n489), .CP(clk), .Q(LogInSquare[73]) );
  FD1 \LogInSquare_reg[77]  ( .D(n487), .CP(clk), .Q(LogInSquare[77]) );
  FD1 \LogInSquare_reg[80]  ( .D(n485), .CP(clk), .Q(LogInSquare[80]) );
  MUX21L \LogInSquare_reg[88]/U5  ( .A(LogInSquare[88]), .B(N97), .S(n5048), 
        .Z(n482) );
  FD1 \LogInSquare_reg[88]  ( .D(n483), .CP(clk), .Q(LogInSquare[88]) );
  MUX21L \LogInSquare_reg[87]/U5  ( .A(LogInSquare[87]), .B(N96), .S(n5048), 
        .Z(n480) );
  FD1 \LogInSquare_reg[87]  ( .D(n481), .CP(clk), .Q(LogInSquare[87]) );
  MUX21L \LogInSquare_reg[86]/U5  ( .A(LogInSquare[86]), .B(N95), .S(n5048), 
        .Z(n478) );
  FD1 \LogInSquare_reg[86]  ( .D(n479), .CP(clk), .Q(LogInSquare[86]) );
  MUX21L \LogInSquare_reg[83]/U5  ( .A(LogInSquare[83]), .B(N92), .S(n5047), 
        .Z(n476) );
  FD1 \LogInSquare_reg[83]  ( .D(n477), .CP(clk), .Q(LogInSquare[83]) );
  MUX21L \LogInSquare_reg[64]/U5  ( .A(LogInSquare[64]), .B(N73), .S(n5046), 
        .Z(n474) );
  FD1 \LogInSquare_reg[64]  ( .D(n475), .CP(clk), .Q(LogInSquare[64]) );
  FD1 \LogInSquare_reg[81]  ( .D(n473), .CP(clk), .Q(LogInSquare[81]) );
  MUX21L \LogInSquare_reg[85]/U5  ( .A(LogInSquare[85]), .B(N94), .S(n5048), 
        .Z(n470) );
  FD1 \LogInSquare_reg[85]  ( .D(n471), .CP(clk), .Q(LogInSquare[85]) );
  MUX21L \LogInSquare_reg[84]/U5  ( .A(LogInSquare[84]), .B(N93), .S(n5048), 
        .Z(n468) );
  FD1 \LogInSquare_reg[84]  ( .D(n469), .CP(clk), .Q(LogInSquare[84]) );
  FD1 \LogInSquare_reg[69]  ( .D(n467), .CP(clk), .Q(LogInSquare[69]) );
  MUX21L \LogInSquare_reg[89]/U5  ( .A(LogInSquare[89]), .B(N98), .S(n5048), 
        .Z(n464) );
  FD1 \LogInSquare_reg[89]  ( .D(n465), .CP(clk), .Q(LogInSquare[89]) );
  FD1 \LogInSquare_reg[95]  ( .D(n463), .CP(clk), .Q(LogInSquare[95]) );
  FD1 \LogInSquare_reg[65]  ( .D(n461), .CP(clk), .Q(LogInSquare[65]) );
  FD1 \LogInSquare_reg[94]  ( .D(n459), .CP(clk), .Q(LogInSquare[94]) );
  FD1 \LogInSquare_reg[93]  ( .D(n457), .CP(clk), .Q(LogInSquare[93]) );
  FD1 \LogInSquare_reg[92]  ( .D(n455), .CP(clk), .Q(LogInSquare[92]) );
  FD1 \LogInSquare_reg[91]  ( .D(n453), .CP(clk), .Q(LogInSquare[91]) );
  FD1 \LogInSquare_reg[90]  ( .D(n451), .CP(clk), .Q(LogInSquare[90]) );
  FD1 \LogInSquare_reg[61]  ( .D(n449), .CP(clk), .Q(LogInSquare[61]) );
  FDS2L \LogInSquare_reg[72]  ( .CR(1'b1), .D(N81), .LD(n5047), .CP(clk), .Q(
        LogInSquare[72]) );
  FDS2L \Term2_reg[60]  ( .CR(1'b1), .D(N209), .LD(n5037), .CP(clk), .Q(
        Term2[60]) );
  FDS2L \Term2_reg[59]  ( .CR(1'b1), .D(N208), .LD(n5037), .CP(clk), .Q(
        Term2[59]) );
  FDS2L \Term1_reg[111]  ( .CR(1'b1), .D(N157), .LD(n5040), .CP(clk), .Q(
        Term1[111]), .QN(n446) );
  FDS2L \Term3_reg[23]  ( .CR(1'b1), .D(N220), .LD(n5030), .CP(clk), .Q(
        Term3[23]), .QN(n447) );
  FDS2L \Term2_reg[58]  ( .CR(1'b1), .D(N207), .LD(n5037), .CP(clk), .Q(
        Term2[58]) );
  FDS2L \Term1_reg[110]  ( .CR(1'b1), .D(N156), .LD(n5040), .CP(clk), .Q(
        Term1[110]) );
  FDS2L \Term2_reg[57]  ( .CR(1'b1), .D(N206), .LD(n5037), .CP(clk), .Q(
        Term2[57]) );
  FDS2L \Term3_reg[22]  ( .CR(1'b1), .D(N221), .LD(n5030), .CP(clk), .Q(
        Term3[22]) );
  FDS2L \Term2_reg[56]  ( .CR(1'b1), .D(N205), .LD(n5037), .CP(clk), .Q(
        Term2[56]) );
  FDS2L \Term1_reg[109]  ( .CR(1'b1), .D(N155), .LD(n5040), .CP(clk), .Q(
        Term1[109]) );
  FDS2L \Term2_reg[55]  ( .CR(1'b1), .D(N204), .LD(n5037), .CP(clk), .Q(
        Term2[55]) );
  FDS2L \Term3_reg[21]  ( .CR(1'b1), .D(N222), .LD(n5030), .CP(clk), .Q(
        Term3[21]) );
  FDS2L \FractionBit_reg[23]  ( .CR(1'b1), .D(N277), .LD(n5034), .CP(clk), .Q(
        FractionBit[23]) );
  FDS2L \Term2_reg[54]  ( .CR(1'b1), .D(N203), .LD(n5037), .CP(clk), .Q(
        Term2[54]) );
  FDS2L \Term1_reg[108]  ( .CR(1'b1), .D(N154), .LD(n5040), .CP(clk), .Q(
        Term1[108]) );
  FDS2L \Term2_reg[53]  ( .CR(1'b1), .D(N202), .LD(n5037), .CP(clk), .Q(
        Term2[53]) );
  FDS2L \Term3_reg[20]  ( .CR(1'b1), .D(N223), .LD(n5029), .CP(clk), .Q(
        Term3[20]) );
  FDS2L \Term2_reg[52]  ( .CR(1'b1), .D(N201), .LD(n5037), .CP(clk), .Q(
        Term2[52]) );
  FDS2L \Term1_reg[107]  ( .CR(1'b1), .D(N153), .LD(n5039), .CP(clk), .Q(
        Term1[107]) );
  FDS2L \Term2_reg[51]  ( .CR(1'b1), .D(N200), .LD(n5037), .CP(clk), .Q(
        Term2[51]) );
  FDS2L \Term3_reg[19]  ( .CR(1'b1), .D(N224), .LD(n5029), .CP(clk), .Q(
        Term3[19]) );
  FDS2L \Term1_reg[101]  ( .CR(1'b1), .D(N147), .LD(n5039), .CP(clk), .Q(N242)
         );
  FDS2L \Term1_reg[100]  ( .CR(1'b1), .D(N146), .LD(n5039), .CP(clk), .Q(N241)
         );
  FDS2L \Term1_reg[106]  ( .CR(1'b1), .D(N152), .LD(n5039), .CP(clk), .Q(
        Term1[106]) );
  FDS2L \Term2_reg[50]  ( .CR(1'b1), .D(N199), .LD(n5036), .CP(clk), .Q(
        Term2[50]) );
  FDS2L \Term3_reg[18]  ( .CR(1'b1), .D(N225), .LD(n5029), .CP(clk), .Q(
        Term3[18]) );
  FDS2L \Term2_reg[49]  ( .CR(1'b1), .D(N198), .LD(n5036), .CP(clk), .Q(
        Term2[49]) );
  FDS2L \Term1_reg[99]  ( .CR(1'b1), .D(N145), .LD(n5039), .CP(clk), .Q(N240)
         );
  FDS2L \Term2_reg[48]  ( .CR(1'b1), .D(N197), .LD(n5036), .CP(clk), .Q(
        Term2[48]) );
  FDS2L \Term1_reg[98]  ( .CR(1'b1), .D(N144), .LD(n5039), .CP(clk), .Q(N239)
         );
  FDS2L \Term1_reg[105]  ( .CR(1'b1), .D(N151), .LD(n5039), .CP(clk), .Q(
        Term1[105]) );
  FDS2L \Term2_reg[47]  ( .CR(1'b1), .D(N196), .LD(n5036), .CP(clk), .Q(
        Term2[47]) );
  FDS2L \Term3_reg[17]  ( .CR(1'b1), .D(N226), .LD(n5029), .CP(clk), .Q(
        Term3[17]) );
  FDS2L \Term1_reg[97]  ( .CR(1'b1), .D(N143), .LD(n5039), .CP(clk), .Q(N238)
         );
  FDS2L \Term2_reg[46]  ( .CR(1'b1), .D(N195), .LD(n5036), .CP(clk), .Q(
        Term2[46]) );
  FDS2L \Term1_reg[96]  ( .CR(1'b1), .D(N142), .LD(n5039), .CP(clk), .Q(N237)
         );
  FDS2L \Term1_reg[104]  ( .CR(1'b1), .D(N150), .LD(n5039), .CP(clk), .Q(
        Term1[104]) );
  FDS2L \Term3_reg[16]  ( .CR(1'b1), .D(N227), .LD(n5029), .CP(clk), .Q(
        Term3[16]) );
  FDS2L \Term2_reg[45]  ( .CR(1'b1), .D(N194), .LD(n5036), .CP(clk), .Q(
        Term2[45]) );
  FDS2L \Term1_reg[95]  ( .CR(1'b1), .D(N141), .LD(n5038), .CP(clk), .Q(N236)
         );
  FDS2L \Term2_reg[44]  ( .CR(1'b1), .D(N193), .LD(n5036), .CP(clk), .Q(
        Term2[44]) );
  FDS2L \Term3_reg[15]  ( .CR(1'b1), .D(N228), .LD(n5029), .CP(clk), .Q(
        Term3[15]) );
  FDS2L \Term1_reg[103]  ( .CR(1'b1), .D(N149), .LD(n5039), .CP(clk), .Q(
        Term1[103]) );
  FDS2L \Term1_reg[94]  ( .CR(1'b1), .D(N140), .LD(n5038), .CP(clk), .Q(N235)
         );
  FDS2L \Term3_reg[14]  ( .CR(1'b1), .D(N229), .LD(n5029), .CP(clk), .Q(
        Term3[14]) );
  FDS2L \Term1_reg[102]  ( .CR(1'b1), .D(N148), .LD(n5039), .CP(clk), .Q(
        Term1[102]) );
  FDS2L \Term2_reg[43]  ( .CR(1'b1), .D(N192), .LD(n5036), .CP(clk), .Q(
        Term2[43]) );
  FDS2L \Term1_reg[93]  ( .CR(1'b1), .D(N139), .LD(n5038), .CP(clk), .Q(N234)
         );
  FDS2L \Term2_reg[42]  ( .CR(1'b1), .D(N191), .LD(n5036), .CP(clk), .Q(
        Term2[42]) );
  FDS2L \Term1_reg[92]  ( .CR(1'b1), .D(N138), .LD(n5038), .CP(clk), .Q(N233)
         );
  FDS2L \Term2_reg[41]  ( .CR(1'b1), .D(N190), .LD(n5036), .CP(clk), .Q(
        Term2[41]) );
  FDS2L \Term1_reg[91]  ( .CR(1'b1), .D(N137), .LD(n5038), .CP(clk), .Q(N232)
         );
  FDS2L \Term2_reg[40]  ( .CR(1'b1), .D(N189), .LD(n5036), .CP(clk), .Q(
        Term2[40]) );
  FDS2L \Term1_reg[89]  ( .CR(1'b1), .D(N135), .LD(n5038), .CP(clk), .Q(N230)
         );
  FDS2L \Term1_reg[90]  ( .CR(1'b1), .D(N136), .LD(n5038), .CP(clk), .Q(N231)
         );
  FDS2L \Term2_reg[39]  ( .CR(1'b1), .D(N188), .LD(n5036), .CP(clk), .Q(
        Term2[39]) );
  FDS2L \Term2_reg[38]  ( .CR(1'b1), .D(N187), .LD(n5035), .CP(clk), .Q(
        Term2[38]) );
  FDS2L \LogIn2_reg[39]  ( .CR(1'b1), .D(LogIn[39]), .LD(n5044), .CP(clk), .Q(
        LogIn2[39]) );
  FDS2L \LogIn2_reg[38]  ( .CR(1'b1), .D(LogIn[38]), .LD(n5044), .CP(clk), .Q(
        LogIn2[38]) );
  FDS2L \LogIn2_reg[37]  ( .CR(1'b1), .D(LogIn[37]), .LD(n5044), .CP(clk), .Q(
        LogIn2[37]) );
  FDS2L \LogIn2_reg[36]  ( .CR(1'b1), .D(LogIn[36]), .LD(n5043), .CP(clk), .Q(
        LogIn2[36]) );
  FDS2L \LogIn2_reg[35]  ( .CR(1'b1), .D(LogIn[35]), .LD(n5043), .CP(clk), .Q(
        LogIn2[35]) );
  FDS2L \LogIn2_reg[34]  ( .CR(1'b1), .D(LogIn[34]), .LD(n5043), .CP(clk), .Q(
        LogIn2[34]) );
  FDS2L \LogIn2_reg[33]  ( .CR(1'b1), .D(LogIn[33]), .LD(n5043), .CP(clk), .Q(
        LogIn2[33]) );
  FDS2L \LogIn2_reg[32]  ( .CR(1'b1), .D(LogIn[32]), .LD(n5043), .CP(clk), .Q(
        LogIn2[32]) );
  FDS2L \LogIn2_reg[31]  ( .CR(1'b1), .D(LogIn[31]), .LD(n5043), .CP(clk), .Q(
        LogIn2[31]) );
  FDS2L \LogIn2_reg[30]  ( .CR(1'b1), .D(LogIn[30]), .LD(n5043), .CP(clk), .Q(
        LogIn2[30]) );
  FDS2L \LogIn2_reg[29]  ( .CR(1'b1), .D(LogIn[29]), .LD(n5043), .CP(clk), .Q(
        LogIn2[29]) );
  FDS2L \LogIn2_reg[28]  ( .CR(1'b1), .D(LogIn[28]), .LD(n5043), .CP(clk), .Q(
        LogIn2[28]) );
  FDS2L \LogIn2_reg[27]  ( .CR(1'b1), .D(LogIn[27]), .LD(n5043), .CP(clk), .Q(
        LogIn2[27]) );
  FDS2L \LogIn2_reg[26]  ( .CR(1'b1), .D(LogIn[26]), .LD(n5043), .CP(clk), .Q(
        LogIn2[26]) );
  FDS2L \LogIn2_reg[25]  ( .CR(1'b1), .D(LogIn[25]), .LD(n5043), .CP(clk), .Q(
        LogIn2[25]) );
  FDS2L \LogIn2_reg[24]  ( .CR(1'b1), .D(LogIn[24]), .LD(n5042), .CP(clk), .Q(
        LogIn2[24]) );
  FDS2L \LogIn2_reg[23]  ( .CR(1'b1), .D(LogIn[23]), .LD(n5042), .CP(clk), .Q(
        LogIn2[23]) );
  FDS2L \LogIn2_reg[22]  ( .CR(1'b1), .D(LogIn[22]), .LD(n5042), .CP(clk), .Q(
        LogIn2[22]) );
  FDS2L \LogIn2_reg[21]  ( .CR(1'b1), .D(LogIn[21]), .LD(n5042), .CP(clk), .Q(
        LogIn2[21]) );
  FDS2L \LogIn2_reg[20]  ( .CR(1'b1), .D(LogIn[20]), .LD(n5042), .CP(clk), .Q(
        LogIn2[20]) );
  FDS2L \LogIn2_reg[19]  ( .CR(1'b1), .D(LogIn[19]), .LD(n5042), .CP(clk), .Q(
        LogIn2[19]) );
  FDS2L \LogIn2_reg[18]  ( .CR(1'b1), .D(LogIn[18]), .LD(n5042), .CP(clk), .Q(
        LogIn2[18]) );
  FDS2L \LogIn2_reg[17]  ( .CR(1'b1), .D(LogIn[17]), .LD(n5042), .CP(clk), .Q(
        LogIn2[17]) );
  FDS2L \LogIn2_reg[16]  ( .CR(1'b1), .D(LogIn[16]), .LD(n5042), .CP(clk), .Q(
        LogIn2[16]) );
  FDS2L \LogIn2_reg[15]  ( .CR(1'b1), .D(LogIn[15]), .LD(n5042), .CP(clk), .Q(
        LogIn2[15]) );
  FDS2L \LogIn2_reg[14]  ( .CR(1'b1), .D(LogIn[14]), .LD(n5042), .CP(clk), .Q(
        LogIn2[14]) );
  FDS2L \LogIn2_reg[13]  ( .CR(1'b1), .D(LogIn[13]), .LD(n5042), .CP(clk), .Q(
        LogIn2[13]) );
  FDS2L \LogIn2_reg[11]  ( .CR(1'b1), .D(LogIn[11]), .LD(n5041), .CP(clk), .Q(
        LogIn2[11]) );
  FDS2L \LogIn2_reg[10]  ( .CR(1'b1), .D(LogIn[10]), .LD(n5041), .CP(clk), .Q(
        LogIn2[10]) );
  FDS2L \LogIn2_reg[9]  ( .CR(1'b1), .D(LogIn[9]), .LD(n5041), .CP(clk), .Q(
        LogIn2[9]) );
  FDS2L \LogIn2_reg[8]  ( .CR(1'b1), .D(LogIn[8]), .LD(n5041), .CP(clk), .Q(
        LogIn2[8]) );
  FDS2L \LogInSquare_reg[82]  ( .CR(1'b1), .D(N91), .LD(n5047), .CP(clk), .Q(
        LogInSquare[82]) );
  FDS2L \LogIn2_reg[7]  ( .CR(1'b1), .D(n22), .LD(n5041), .CP(clk), .Q(
        LogIn2[7]) );
  FDS2L \LogInSquare_reg[76]  ( .CR(1'b1), .D(N85), .LD(n5047), .CP(clk), .Q(
        LogInSquare[76]) );
  FDS2L \LogIn2_reg[6]  ( .CR(1'b1), .D(LogIn[6]), .LD(n5041), .CP(clk), .Q(
        LogIn2[6]) );
  FDS2L \LogInSquare_reg[79]  ( .CR(1'b1), .D(N88), .LD(n5047), .CP(clk), .Q(
        LogInSquare[79]) );
  FDS2L \LogInSquare_reg[78]  ( .CR(1'b1), .D(N87), .LD(n5047), .CP(clk), .Q(
        LogInSquare[78]) );
  FDS2L \LogInSquare_reg[75]  ( .CR(1'b1), .D(N84), .LD(n5047), .CP(clk), .Q(
        LogInSquare[75]) );
  FDS2L \LogInSquare_reg[74]  ( .CR(1'b1), .D(N83), .LD(n5047), .CP(clk), .Q(
        LogInSquare[74]) );
  FDS2L \LogInSquare_reg[71]  ( .CR(1'b1), .D(N80), .LD(n5046), .CP(clk), .Q(
        LogInSquare[71]) );
  FDS2L \LogInSquare_reg[70]  ( .CR(1'b1), .D(N79), .LD(n5046), .CP(clk), .Q(
        LogInSquare[70]) );
  FDS2L \LogInSquare_reg[57]  ( .CR(1'b1), .D(N66), .LD(n5045), .CP(clk), .Q(
        LogInSquare[57]) );
  FDS2L \LogInSquare_reg[56]  ( .CR(1'b1), .D(N65), .LD(n5045), .CP(clk), .Q(
        LogInSquare[56]) );
  FDS2L \LogInSquare_reg[30]  ( .CR(1'b1), .D(N39), .LD(n5027), .CP(clk), .Q(
        LogInSquare[30]) );
  FDS2L \LogInSquare_reg[1]  ( .CR(1'b1), .D(1'b0), .LD(n5025), .CP(clk), .Q(
        LogInSquare[1]) );
  FDS2L \LogInSquare_reg[67]  ( .CR(1'b1), .D(N76), .LD(n5046), .CP(clk), .Q(
        LogInSquare[67]) );
  FDS2L \LogInSquare_reg[66]  ( .CR(1'b1), .D(N75), .LD(n5046), .CP(clk), .Q(
        LogInSquare[66]) );
  FDS2L \LogInSquare_reg[63]  ( .CR(1'b1), .D(N72), .LD(n5046), .CP(clk), .Q(
        LogInSquare[63]) );
  FDS2L \LogInSquare_reg[62]  ( .CR(1'b1), .D(N71), .LD(n5046), .CP(clk), .Q(
        LogInSquare[62]) );
  FDS2L \LogInSquare_reg[60]  ( .CR(1'b1), .D(N69), .LD(n5046), .CP(clk), .Q(
        LogInSquare[60]) );
  FDS2L \LogInSquare_reg[55]  ( .CR(1'b1), .D(N64), .LD(n5045), .CP(clk), .Q(
        LogInSquare[55]) );
  FDS2L \LogIn2_reg[5]  ( .CR(1'b1), .D(LogIn[5]), .LD(n5041), .CP(clk), .Q(
        LogIn2[5]) );
  FDS2L \LogInSquare_reg[59]  ( .CR(1'b1), .D(N68), .LD(n5045), .CP(clk), .Q(
        LogInSquare[59]) );
  FDS2L \LogInSquare_reg[58]  ( .CR(1'b1), .D(N67), .LD(n5045), .CP(clk), .Q(
        LogInSquare[58]) );
  FDS2L \LogInSquare_reg[54]  ( .CR(1'b1), .D(N63), .LD(n5045), .CP(clk), .Q(
        LogInSquare[54]) );
  FDS2L \LogInSquare_reg[44]  ( .CR(1'b1), .D(N53), .LD(n5044), .CP(clk), .Q(
        LogInSquare[44]) );
  FDS2L \LogInSquare_reg[43]  ( .CR(1'b1), .D(N52), .LD(n5044), .CP(clk), .Q(
        LogInSquare[43]) );
  FDS2L \LogInSquare_reg[42]  ( .CR(1'b1), .D(N51), .LD(n5044), .CP(clk), .Q(
        LogInSquare[42]) );
  FDS2L \LogInSquare_reg[41]  ( .CR(1'b1), .D(N50), .LD(n5044), .CP(clk), .Q(
        LogInSquare[41]) );
  FDS2L \LogInSquare_reg[40]  ( .CR(1'b1), .D(N49), .LD(n5044), .CP(clk), .Q(
        LogInSquare[40]) );
  FDS2L \LogInSquare_reg[39]  ( .CR(1'b1), .D(N48), .LD(n5044), .CP(clk), .Q(
        LogInSquare[39]) );
  FDS2L \LogInSquare_reg[38]  ( .CR(1'b1), .D(N47), .LD(n5028), .CP(clk), .Q(
        LogInSquare[38]) );
  FDS2L \LogInSquare_reg[37]  ( .CR(1'b1), .D(N46), .LD(n5028), .CP(clk), .Q(
        LogInSquare[37]) );
  FDS2L \LogInSquare_reg[36]  ( .CR(1'b1), .D(N45), .LD(n5028), .CP(clk), .Q(
        LogInSquare[36]) );
  FDS2L \LogInSquare_reg[35]  ( .CR(1'b1), .D(N44), .LD(n5027), .CP(clk), .Q(
        LogInSquare[35]) );
  FDS2L \LogInSquare_reg[34]  ( .CR(1'b1), .D(N43), .LD(n5027), .CP(clk), .Q(
        LogInSquare[34]) );
  FDS2L \LogInSquare_reg[32]  ( .CR(1'b1), .D(N41), .LD(n5027), .CP(clk), .Q(
        LogInSquare[32]) );
  FDS2L \LogInSquare_reg[31]  ( .CR(1'b1), .D(N40), .LD(n5027), .CP(clk), .Q(
        LogInSquare[31]) );
  FDS2L \LogInSquare_reg[29]  ( .CR(1'b1), .D(N38), .LD(n5027), .CP(clk), .Q(
        LogInSquare[29]) );
  FDS2L \LogInSquare_reg[28]  ( .CR(1'b1), .D(N37), .LD(n5027), .CP(clk), .Q(
        LogInSquare[28]) );
  FDS2L \LogInSquare_reg[27]  ( .CR(1'b1), .D(N36), .LD(n5027), .CP(clk), .Q(
        LogInSquare[27]) );
  FDS2L \LogInSquare_reg[26]  ( .CR(1'b1), .D(N35), .LD(n5027), .CP(clk), .Q(
        LogInSquare[26]) );
  FDS2L \LogInSquare_reg[25]  ( .CR(1'b1), .D(N34), .LD(n5027), .CP(clk), .Q(
        LogInSquare[25]) );
  FDS2L \LogInSquare_reg[24]  ( .CR(1'b1), .D(N33), .LD(n5027), .CP(clk), .Q(
        LogInSquare[24]) );
  FDS2L \LogInSquare_reg[23]  ( .CR(1'b1), .D(N32), .LD(n5026), .CP(clk), .Q(
        LogInSquare[23]) );
  FDS2L \LogInSquare_reg[8]  ( .CR(1'b1), .D(N17), .LD(n5025), .CP(clk), .Q(
        LogInSquare[8]) );
  FDS2L \LogInSquare_reg[7]  ( .CR(1'b1), .D(N16), .LD(n5025), .CP(clk), .Q(
        LogInSquare[7]) );
  FDS2L \LogInSquare_reg[6]  ( .CR(1'b1), .D(N15), .LD(n5025), .CP(clk), .Q(
        LogInSquare[6]) );
  FDS2L \LogInSquare_reg[4]  ( .CR(1'b1), .D(N13), .LD(n5025), .CP(clk), .Q(
        LogInSquare[4]) );
  FDS2L \LogInSquare_reg[3]  ( .CR(1'b1), .D(N12), .LD(n5025), .CP(clk), .Q(
        LogInSquare[3]) );
  FDS2L \LogInSquare_reg[2]  ( .CR(1'b1), .D(N11), .LD(n5025), .CP(clk), .Q(
        LogInSquare[2]) );
  FDS2L \LogIn2_reg[4]  ( .CR(1'b1), .D(LogIn[4]), .LD(n5041), .CP(clk), .Q(
        LogIn2[4]) );
  FDS2L \LogIn2_reg[3]  ( .CR(1'b1), .D(LogIn[3]), .LD(n5041), .CP(clk), .Q(
        LogIn2[3]) );
  FDS2L \LogIn2_reg[2]  ( .CR(1'b1), .D(LogIn[2]), .LD(n5041), .CP(clk), .Q(
        LogIn2[2]) );
  FDS2L \LogInSquare_reg[53]  ( .CR(1'b1), .D(N62), .LD(n5045), .CP(clk), .Q(
        LogInSquare[53]) );
  FDS2L \LogInSquare_reg[52]  ( .CR(1'b1), .D(N61), .LD(n5045), .CP(clk), .Q(
        LogInSquare[52]) );
  FDS2L \LogInSquare_reg[51]  ( .CR(1'b1), .D(N60), .LD(n5045), .CP(clk), .Q(
        LogInSquare[51]) );
  FDS2L \LogInSquare_reg[50]  ( .CR(1'b1), .D(N59), .LD(n5045), .CP(clk), .Q(
        LogInSquare[50]) );
  FDS2L \LogInSquare_reg[49]  ( .CR(1'b1), .D(N58), .LD(n5045), .CP(clk), .Q(
        LogInSquare[49]) );
  FDS2L \LogInSquare_reg[48]  ( .CR(1'b1), .D(N57), .LD(n5045), .CP(clk), .Q(
        LogInSquare[48]) );
  FDS2L \LogInSquare_reg[47]  ( .CR(1'b1), .D(N56), .LD(n5044), .CP(clk), .Q(
        LogInSquare[47]) );
  FDS2L \LogInSquare_reg[46]  ( .CR(1'b1), .D(N55), .LD(n5044), .CP(clk), .Q(
        LogInSquare[46]) );
  FDS2L \LogInSquare_reg[45]  ( .CR(1'b1), .D(N54), .LD(n5044), .CP(clk), .Q(
        LogInSquare[45]) );
  FDS2L \LogInSquare_reg[22]  ( .CR(1'b1), .D(N31), .LD(n5026), .CP(clk), .Q(
        LogInSquare[22]) );
  FDS2L \LogInSquare_reg[21]  ( .CR(1'b1), .D(N30), .LD(n5026), .CP(clk), .Q(
        LogInSquare[21]) );
  FDS2L \LogInSquare_reg[20]  ( .CR(1'b1), .D(N29), .LD(n5026), .CP(clk), .Q(
        LogInSquare[20]) );
  FDS2L \LogInSquare_reg[18]  ( .CR(1'b1), .D(N27), .LD(n5026), .CP(clk), .Q(
        LogInSquare[18]) );
  FDS2L \LogInSquare_reg[17]  ( .CR(1'b1), .D(N26), .LD(n5026), .CP(clk), .Q(
        LogInSquare[17]) );
  FDS2L \LogInSquare_reg[16]  ( .CR(1'b1), .D(N25), .LD(n5026), .CP(clk), .Q(
        LogInSquare[16]) );
  FDS2L \LogInSquare_reg[15]  ( .CR(1'b1), .D(N24), .LD(n5026), .CP(clk), .Q(
        LogInSquare[15]) );
  FDS2L \LogInSquare_reg[14]  ( .CR(1'b1), .D(N23), .LD(n5026), .CP(clk), .Q(
        LogInSquare[14]) );
  FDS2L \LogInSquare_reg[13]  ( .CR(1'b1), .D(N22), .LD(n5026), .CP(clk), .Q(
        LogInSquare[13]) );
  FDS2L \LogInSquare_reg[12]  ( .CR(1'b1), .D(N21), .LD(n5026), .CP(clk), .Q(
        LogInSquare[12]) );
  FDS2L \LogInSquare_reg[11]  ( .CR(1'b1), .D(N20), .LD(n5025), .CP(clk), .Q(
        LogInSquare[11]) );
  FDS2L \LogInSquare_reg[10]  ( .CR(1'b1), .D(N19), .LD(n5025), .CP(clk), .Q(
        LogInSquare[10]) );
  FDS2L \LogInSquare_reg[9]  ( .CR(1'b1), .D(N18), .LD(n5025), .CP(clk), .Q(
        LogInSquare[9]) );
  FDS2L \LogInSquare_reg[5]  ( .CR(1'b1), .D(N14), .LD(n5025), .CP(clk), .Q(
        LogInSquare[5]) );
  FDS2L \LogInSquare_reg[19]  ( .CR(1'b1), .D(N28), .LD(n5026), .CP(clk), .Q(
        LogInSquare[19]) );
  FDS2L \FractionBit_reg[22]  ( .CR(1'b1), .D(N276), .LD(n5034), .CP(clk), .Q(
        FractionBit[22]) );
  FDS2L \FractionBit_reg[21]  ( .CR(1'b1), .D(N275), .LD(n5034), .CP(clk), .Q(
        FractionBit[21]) );
  FDS2L \FractionBit_reg[20]  ( .CR(1'b1), .D(N274), .LD(n5034), .CP(clk), .Q(
        FractionBit[20]) );
  FDS2L \FractionBit_reg[19]  ( .CR(1'b1), .D(N273), .LD(n5034), .CP(clk), .Q(
        FractionBit[19]) );
  FDS2L \FractionBit_reg[18]  ( .CR(1'b1), .D(N272), .LD(n5034), .CP(clk), .Q(
        FractionBit[18]) );
  FDS2L \FractionBit_reg[17]  ( .CR(1'b1), .D(N271), .LD(n5034), .CP(clk), .Q(
        FractionBit[17]) );
  FDS2L \FractionBit_reg[16]  ( .CR(1'b1), .D(N270), .LD(n5034), .CP(clk), .Q(
        FractionBit[16]) );
  FDS2L \FractionBit_reg[15]  ( .CR(1'b1), .D(N269), .LD(n5034), .CP(clk), .Q(
        FractionBit[15]) );
  FDS2L \FractionBit_reg[14]  ( .CR(1'b1), .D(N268), .LD(n5033), .CP(clk), .Q(
        FractionBit[14]) );
  FDS2L \FractionBit_reg[13]  ( .CR(1'b1), .D(N267), .LD(n5033), .CP(clk), .Q(
        FractionBit[13]) );
  FDS2L \FractionBit_reg[12]  ( .CR(1'b1), .D(N266), .LD(n5033), .CP(clk), .Q(
        FractionBit[12]) );
  FDS2L \FractionBit_reg[11]  ( .CR(1'b1), .D(N265), .LD(n5033), .CP(clk), .Q(
        FractionBit[11]) );
  FDS2L \FractionBit_reg[10]  ( .CR(1'b1), .D(N264), .LD(n5033), .CP(clk), .Q(
        FractionBit[10]) );
  FDS2L \FractionBit_reg[9]  ( .CR(1'b1), .D(N263), .LD(n5033), .CP(clk), .Q(
        FractionBit[9]) );
  FDS2L \FractionBit_reg[8]  ( .CR(1'b1), .D(N262), .LD(n5033), .CP(clk), .Q(
        FractionBit[8]) );
  FDS2L \FractionBit_reg[7]  ( .CR(1'b1), .D(N261), .LD(n5033), .CP(clk), .Q(
        FractionBit[7]) );
  FDS2L \FractionBit_reg[6]  ( .CR(1'b1), .D(N260), .LD(n5033), .CP(clk), .Q(
        FractionBit[6]) );
  FDS2L \FractionBit_reg[5]  ( .CR(1'b1), .D(N259), .LD(n5033), .CP(clk), .Q(
        FractionBit[5]) );
  FDS2L \FractionBit_reg[4]  ( .CR(1'b1), .D(N258), .LD(n5033), .CP(clk), .Q(
        FractionBit[4]) );
  FDS2L \FractionBit_reg[3]  ( .CR(1'b1), .D(N257), .LD(n5033), .CP(clk), .Q(
        FractionBit[3]) );
  FDS2L \FractionBit_reg[2]  ( .CR(1'b1), .D(N256), .LD(n5032), .CP(clk), .Q(
        FractionBit[2]) );
  FDS2L \FractionBit_reg[1]  ( .CR(1'b1), .D(N255), .LD(n5032), .CP(clk), .Q(
        FractionBit[1]) );
  FDS2L \FractionBit_reg[0]  ( .CR(1'b1), .D(N254), .LD(n5032), .CP(clk), .Q(
        FractionBit[0]) );
  FDS2L \IntegerBits_reg[6]  ( .CR(1'b1), .D(N298), .LD(n5032), .CP(clk), .Q(
        IntegerBits[6]) );
  FDS2L \IntegerBits_reg[5]  ( .CR(1'b1), .D(N297), .LD(n5032), .CP(clk), .Q(
        IntegerBits[5]) );
  FDS2L \IntegerBits_reg[4]  ( .CR(1'b1), .D(N296), .LD(n5032), .CP(clk), .Q(
        IntegerBits[4]) );
  FDS2L \IntegerBits_reg[3]  ( .CR(1'b1), .D(N295), .LD(n5032), .CP(clk), .Q(
        IntegerBits[3]) );
  FDS2L \IntegerBits_reg[2]  ( .CR(1'b1), .D(N294), .LD(n5032), .CP(clk), .Q(
        IntegerBits[2]) );
  FDS2L \IntegerBits_reg[1]  ( .CR(1'b1), .D(N293), .LD(n5032), .CP(clk), .Q(
        IntegerBits[1]) );
  FDS2L \IntegerBits_reg[0]  ( .CR(1'b1), .D(N292), .LD(n5032), .CP(clk), .Q(
        IntegerBits[0]) );
  FDS2L \Term1_reg[118]  ( .CR(1'b1), .D(N164), .LD(n5040), .CP(clk), .Q(
        Term1[118]) );
  FDS2L \Term1_reg[117]  ( .CR(1'b1), .D(N163), .LD(n5040), .CP(clk), .Q(
        Term1[117]) );
  FDS2L \Term1_reg[116]  ( .CR(1'b1), .D(N162), .LD(n5040), .CP(clk), .Q(
        Term1[116]) );
  FDS2L \Term1_reg[115]  ( .CR(1'b1), .D(N161), .LD(n5040), .CP(clk), .Q(
        Term1[115]) );
  FDS2L \Term1_reg[114]  ( .CR(1'b1), .D(N160), .LD(n5040), .CP(clk), .Q(
        Term1[114]) );
  FDS2L \Term1_reg[113]  ( .CR(1'b1), .D(N159), .LD(n5040), .CP(clk), .Q(
        Term1[113]) );
  FDS2L \Term1_reg[112]  ( .CR(1'b1), .D(N158), .LD(n5040), .CP(clk), .Q(
        Term1[112]) );
  FDS2L \Term2_reg[67]  ( .CR(1'b1), .D(N216), .LD(n5038), .CP(clk), .Q(
        Term2[67]) );
  FDS2L \Term2_reg[66]  ( .CR(1'b1), .D(N215), .LD(n5038), .CP(clk), .Q(
        Term2[66]) );
  FDS2L \Term2_reg[65]  ( .CR(1'b1), .D(N214), .LD(n5038), .CP(clk), .Q(
        Term2[65]) );
  FDS2L \Term2_reg[64]  ( .CR(1'b1), .D(N213), .LD(n5038), .CP(clk), .Q(
        Term2[64]) );
  FDS2L \Term2_reg[63]  ( .CR(1'b1), .D(N212), .LD(n5038), .CP(clk), .Q(
        Term2[63]) );
  FDS2L \Term2_reg[62]  ( .CR(1'b1), .D(N211), .LD(n5037), .CP(clk), .Q(
        Term2[62]) );
  FDS2L \Term2_reg[61]  ( .CR(1'b1), .D(N210), .LD(n5037), .CP(clk), .Q(
        Term2[61]) );
  FDS2L \Term3_reg[26]  ( .CR(1'b1), .D(n129), .LD(n5028), .CP(clk), .Q(
        Term3[26]) );
  FDS2L \Term3_reg[25]  ( .CR(1'b1), .D(N218), .LD(n5029), .CP(clk), .Q(
        Term3[25]) );
  FDS2L \Term3_reg[24]  ( .CR(1'b1), .D(N219), .LD(n5029), .CP(clk), .Q(
        Term3[24]) );
  FDS2L \LogOut_reg[20]  ( .CR(1'b1), .D(Log[19]), .LD(n5031), .CP(clk), .Q(
        LogOut[20]) );
  FDS2L \LogOut_reg[19]  ( .CR(1'b1), .D(Log[18]), .LD(n5031), .CP(clk), .Q(
        LogOut[19]) );
  FDS2L \LogOut_reg[18]  ( .CR(1'b1), .D(Log[17]), .LD(n5031), .CP(clk), .Q(
        LogOut[18]) );
  FDS2L \LogOut_reg[17]  ( .CR(1'b1), .D(Log[16]), .LD(n5031), .CP(clk), .Q(
        LogOut[17]) );
  FDS2L \LogOut_reg[16]  ( .CR(1'b1), .D(Log[15]), .LD(n5031), .CP(clk), .Q(
        LogOut[16]) );
  FDS2L \LogOut_reg[15]  ( .CR(1'b1), .D(Log[14]), .LD(n5031), .CP(clk), .Q(
        LogOut[15]) );
  FDS2L \LogOut_reg[14]  ( .CR(1'b1), .D(Log[13]), .LD(n5031), .CP(clk), .Q(
        LogOut[14]) );
  FDS2L \LogOut_reg[13]  ( .CR(1'b1), .D(Log[12]), .LD(n5031), .CP(clk), .Q(
        LogOut[13]) );
  FDS2L \LogOut_reg[12]  ( .CR(1'b1), .D(Log[11]), .LD(n5031), .CP(clk), .Q(
        LogOut[12]) );
  FDS2L \LogOut_reg[11]  ( .CR(1'b1), .D(Log[10]), .LD(n5031), .CP(clk), .Q(
        LogOut[11]) );
  FDS2L \LogOut_reg[10]  ( .CR(1'b1), .D(Log[9]), .LD(n5031), .CP(clk), .Q(
        LogOut[10]) );
  FDS2L \LogOut_reg[9]  ( .CR(1'b1), .D(Log[8]), .LD(n5030), .CP(clk), .Q(
        LogOut[9]) );
  FDS2L \LogOut_reg[8]  ( .CR(1'b1), .D(Log[7]), .LD(n5030), .CP(clk), .Q(
        LogOut[8]) );
  FDS2L \LogOut_reg[7]  ( .CR(1'b1), .D(Log[6]), .LD(n5030), .CP(clk), .Q(
        LogOut[7]) );
  FDS2L \LogOut_reg[6]  ( .CR(1'b1), .D(Log[5]), .LD(n5030), .CP(clk), .Q(
        LogOut[6]) );
  FDS2L \LogOut_reg[5]  ( .CR(1'b1), .D(Log[4]), .LD(n5030), .CP(clk), .Q(
        LogOut[5]) );
  FDS2L \LogOut_reg[4]  ( .CR(1'b1), .D(Log[3]), .LD(n5030), .CP(clk), .Q(
        LogOut[4]) );
  FDS2L \LogOut_reg[3]  ( .CR(1'b1), .D(Log[2]), .LD(n5030), .CP(clk), .Q(
        LogOut[3]) );
  FDS2L \LogOut_reg[2]  ( .CR(1'b1), .D(Log[1]), .LD(n5030), .CP(clk), .Q(
        LogOut[2]) );
  FDS2L \LogOut_reg[1]  ( .CR(1'b1), .D(Log[0]), .LD(n5030), .CP(clk), .Q(
        LogOut[1]) );
  FDS2L \LogIn2_reg[47]  ( .CR(1'b1), .D(LogIn[47]), .LD(n5071), .CP(clk), .Q(
        LogIn2[47]), .QN(n26) );
  FDS2L \LogIn2_reg[46]  ( .CR(1'b1), .D(LogIn[46]), .LD(n5071), .CP(clk), .Q(
        LogIn2[46]), .QN(n24) );
  FDS2L \LogIn2_reg[45]  ( .CR(1'b1), .D(LogIn[45]), .LD(n5071), .CP(clk), .Q(
        LogIn2[45]), .QN(n3932) );
  FDS2L \LogIn2_reg[44]  ( .CR(1'b1), .D(LogIn[44]), .LD(n5071), .CP(clk), .Q(
        LogIn2[44]), .QN(n23) );
  FDS2L \LogIn2_reg[43]  ( .CR(1'b1), .D(LogIn[43]), .LD(n5071), .CP(clk), .Q(
        LogIn2[43]) );
  FDS2L \LogIn2_reg[42]  ( .CR(1'b1), .D(LogIn[42]), .LD(n5071), .CP(clk), .Q(
        LogIn2[42]) );
  FDS2L \LogIn2_reg[41]  ( .CR(1'b1), .D(LogIn[41]), .LD(n5071), .CP(clk), .Q(
        LogIn2[41]) );
  FDS2L \LogIn2_reg[40]  ( .CR(1'b1), .D(LogIn[40]), .LD(n5071), .CP(clk), .Q(
        LogIn2[40]), .QN(n25) );
  FDS2L \LogInSquare_reg[0]  ( .CR(1'b1), .D(N9), .LD(n5071), .CP(clk), .Q(
        LogInSquare[0]) );
  FDS2L \Term31_reg[26]  ( .CR(1'b1), .D(Term3[26]), .LD(n5071), .CP(clk), .Q(
        Term31[26]) );
  FDS2L \Term31_reg[25]  ( .CR(1'b1), .D(Term3[25]), .LD(n5071), .CP(clk), .Q(
        Term31[25]) );
  FDS2L \Term31_reg[24]  ( .CR(1'b1), .D(Term3[24]), .LD(n5071), .CP(clk), .Q(
        Term31[24]) );
  FDS2L \Term21_reg[67]  ( .CR(1'b1), .D(Term2[67]), .LD(n5071), .CP(clk), .Q(
        Term21[67]) );
  FDS2L \Term21_reg[66]  ( .CR(1'b1), .D(Term2[66]), .LD(n5071), .CP(clk), .Q(
        Term21[66]) );
  FDS2L \Term21_reg[65]  ( .CR(1'b1), .D(Term2[65]), .LD(n5071), .CP(clk), .Q(
        Term21[65]) );
  FDS2L \Term21_reg[64]  ( .CR(1'b1), .D(Term2[64]), .LD(n5071), .CP(clk), .Q(
        Term21[64]) );
  FDS2L \Term21_reg[63]  ( .CR(1'b1), .D(Term2[63]), .LD(n5071), .CP(clk), .Q(
        Term21[63]) );
  FDS2L \Term21_reg[62]  ( .CR(1'b1), .D(Term2[62]), .LD(n5071), .CP(clk), .Q(
        Term21[62]) );
  FDS2L \Term21_reg[61]  ( .CR(1'b1), .D(Term2[61]), .LD(n5071), .CP(clk), .Q(
        Term21[61]) );
  FDS2L \Term11_reg[118]  ( .CR(1'b1), .D(Term1[118]), .LD(n5071), .CP(clk), 
        .Q(Term11[118]) );
  FDS2L \Term11_reg[117]  ( .CR(1'b1), .D(Term1[117]), .LD(n5071), .CP(clk), 
        .Q(Term11[117]) );
  FDS2L \Term11_reg[116]  ( .CR(1'b1), .D(Term1[116]), .LD(n5071), .CP(clk), 
        .Q(Term11[116]) );
  FDS2L \Term11_reg[115]  ( .CR(1'b1), .D(Term1[115]), .LD(n5071), .CP(clk), 
        .Q(Term11[115]) );
  FDS2L \Term11_reg[114]  ( .CR(1'b1), .D(Term1[114]), .LD(n5071), .CP(clk), 
        .Q(Term11[114]) );
  FDS2L \Term11_reg[113]  ( .CR(1'b1), .D(Term1[113]), .LD(n5071), .CP(clk), 
        .Q(Term11[113]) );
  FDS2L \Term11_reg[112]  ( .CR(1'b1), .D(Term1[112]), .LD(n5071), .CP(clk), 
        .Q(Term11[112]) );
  FDS2L \Log_reg[29]  ( .CR(1'b1), .D(IntegerBits[6]), .LD(n5071), .CP(clk), 
        .Q(Log[29]) );
  FDS2L \Log_reg[28]  ( .CR(1'b1), .D(IntegerBits[5]), .LD(n5071), .CP(clk), 
        .Q(Log[28]) );
  FDS2L \Log_reg[27]  ( .CR(1'b1), .D(IntegerBits[4]), .LD(n5071), .CP(clk), 
        .Q(Log[27]) );
  FDS2L \Log_reg[26]  ( .CR(1'b1), .D(IntegerBits[3]), .LD(n5071), .CP(clk), 
        .Q(Log[26]) );
  FDS2L \Log_reg[25]  ( .CR(1'b1), .D(IntegerBits[2]), .LD(n5071), .CP(clk), 
        .Q(Log[25]) );
  FDS2L \Log_reg[24]  ( .CR(1'b1), .D(IntegerBits[1]), .LD(n5071), .CP(clk), 
        .Q(Log[24]) );
  FDS2L \Log_reg[23]  ( .CR(1'b1), .D(IntegerBits[0]), .LD(n5071), .CP(clk), 
        .Q(Log[23]) );
  FDS2L \Log_reg[22]  ( .CR(1'b1), .D(LogPipe[22]), .LD(n5071), .CP(clk), .Q(
        Log[22]) );
  FDS2L \Log_reg[21]  ( .CR(1'b1), .D(LogPipe[21]), .LD(n5071), .CP(clk), .Q(
        Log[21]) );
  FDS2L \Log_reg[20]  ( .CR(1'b1), .D(LogPipe[20]), .LD(n5071), .CP(clk), .Q(
        Log[20]) );
  FDS2L \Log_reg[19]  ( .CR(1'b1), .D(LogPipe[19]), .LD(n5071), .CP(clk), .Q(
        Log[19]) );
  FDS2L \Log_reg[18]  ( .CR(1'b1), .D(LogPipe[18]), .LD(n5071), .CP(clk), .Q(
        Log[18]) );
  FDS2L \Log_reg[17]  ( .CR(1'b1), .D(LogPipe[17]), .LD(n5071), .CP(clk), .Q(
        Log[17]) );
  FDS2L \Log_reg[16]  ( .CR(1'b1), .D(LogPipe[16]), .LD(n5071), .CP(clk), .Q(
        Log[16]) );
  FDS2L \Log_reg[15]  ( .CR(1'b1), .D(LogPipe[15]), .LD(n5071), .CP(clk), .Q(
        Log[15]) );
  FDS2L \Log_reg[14]  ( .CR(1'b1), .D(LogPipe[14]), .LD(n5071), .CP(clk), .Q(
        Log[14]) );
  FDS2L \Log_reg[13]  ( .CR(1'b1), .D(LogPipe[13]), .LD(n5071), .CP(clk), .Q(
        Log[13]) );
  FDS2L \Log_reg[12]  ( .CR(1'b1), .D(LogPipe[12]), .LD(n5071), .CP(clk), .Q(
        Log[12]) );
  FDS2L \Log_reg[11]  ( .CR(1'b1), .D(LogPipe[11]), .LD(n5071), .CP(clk), .Q(
        Log[11]) );
  FDS2L \Log_reg[10]  ( .CR(1'b1), .D(LogPipe[10]), .LD(n5071), .CP(clk), .Q(
        Log[10]) );
  FDS2L \Log_reg[9]  ( .CR(1'b1), .D(LogPipe[9]), .LD(n5071), .CP(clk), .Q(
        Log[9]) );
  FDS2L \Log_reg[8]  ( .CR(1'b1), .D(LogPipe[8]), .LD(n5071), .CP(clk), .Q(
        Log[8]) );
  FDS2L \Log_reg[7]  ( .CR(1'b1), .D(LogPipe[7]), .LD(n5071), .CP(clk), .Q(
        Log[7]) );
  FDS2L \Log_reg[6]  ( .CR(1'b1), .D(LogPipe[6]), .LD(n5071), .CP(clk), .Q(
        Log[6]) );
  FDS2L \Log_reg[5]  ( .CR(1'b1), .D(LogPipe[5]), .LD(n5071), .CP(clk), .Q(
        Log[5]) );
  FDS2L \Log_reg[4]  ( .CR(1'b1), .D(LogPipe[4]), .LD(n5071), .CP(clk), .Q(
        Log[4]) );
  FDS2L \Log_reg[3]  ( .CR(1'b1), .D(LogPipe[3]), .LD(n5071), .CP(clk), .Q(
        Log[3]) );
  FDS2L \Log_reg[2]  ( .CR(1'b1), .D(LogPipe[2]), .LD(n5071), .CP(clk), .Q(
        Log[2]) );
  FDS2L \Log_reg[1]  ( .CR(1'b1), .D(LogPipe[1]), .LD(n5071), .CP(clk), .Q(
        Log[1]) );
  FDS2L \Log_reg[0]  ( .CR(1'b1), .D(LogPipe[0]), .LD(n5071), .CP(clk), .Q(
        Log[0]) );
  FDS2L \LogPipe_reg[22]  ( .CR(1'b1), .D(FractionBit[22]), .LD(n5071), .CP(
        clk), .Q(LogPipe[22]) );
  FDS2L \LogPipe_reg[21]  ( .CR(1'b1), .D(FractionBit[21]), .LD(n5071), .CP(
        clk), .Q(LogPipe[21]) );
  FDS2L \LogPipe_reg[20]  ( .CR(1'b1), .D(FractionBit[20]), .LD(n5071), .CP(
        clk), .Q(LogPipe[20]) );
  FDS2L \LogPipe_reg[19]  ( .CR(1'b1), .D(FractionBit[19]), .LD(n5071), .CP(
        clk), .Q(LogPipe[19]) );
  FDS2L \LogPipe_reg[18]  ( .CR(1'b1), .D(FractionBit[18]), .LD(n5071), .CP(
        clk), .Q(LogPipe[18]) );
  FDS2L \LogPipe_reg[17]  ( .CR(1'b1), .D(FractionBit[17]), .LD(n5071), .CP(
        clk), .Q(LogPipe[17]) );
  FDS2L \LogPipe_reg[16]  ( .CR(1'b1), .D(FractionBit[16]), .LD(n5071), .CP(
        clk), .Q(LogPipe[16]) );
  FDS2L \LogPipe_reg[15]  ( .CR(1'b1), .D(FractionBit[15]), .LD(n5071), .CP(
        clk), .Q(LogPipe[15]) );
  FDS2L \LogPipe_reg[14]  ( .CR(1'b1), .D(FractionBit[14]), .LD(n5071), .CP(
        clk), .Q(LogPipe[14]) );
  FDS2L \LogPipe_reg[13]  ( .CR(1'b1), .D(FractionBit[13]), .LD(n5071), .CP(
        clk), .Q(LogPipe[13]) );
  FDS2L \LogPipe_reg[12]  ( .CR(1'b1), .D(FractionBit[12]), .LD(n5071), .CP(
        clk), .Q(LogPipe[12]) );
  FDS2L \LogPipe_reg[11]  ( .CR(1'b1), .D(FractionBit[11]), .LD(n5071), .CP(
        clk), .Q(LogPipe[11]) );
  FDS2L \LogPipe_reg[10]  ( .CR(1'b1), .D(FractionBit[10]), .LD(n5071), .CP(
        clk), .Q(LogPipe[10]) );
  FDS2L \LogPipe_reg[9]  ( .CR(1'b1), .D(FractionBit[9]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[9]) );
  FDS2L \LogPipe_reg[8]  ( .CR(1'b1), .D(FractionBit[8]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[8]) );
  FDS2L \LogPipe_reg[7]  ( .CR(1'b1), .D(FractionBit[7]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[7]) );
  FDS2L \LogPipe_reg[6]  ( .CR(1'b1), .D(FractionBit[6]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[6]) );
  FDS2L \LogPipe_reg[5]  ( .CR(1'b1), .D(FractionBit[5]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[5]) );
  FDS2L \LogPipe_reg[4]  ( .CR(1'b1), .D(FractionBit[4]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[4]) );
  FDS2L \LogPipe_reg[3]  ( .CR(1'b1), .D(FractionBit[3]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[3]) );
  FDS2L \LogPipe_reg[2]  ( .CR(1'b1), .D(FractionBit[2]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[2]) );
  FDS2L \LogPipe_reg[1]  ( .CR(1'b1), .D(FractionBit[1]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[1]) );
  FDS2L \LogPipe_reg[0]  ( .CR(1'b1), .D(FractionBit[0]), .LD(n5071), .CP(clk), 
        .Q(LogPipe[0]) );
  FDS2L \LogOut_reg[30]  ( .CR(1'b1), .D(Log[29]), .LD(n5071), .CP(clk), .Q(
        LogOut[30]) );
  FDS2L \LogOut_reg[29]  ( .CR(1'b1), .D(Log[28]), .LD(n5071), .CP(clk), .Q(
        LogOut[29]) );
  FDS2L \LogOut_reg[28]  ( .CR(1'b1), .D(Log[27]), .LD(n5071), .CP(clk), .Q(
        LogOut[28]) );
  FDS2L \LogOut_reg[27]  ( .CR(1'b1), .D(Log[26]), .LD(n5071), .CP(clk), .Q(
        LogOut[27]) );
  FDS2L \LogOut_reg[26]  ( .CR(1'b1), .D(Log[25]), .LD(n5071), .CP(clk), .Q(
        LogOut[26]) );
  FDS2L \LogOut_reg[25]  ( .CR(1'b1), .D(Log[24]), .LD(n5071), .CP(clk), .Q(
        LogOut[25]) );
  FDS2L \LogOut_reg[24]  ( .CR(1'b1), .D(Log[23]), .LD(n5071), .CP(clk), .Q(
        LogOut[24]) );
  FDS2L \LogOut_reg[23]  ( .CR(1'b1), .D(Log[22]), .LD(n5071), .CP(clk), .Q(
        LogOut[23]) );
  FDS2L \LogOut_reg[22]  ( .CR(1'b1), .D(Log[21]), .LD(n5071), .CP(clk), .Q(
        LogOut[22]) );
  FDS2L \LogOut_reg[21]  ( .CR(1'b1), .D(Log[20]), .LD(n5071), .CP(clk), .Q(
        LogOut[21]) );
  MUX21LP U3 ( .A(LogInSquare[61]), .B(N70), .S(n5046), .Z(n448) );
  MUX21LP U4 ( .A(LogInSquare[65]), .B(N74), .S(n5046), .Z(n460) );
  B2I U5 ( .A(LogIn[0]), .Z2(n35) );
  MUX21LP U6 ( .A(LogInSquare[69]), .B(N78), .S(n5046), .Z(n466) );
  B5I U7 ( .A(n462), .Z(n463) );
  MUX21LP U8 ( .A(LogInSquare[95]), .B(N104), .S(n5048), .Z(n462) );
  B5I U9 ( .A(LogIn[7]), .Z(n21) );
  B4IP U10 ( .A(n21), .Z(n22) );
  NR3 U11 ( .A(n4015), .B(n437), .C(n3930), .Z(n3398) );
  NR3 U12 ( .A(n3925), .B(n4002), .C(n435), .Z(n3651) );
  NR2 U13 ( .A(n3999), .B(n436), .Z(n3781) );
  NR3 U14 ( .A(n3998), .B(n441), .C(n3928), .Z(n3502) );
  NR2 U15 ( .A(n3953), .B(n442), .Z(n3501) );
  NR2 U16 ( .A(n3929), .B(n440), .Z(n3443) );
  NR2 U17 ( .A(n4014), .B(n438), .Z(n3350) );
  NR2 U18 ( .A(n3928), .B(n439), .Z(n3465) );
  NR3 U19 ( .A(n443), .B(n4000), .C(n3955), .Z(n3590) );
  IVP U20 ( .A(n450), .Z(n451) );
  IVP U21 ( .A(n452), .Z(n453) );
  IVP U22 ( .A(n454), .Z(n455) );
  IVP U23 ( .A(n456), .Z(n457) );
  IVP U24 ( .A(n458), .Z(n459) );
  IVP U25 ( .A(n460), .Z(n461) );
  IVP U26 ( .A(n466), .Z(n467) );
  IVP U27 ( .A(n472), .Z(n473) );
  IVP U28 ( .A(n484), .Z(n485) );
  IVP U29 ( .A(n486), .Z(n487) );
  MUX21L U30 ( .A(LogInSquare[77]), .B(N86), .S(n5047), .Z(n486) );
  IVP U31 ( .A(n488), .Z(n489) );
  MUX21L U32 ( .A(LogInSquare[73]), .B(N82), .S(n5047), .Z(n488) );
  AN3 U33 ( .A(n3866), .B(n3875), .C(n75), .Z(n27) );
  AN3 U34 ( .A(n3866), .B(n3875), .C(n77), .Z(n28) );
  AN3 U35 ( .A(n3865), .B(n3874), .C(n78), .Z(n29) );
  AN3 U36 ( .A(n3868), .B(n3874), .C(n82), .Z(n30) );
  AN3 U37 ( .A(n3868), .B(n3874), .C(n83), .Z(n31) );
  AN3 U38 ( .A(n3868), .B(n3878), .C(n115), .Z(n32) );
  AN3 U39 ( .A(n3868), .B(n3878), .C(n116), .Z(n33) );
  AN3 U40 ( .A(n3868), .B(n3877), .C(n117), .Z(n34) );
  MUX21H U41 ( .A(LogInSquare[68]), .B(N77), .S(n5046), .Z(n36) );
  AN2P U42 ( .A(n2648), .B(n2647), .Z(n37) );
  AN2P U43 ( .A(n2522), .B(n2521), .Z(n38) );
  AN2P U44 ( .A(n2786), .B(n2785), .Z(n39) );
  AN2P U45 ( .A(n2092), .B(n4191), .Z(n40) );
  AN2P U46 ( .A(n2561), .B(n2560), .Z(n41) );
  MUX21H U47 ( .A(n2677), .B(n2676), .S(n4902), .Z(n42) );
  MUX21H U48 ( .A(n2181), .B(n4140), .S(n4567), .Z(n43) );
  MUX21H U49 ( .A(n4295), .B(n1979), .S(n4924), .Z(n44) );
  AN2P U50 ( .A(n1992), .B(n1991), .Z(n45) );
  AN2P U51 ( .A(n1825), .B(n1824), .Z(n46) );
  AN2P U52 ( .A(n2183), .B(n2182), .Z(n47) );
  AN2P U53 ( .A(n2317), .B(n2316), .Z(n48) );
  MUX21H U54 ( .A(n2756), .B(n2755), .S(n4244), .Z(n49) );
  AN3 U55 ( .A(n2547), .B(n2546), .C(n2545), .Z(n50) );
  AN3 U56 ( .A(n3150), .B(n3149), .C(n3148), .Z(n51) );
  AN2P U57 ( .A(n3222), .B(n3221), .Z(n52) );
  AN2P U58 ( .A(n1965), .B(n1964), .Z(n53) );
  AN2P U59 ( .A(n2017), .B(n4197), .Z(n54) );
  AN2P U60 ( .A(n1939), .B(n1938), .Z(n55) );
  MUX21H U61 ( .A(n4537), .B(n1976), .S(n4294), .Z(n56) );
  AN3 U62 ( .A(n2733), .B(n2732), .C(n2731), .Z(n57) );
  AN2P U63 ( .A(n4197), .B(n4541), .Z(n58) );
  AN3 U64 ( .A(n3929), .B(n3421), .C(n3420), .Z(n59) );
  AN2P U65 ( .A(n2692), .B(n2691), .Z(n60) );
  MUX21H U66 ( .A(n4480), .B(n2707), .S(n4213), .Z(n61) );
  AN2P U67 ( .A(n3296), .B(n3295), .Z(n62) );
  AN3 U68 ( .A(n3867), .B(n3877), .C(n760), .Z(n63) );
  AN3 U69 ( .A(n3866), .B(n3876), .C(n757), .Z(n64) );
  AN2P U70 ( .A(n3244), .B(n3243), .Z(n65) );
  MUX21H U71 ( .A(n3161), .B(n3160), .S(n4908), .Z(n66) );
  AN3 U72 ( .A(n3869), .B(n3880), .C(n1172), .Z(n67) );
  AN2P U73 ( .A(n3223), .B(n4587), .Z(n68) );
  AN3 U74 ( .A(n3869), .B(n3880), .C(n1167), .Z(n69) );
  AN3 U75 ( .A(n3866), .B(n3876), .C(n755), .Z(n70) );
  MUX21H U76 ( .A(n4253), .B(n4446), .S(n4906), .Z(n71) );
  AN3 U77 ( .A(n3869), .B(n3874), .C(n1164), .Z(n72) );
  MUX21H U78 ( .A(n4254), .B(n3113), .S(n4582), .Z(n73) );
  MUX21H U79 ( .A(n3225), .B(n3224), .S(n4911), .Z(n74) );
  AN4P U80 ( .A(n753), .B(n3896), .C(n3943), .D(n3979), .Z(n75) );
  MUX21H U81 ( .A(n4782), .B(n4233), .S(n4584), .Z(n76) );
  AN4P U82 ( .A(n752), .B(n3894), .C(n3946), .D(n3980), .Z(n77) );
  AN4P U83 ( .A(n751), .B(n3895), .C(n3943), .D(n3980), .Z(n78) );
  AN4P U84 ( .A(n4001), .B(n1161), .C(n3900), .D(n3944), .Z(n79) );
  AN3 U85 ( .A(n3868), .B(n3879), .C(n1159), .Z(n80) );
  AN3 U86 ( .A(n3868), .B(n3879), .C(n1157), .Z(n81) );
  AN4P U87 ( .A(n1154), .B(n3899), .C(n3950), .D(n3982), .Z(n82) );
  AN4P U88 ( .A(n1153), .B(n3898), .C(n3944), .D(n3982), .Z(n83) );
  AN4P U89 ( .A(n1152), .B(n3898), .C(n3946), .D(n3982), .Z(n115) );
  AN4P U90 ( .A(n1151), .B(n3897), .C(n3944), .D(n3981), .Z(n116) );
  AN4P U91 ( .A(n1150), .B(n3897), .C(n3947), .D(n3981), .Z(n117) );
  AN2P U92 ( .A(Term3[14]), .B(Term1[102]), .Z(n118) );
  AN4P U93 ( .A(n3673), .B(n3672), .C(n3671), .D(n3670), .Z(n119) );
  AN2P U94 ( .A(n1998), .B(n1997), .Z(n120) );
  AN2P U95 ( .A(n3256), .B(n3255), .Z(n121) );
  AN4P U96 ( .A(n3683), .B(n3682), .C(n3681), .D(n3680), .Z(n122) );
  MUX21H U97 ( .A(n4589), .B(n4239), .S(n4912), .Z(n123) );
  AN2P U98 ( .A(n2160), .B(n2159), .Z(n124) );
  MUX21H U99 ( .A(n2323), .B(n4633), .S(n4288), .Z(n125) );
  AN3 U100 ( .A(n2001), .B(n2000), .C(n1999), .Z(n126) );
  MUX21H U101 ( .A(n2011), .B(n2010), .S(n4925), .Z(n127) );
  AN4P U102 ( .A(n508), .B(n3908), .C(n3949), .D(n3990), .Z(n128) );
  AN3 U103 ( .A(n3865), .B(n3874), .C(n490), .Z(n129) );
  MUX21LP U193 ( .A(LogInSquare[80]), .B(N89), .S(n5047), .Z(n484) );
  B2I U194 ( .A(LogIn[1]), .Z2(n405) );
  MUX21LP U195 ( .A(LogInSquare[81]), .B(N90), .S(n5047), .Z(n472) );
  MUX21LP U196 ( .A(LogInSquare[94]), .B(N103), .S(n5048), .Z(n458) );
  MUX21LP U197 ( .A(LogInSquare[93]), .B(N102), .S(n5048), .Z(n456) );
  MUX21LP U198 ( .A(LogInSquare[91]), .B(N100), .S(n5048), .Z(n452) );
  MUX21LP U199 ( .A(LogInSquare[92]), .B(N101), .S(n5048), .Z(n454) );
  MUX21LP U200 ( .A(LogInSquare[90]), .B(N99), .S(n5048), .Z(n450) );
  ND2 U201 ( .A(n2620), .B(n2619), .Z(n1642) );
  ND2 U202 ( .A(n4949), .B(n4213), .Z(n2619) );
  EN U203 ( .A(n4563), .B(n4211), .Z(n2620) );
  NR2 U204 ( .A(n4946), .B(n4595), .Z(n2520) );
  EO U205 ( .A(n4888), .B(n4273), .Z(n1684) );
  EN U206 ( .A(n4566), .B(n4223), .Z(n2419) );
  ND2 U207 ( .A(n4941), .B(n4223), .Z(n2418) );
  ND2 U208 ( .A(n1691), .B(n1690), .Z(n1622) );
  EN U209 ( .A(n4565), .B(n4291), .Z(n1691) );
  EN U210 ( .A(n4890), .B(n4291), .Z(n1690) );
  ND2 U211 ( .A(n1930), .B(n1929), .Z(n1628) );
  ND2 U212 ( .A(n1926), .B(n4940), .Z(n1929) );
  MUX21L U213 ( .A(n1927), .B(n1928), .S(n4291), .Z(n1930) );
  NR2 U214 ( .A(n4626), .B(n4291), .Z(n1926) );
  NR2 U215 ( .A(n4901), .B(n4243), .Z(n2749) );
  NR2 U216 ( .A(n4922), .B(n4626), .Z(n1928) );
  EO U217 ( .A(n4888), .B(n4580), .Z(n1093) );
  EN U218 ( .A(n4562), .B(n4231), .Z(n1618) );
  EN U219 ( .A(n4888), .B(n4247), .Z(n1613) );
  ND2 U220 ( .A(n3257), .B(n4239), .Z(n1688) );
  EO U221 ( .A(n4892), .B(n4589), .Z(n3257) );
  ND2 U222 ( .A(n3121), .B(n3120), .Z(n1686) );
  EN U223 ( .A(n4884), .B(n4254), .Z(n3121) );
  ND2 U224 ( .A(n4582), .B(n4248), .Z(n3120) );
  ND2 U225 ( .A(n2742), .B(n2741), .Z(n1138) );
  ND2 U226 ( .A(n4604), .B(n4243), .Z(n2741) );
  MUX21L U227 ( .A(n2740), .B(n4243), .S(n4898), .Z(n2742) );
  NR2 U228 ( .A(n4604), .B(n4243), .Z(n2740) );
  ND2 U229 ( .A(n2500), .B(n4227), .Z(n1134) );
  EO U230 ( .A(n4893), .B(n4594), .Z(n2500) );
  ND2 U231 ( .A(n1780), .B(n1779), .Z(n1118) );
  ND2 U232 ( .A(n1776), .B(n4935), .Z(n1779) );
  MUX21L U233 ( .A(n1777), .B(n1778), .S(n4935), .Z(n1780) );
  NR2 U234 ( .A(n4575), .B(n4264), .Z(n1776) );
  ND2 U235 ( .A(n2467), .B(n2466), .Z(n1100) );
  EN U236 ( .A(n4885), .B(n4225), .Z(n2467) );
  EO U237 ( .A(n4566), .B(n4225), .Z(n2466) );
  ND2 U238 ( .A(n4577), .B(n4262), .Z(n1820) );
  ND2 U239 ( .A(n2587), .B(n2586), .Z(n1610) );
  MUX21L U240 ( .A(n2584), .B(n2585), .S(n4948), .Z(n2586) );
  MUX21L U241 ( .A(n2582), .B(n2583), .S(n4632), .Z(n2587) );
  NR2 U242 ( .A(n4631), .B(n4213), .Z(n2584) );
  ND2 U243 ( .A(n3258), .B(n4589), .Z(n1620) );
  EO U244 ( .A(n4891), .B(n4240), .Z(n3258) );
  MUX21L U245 ( .A(n4299), .B(n4927), .S(n4640), .Z(n1665) );
  AO4 U246 ( .A(n4636), .B(n4285), .C(n4953), .D(n4285), .Z(n1095) );
  NR2 U247 ( .A(n4577), .B(n4278), .Z(n2095) );
  NR2 U248 ( .A(n4939), .B(n4628), .Z(n1595) );
  EO U249 ( .A(n4890), .B(n4571), .Z(n1591) );
  EO U250 ( .A(n4562), .B(n4245), .Z(n2786) );
  ND3 U251 ( .A(n2784), .B(n2783), .C(n2782), .Z(n1105) );
  ND2 U252 ( .A(n4601), .B(n4902), .Z(n2784) );
  ND2 U253 ( .A(n4902), .B(n4245), .Z(n2783) );
  ND2 U254 ( .A(n4601), .B(n4245), .Z(n2782) );
  ND2 U255 ( .A(n4577), .B(n4262), .Z(n1812) );
  ND2 U256 ( .A(n4617), .B(n4251), .Z(n2875) );
  ND2 U257 ( .A(n4907), .B(n3124), .Z(n1112) );
  ND2 U258 ( .A(n4582), .B(n4231), .Z(n3124) );
  ND2 U259 ( .A(n4283), .B(n2225), .Z(n1603) );
  ND2 U260 ( .A(n4952), .B(n4637), .Z(n2225) );
  ND2 U261 ( .A(n4607), .B(n4215), .Z(n2676) );
  ND2 U262 ( .A(n3011), .B(n3010), .Z(n1077) );
  ND2 U263 ( .A(n3007), .B(n4920), .Z(n3010) );
  MUX21L U264 ( .A(n3008), .B(n3009), .S(n4269), .Z(n3011) );
  NR2 U265 ( .A(n4598), .B(n4268), .Z(n3007) );
  AN2P U266 ( .A(n4607), .B(n4216), .Z(n406) );
  MUX21L U267 ( .A(n4923), .B(n4624), .S(n4294), .Z(n1123) );
  MUX21L U268 ( .A(n4224), .B(n2447), .S(n4592), .Z(n1608) );
  ND2 U269 ( .A(n4942), .B(n4224), .Z(n2447) );
  MUX21L U270 ( .A(n4264), .B(n1775), .S(n4935), .Z(n1592) );
  ND2 U271 ( .A(n4575), .B(n4264), .Z(n1775) );
  NR2 U272 ( .A(n4580), .B(n4256), .Z(n2147) );
  NR2 U273 ( .A(n4920), .B(n4598), .Z(n3009) );
  ND2 U274 ( .A(n1707), .B(n1706), .Z(n1555) );
  MUX21L U275 ( .A(n1704), .B(n1705), .S(n4932), .Z(n1706) );
  MUX21L U276 ( .A(n1702), .B(n1703), .S(n4571), .Z(n1707) );
  NR2 U277 ( .A(n4571), .B(n4290), .Z(n1704) );
  ND2 U278 ( .A(n1867), .B(n4259), .Z(n1056) );
  EO U279 ( .A(n4893), .B(n4629), .Z(n1867) );
  ND2 U280 ( .A(n2833), .B(n2832), .Z(n1074) );
  ND2 U281 ( .A(n4248), .B(n4619), .Z(n2832) );
  MUX21L U282 ( .A(n2831), .B(n4619), .S(n4896), .Z(n2833) );
  NR2 U283 ( .A(n4619), .B(n4248), .Z(n2831) );
  AO4 U284 ( .A(n4593), .B(n4225), .C(n4943), .D(n4225), .Z(n1574) );
  NR2 U285 ( .A(n4916), .B(n4275), .Z(n2922) );
  NR2 U286 ( .A(n4921), .B(n4267), .Z(n3042) );
  NR2 U287 ( .A(n4947), .B(n4229), .Z(n2551) );
  NR2 U288 ( .A(n4900), .B(n4246), .Z(n2803) );
  EN U289 ( .A(n4887), .B(n4300), .Z(n2062) );
  MUX21L U290 ( .A(n2055), .B(n4927), .S(n4299), .Z(n1564) );
  ND2 U291 ( .A(n4927), .B(n4640), .Z(n2055) );
  ND2 U292 ( .A(n2074), .B(n2073), .Z(n1028) );
  ND2 U293 ( .A(n2070), .B(n4928), .Z(n2073) );
  MUX21L U294 ( .A(n2071), .B(n2072), .S(n4928), .Z(n2074) );
  NR2 U295 ( .A(n4639), .B(n4295), .Z(n2070) );
  AO4 U296 ( .A(n4580), .B(n4291), .C(n4932), .D(n4291), .Z(n1018) );
  AO7 U297 ( .A(n4900), .B(n4217), .C(n4605), .Z(n1042) );
  NR2 U298 ( .A(n4940), .B(n4569), .Z(n2387) );
  NR2 U299 ( .A(n4935), .B(n4265), .Z(n1758) );
  EO U300 ( .A(n4564), .B(n4223), .Z(n1537) );
  ND2 U301 ( .A(n3212), .B(n4911), .Z(n1552) );
  EN U302 ( .A(n4565), .B(n4237), .Z(n3212) );
  ND2 U303 ( .A(n1832), .B(n4261), .Z(n1524) );
  EN U304 ( .A(n4892), .B(n4631), .Z(n1832) );
  ND2 U305 ( .A(n4568), .B(n4222), .Z(n1036) );
  NR2 U306 ( .A(n4581), .B(n4252), .Z(n3075) );
  NR2 U307 ( .A(n4905), .B(n4581), .Z(n3077) );
  ND2 U308 ( .A(n3012), .B(n4268), .Z(n1014) );
  EN U309 ( .A(n4886), .B(n4598), .Z(n3012) );
  ND2 U310 ( .A(n2243), .B(n2242), .Z(n997) );
  EN U311 ( .A(n4889), .B(n4284), .Z(n2243) );
  EO U312 ( .A(n4566), .B(n4284), .Z(n2242) );
  ND2 U313 ( .A(n2264), .B(n2263), .Z(n998) );
  EN U314 ( .A(n4566), .B(n4285), .Z(n2264) );
  EN U315 ( .A(n4889), .B(n4285), .Z(n2263) );
  MUX21L U316 ( .A(n2754), .B(n4603), .S(n4244), .Z(n1008) );
  ND2 U317 ( .A(n4902), .B(n4603), .Z(n2754) );
  MUX21L U318 ( .A(n4597), .B(n4270), .S(n4919), .Z(n1549) );
  ND2 U319 ( .A(n1888), .B(n1887), .Z(n1489) );
  ND2 U320 ( .A(n4628), .B(n4258), .Z(n1887) );
  EO U321 ( .A(n4893), .B(n4258), .Z(n1888) );
  EN U322 ( .A(n4890), .B(n4240), .Z(n1518) );
  ND2 U323 ( .A(n4627), .B(n4257), .Z(n990) );
  NR2 U324 ( .A(n4573), .B(n4260), .Z(n1744) );
  ND2 U325 ( .A(n2099), .B(n4577), .Z(n1496) );
  EN U326 ( .A(n4887), .B(n4279), .Z(n2099) );
  ND2 U327 ( .A(n4940), .B(n4257), .Z(n1919) );
  MUX21L U328 ( .A(n4255), .B(n2167), .S(n4950), .Z(n1497) );
  ND2 U329 ( .A(n4576), .B(n4255), .Z(n2167) );
  ND2 U330 ( .A(n4919), .B(n4270), .Z(n1515) );
  NR2 U331 ( .A(n4595), .B(n4228), .Z(n2526) );
  ND2 U332 ( .A(n4586), .B(n3191), .Z(n985) );
  ND2 U333 ( .A(n4910), .B(n4235), .Z(n3191) );
  ND2 U334 ( .A(n2504), .B(n2503), .Z(n974) );
  ND2 U335 ( .A(n4594), .B(n4945), .Z(n2504) );
  ND2 U336 ( .A(n4945), .B(n4227), .Z(n2503) );
  ND2 U337 ( .A(n2628), .B(n2627), .Z(n1473) );
  ND2 U338 ( .A(n4609), .B(n4212), .Z(n2627) );
  EN U339 ( .A(n4890), .B(n4212), .Z(n2628) );
  ND2 U340 ( .A(n2737), .B(n4896), .Z(n1475) );
  EO U341 ( .A(n4561), .B(n4242), .Z(n2737) );
  ND2 U342 ( .A(n2781), .B(n4902), .Z(n1476) );
  EO U343 ( .A(n4562), .B(n4245), .Z(n2781) );
  ND2 U344 ( .A(n1890), .B(n1889), .Z(n1457) );
  ND2 U345 ( .A(n4939), .B(n4258), .Z(n1889) );
  EO U346 ( .A(n4565), .B(n4258), .Z(n1890) );
  EO U347 ( .A(n4891), .B(n4266), .Z(n1455) );
  ND2 U348 ( .A(n2824), .B(n4619), .Z(n1478) );
  EO U349 ( .A(n4888), .B(n4248), .Z(n2824) );
  ND2 U350 ( .A(n4573), .B(n4934), .Z(n1734) );
  ND2 U351 ( .A(n2169), .B(n2168), .Z(n1464) );
  ND2 U352 ( .A(n4950), .B(n4255), .Z(n2168) );
  ND2 U353 ( .A(n4567), .B(n4950), .Z(n2169) );
  MUX21L U354 ( .A(n4235), .B(n3190), .S(n4909), .Z(n1483) );
  ND2 U355 ( .A(n4585), .B(n4235), .Z(n3190) );
  ND2 U356 ( .A(n4899), .B(n4605), .Z(n978) );
  NR2 U357 ( .A(n4934), .B(n4265), .Z(n1748) );
  NR2 U358 ( .A(n4622), .B(n4297), .Z(n1461) );
  ND2 U359 ( .A(n2577), .B(n2576), .Z(n944) );
  ND2 U360 ( .A(n4632), .B(n4225), .Z(n2576) );
  EO U361 ( .A(n4891), .B(n4210), .Z(n2577) );
  EN U362 ( .A(n4892), .B(n4262), .Z(n931) );
  ND2 U363 ( .A(n4927), .B(n4299), .Z(n1462) );
  ND2 U364 ( .A(n4951), .B(n4271), .Z(n2182) );
  ND2 U365 ( .A(n4924), .B(n4624), .Z(n1980) );
  MUX21L U366 ( .A(n4217), .B(n4605), .S(n4897), .Z(n946) );
  ND2 U367 ( .A(n1740), .B(n1739), .Z(n1421) );
  ND2 U368 ( .A(n1736), .B(n4934), .Z(n1739) );
  MUX21L U369 ( .A(n1737), .B(n1738), .S(n4934), .Z(n1740) );
  NR2 U370 ( .A(n4573), .B(n4289), .Z(n1736) );
  NR2 U371 ( .A(n4901), .B(n4601), .Z(n2791) );
  ND2 U372 ( .A(n2999), .B(n4597), .Z(n1448) );
  EN U373 ( .A(n4887), .B(n4269), .Z(n2999) );
  ND2 U374 ( .A(n3129), .B(n3128), .Z(n1449) );
  ND2 U375 ( .A(n4907), .B(n4231), .Z(n3128) );
  EN U376 ( .A(n4884), .B(n4583), .Z(n3129) );
  ND2 U377 ( .A(n2669), .B(n4607), .Z(n1440) );
  EO U378 ( .A(n4891), .B(n4215), .Z(n2669) );
  ND2 U379 ( .A(n4589), .B(n3261), .Z(n1451) );
  ND2 U380 ( .A(n4912), .B(n4240), .Z(n3261) );
  ND2 U381 ( .A(n2622), .B(n2621), .Z(n1439) );
  ND2 U382 ( .A(n4610), .B(n4949), .Z(n2622) );
  ND2 U383 ( .A(n4949), .B(n4211), .Z(n2621) );
  ND2 U384 ( .A(n2231), .B(n4952), .Z(n2234) );
  NR2 U385 ( .A(n4637), .B(n4283), .Z(n2231) );
  AO4 U386 ( .A(n4946), .B(n4228), .C(n4946), .D(n4595), .Z(n1438) );
  NR2 U387 ( .A(n4937), .B(n4260), .Z(n1843) );
  ND2 U388 ( .A(n4603), .B(n4902), .Z(n2756) );
  ND2 U389 ( .A(n3272), .B(n3271), .Z(n927) );
  ND2 U390 ( .A(n4240), .B(n4913), .Z(n3271) );
  MUX21L U391 ( .A(n3270), .B(n4590), .S(n4913), .Z(n3272) );
  NR2 U392 ( .A(n4590), .B(n4240), .Z(n3270) );
  AO4 U393 ( .A(n4621), .B(n4247), .C(n4899), .D(n4621), .Z(n921) );
  EO U394 ( .A(n4885), .B(n4243), .Z(n1410) );
  EO U395 ( .A(n4886), .B(n4622), .Z(n1396) );
  ND2 U396 ( .A(n2469), .B(n2468), .Z(n1405) );
  ND2 U397 ( .A(n4943), .B(n4225), .Z(n2468) );
  EN U398 ( .A(n4885), .B(n4592), .Z(n2469) );
  ND2 U399 ( .A(n4274), .B(n2928), .Z(n923) );
  ND2 U400 ( .A(n4916), .B(n4614), .Z(n2928) );
  MUX21L U401 ( .A(n4598), .B(n4268), .S(n4920), .Z(n925) );
  NR2 U402 ( .A(n4894), .B(n4250), .Z(n2857) );
  NR2 U403 ( .A(n4944), .B(n4226), .Z(n2492) );
  ND3 U404 ( .A(n2684), .B(n2683), .C(n2682), .Z(n1408) );
  ND2 U405 ( .A(n4903), .B(n4216), .Z(n2683) );
  ND2 U406 ( .A(n4607), .B(n4903), .Z(n2684) );
  ND2 U407 ( .A(n4607), .B(n4216), .Z(n2682) );
  ND3 U408 ( .A(n4601), .B(n4246), .C(n4901), .Z(n1412) );
  ND2 U409 ( .A(n4928), .B(n2077), .Z(n1397) );
  ND2 U410 ( .A(n4639), .B(n4277), .Z(n2077) );
  ND2 U411 ( .A(n1892), .B(n1891), .Z(n875) );
  ND2 U412 ( .A(n4939), .B(n4258), .Z(n1891) );
  EO U413 ( .A(n4565), .B(n4258), .Z(n1892) );
  ND2 U414 ( .A(n3287), .B(n3286), .Z(n899) );
  EN U415 ( .A(n4890), .B(n4241), .Z(n3287) );
  EO U416 ( .A(n4564), .B(n4241), .Z(n3286) );
  ND2 U417 ( .A(n2177), .B(n2176), .Z(n882) );
  ND2 U418 ( .A(n2173), .B(n4951), .Z(n2176) );
  MUX21L U419 ( .A(n2174), .B(n2175), .S(n4951), .Z(n2177) );
  NR2 U420 ( .A(n4567), .B(n4254), .Z(n2173) );
  ND2 U421 ( .A(n4281), .B(n4579), .Z(n2139) );
  ND2 U422 ( .A(n4927), .B(n4641), .Z(n2042) );
  MUX21L U423 ( .A(n2138), .B(n4579), .S(n4931), .Z(n2140) );
  NR2 U424 ( .A(n4579), .B(n4281), .Z(n2138) );
  MUX21L U425 ( .A(n4250), .B(n2868), .S(n4617), .Z(n894) );
  ND2 U426 ( .A(n4893), .B(n4250), .Z(n2868) );
  ND2 U427 ( .A(n3204), .B(n3203), .Z(n1387) );
  ND2 U428 ( .A(n4910), .B(n4236), .Z(n3203) );
  EO U429 ( .A(n4565), .B(n4236), .Z(n3204) );
  EN U430 ( .A(n4566), .B(n4274), .Z(n1383) );
  ND2 U431 ( .A(n2637), .B(n2636), .Z(n1377) );
  ND2 U432 ( .A(n4940), .B(n4213), .Z(n2636) );
  EO U433 ( .A(n4561), .B(n4213), .Z(n2637) );
  ND2 U434 ( .A(n2450), .B(n4592), .Z(n1374) );
  EO U435 ( .A(n4886), .B(n4224), .Z(n2450) );
  EO U436 ( .A(n4563), .B(n4281), .Z(n1369) );
  EO U437 ( .A(n4887), .B(n4640), .Z(n1367) );
  ND2 U438 ( .A(n4905), .B(n4600), .Z(n3070) );
  ND2 U439 ( .A(n4263), .B(n4575), .Z(n1788) );
  MUX21L U440 ( .A(n1787), .B(n4575), .S(n4935), .Z(n1789) );
  NR2 U441 ( .A(n4575), .B(n4263), .Z(n1787) );
  ND2 U442 ( .A(n1987), .B(n1986), .Z(n1364) );
  ND2 U443 ( .A(n4295), .B(n4924), .Z(n1986) );
  MUX21L U444 ( .A(n1985), .B(n4623), .S(n4924), .Z(n1987) );
  NR2 U445 ( .A(n4623), .B(n4295), .Z(n1985) );
  EN U446 ( .A(n4892), .B(n4215), .Z(n861) );
  ND2 U447 ( .A(n4625), .B(n4293), .Z(n1964) );
  ND2 U448 ( .A(n4896), .B(n4619), .Z(n2834) );
  ND2 U449 ( .A(n3274), .B(n3273), .Z(n870) );
  EN U450 ( .A(n4565), .B(n4240), .Z(n3274) );
  EO U451 ( .A(n4890), .B(n4240), .Z(n3273) );
  MUX21L U452 ( .A(n2120), .B(n4578), .S(n4280), .Z(n852) );
  ND2 U453 ( .A(n4930), .B(n4578), .Z(n2120) );
  ND2 U454 ( .A(n2509), .B(n2508), .Z(n859) );
  ND2 U455 ( .A(n2505), .B(n4945), .Z(n2508) );
  MUX21L U456 ( .A(n2506), .B(n2507), .S(n4945), .Z(n2509) );
  NR2 U457 ( .A(n4594), .B(n4227), .Z(n2505) );
  NR2 U458 ( .A(n4941), .B(n4223), .Z(n2425) );
  NR2 U459 ( .A(n4627), .B(n4257), .Z(n848) );
  ND2 U460 ( .A(n1827), .B(n1826), .Z(n1332) );
  ND2 U461 ( .A(n4937), .B(n4261), .Z(n1826) );
  EO U462 ( .A(n4565), .B(n4261), .Z(n1827) );
  EO U463 ( .A(n4884), .B(n4626), .Z(n1335) );
  ND2 U464 ( .A(n4949), .B(n4212), .Z(n2623) );
  MUX21L U465 ( .A(n1753), .B(n4574), .S(n4265), .Z(n1331) );
  ND2 U466 ( .A(n4935), .B(n4574), .Z(n1753) );
  ND2 U467 ( .A(n4603), .B(n4244), .Z(n863) );
  ND2 U468 ( .A(n2730), .B(n2729), .Z(n834) );
  ND2 U469 ( .A(n2726), .B(n4894), .Z(n2729) );
  MUX21L U470 ( .A(n2727), .B(n2728), .S(n4894), .Z(n2730) );
  NR2 U471 ( .A(n4604), .B(n4219), .Z(n2726) );
  ND2 U472 ( .A(n2989), .B(n2988), .Z(n839) );
  ND2 U473 ( .A(n4611), .B(n4919), .Z(n2989) );
  ND2 U474 ( .A(n4919), .B(n4270), .Z(n2988) );
  AN2P U475 ( .A(n4637), .B(n4284), .Z(n407) );
  EO U476 ( .A(n4889), .B(n4287), .Z(n1309) );
  ND2 U477 ( .A(n2596), .B(n2595), .Z(n1316) );
  MUX21L U478 ( .A(n2593), .B(n2594), .S(n4948), .Z(n2595) );
  MUX21L U479 ( .A(n2591), .B(n2592), .S(n4606), .Z(n2596) );
  NR2 U480 ( .A(n4611), .B(n4212), .Z(n2593) );
  ND2 U481 ( .A(n3289), .B(n3288), .Z(n1328) );
  EO U482 ( .A(n4890), .B(n4241), .Z(n3289) );
  EO U483 ( .A(n4564), .B(n4241), .Z(n3288) );
  NR2 U484 ( .A(n4914), .B(n4616), .Z(n1323) );
  NR2 U485 ( .A(n4609), .B(n4214), .Z(n2638) );
  NR2 U486 ( .A(n4639), .B(n4300), .Z(n825) );
  EN U487 ( .A(n4891), .B(n4605), .Z(n1318) );
  EO U488 ( .A(n4889), .B(n4249), .Z(n814) );
  ND2 U489 ( .A(n4948), .B(n4632), .Z(n2579) );
  ND2 U490 ( .A(n2083), .B(n2082), .Z(n1305) );
  ND2 U491 ( .A(n4928), .B(n4278), .Z(n2082) );
  EO U492 ( .A(n4562), .B(n4278), .Z(n2083) );
  ND2 U493 ( .A(n4931), .B(n4580), .Z(n2143) );
  ND2 U494 ( .A(n4625), .B(n4294), .Z(n1968) );
  ND2 U495 ( .A(n4923), .B(n4294), .Z(n1969) );
  ND2 U496 ( .A(n2688), .B(n2687), .Z(n810) );
  ND2 U497 ( .A(n4904), .B(n4216), .Z(n2687) );
  EO U498 ( .A(n4563), .B(n4216), .Z(n2688) );
  ND2 U499 ( .A(n3294), .B(n3293), .Z(n819) );
  ND2 U500 ( .A(n4590), .B(n4242), .Z(n3293) );
  EO U501 ( .A(n4890), .B(n4242), .Z(n3294) );
  EN U502 ( .A(n4565), .B(n4230), .Z(n808) );
  MUX21L U503 ( .A(n3151), .B(n4908), .S(n4233), .Z(n1327) );
  ND2 U504 ( .A(n4908), .B(n4583), .Z(n3151) );
  MUX21L U505 ( .A(n2021), .B(n4622), .S(n4297), .Z(n1304) );
  ND2 U506 ( .A(n4926), .B(n4622), .Z(n2021) );
  NR2 U507 ( .A(n4942), .B(n4223), .Z(n2429) );
  AO4 U508 ( .A(n4621), .B(n4297), .C(n4926), .D(n4297), .Z(n1272) );
  NR3 U509 ( .A(n4290), .B(n4933), .C(n4572), .Z(n1267) );
  EO U510 ( .A(n4561), .B(n4214), .Z(n1285) );
  EN U511 ( .A(n4892), .B(n4585), .Z(n1295) );
  EO U512 ( .A(n4563), .B(n4282), .Z(n1276) );
  EO U513 ( .A(n4560), .B(n4256), .Z(n1275) );
  ND2 U514 ( .A(n2705), .B(n4606), .Z(n1286) );
  EN U515 ( .A(n4893), .B(n4217), .Z(n2705) );
  ND2 U516 ( .A(n2085), .B(n2084), .Z(n1273) );
  ND2 U517 ( .A(n4929), .B(n4278), .Z(n2085) );
  ND2 U518 ( .A(n4577), .B(n4278), .Z(n2084) );
  ND2 U519 ( .A(n4607), .B(n4216), .Z(n2689) );
  ND2 U520 ( .A(n4904), .B(n4216), .Z(n2690) );
  OR3 U521 ( .A(n4292), .B(n4922), .C(n4626), .Z(n408) );
  NR2 U522 ( .A(n410), .B(n411), .Z(n409) );
  EO U523 ( .A(n4560), .B(n4218), .Z(n410) );
  EO U524 ( .A(n4893), .B(n4218), .Z(n411) );
  MUX21L U525 ( .A(n2747), .B(n4900), .S(n4243), .Z(n1287) );
  ND2 U526 ( .A(n4900), .B(n4604), .Z(n2747) );
  EN U527 ( .A(n4887), .B(n4270), .Z(n794) );
  EN U528 ( .A(n4888), .B(n4614), .Z(n793) );
  AN2P U529 ( .A(n4632), .B(n4230), .Z(n412) );
  NR2 U530 ( .A(n4905), .B(n4581), .Z(n3072) );
  EN U531 ( .A(n4893), .B(n4595), .Z(n2517) );
  EO U532 ( .A(n4887), .B(n4598), .Z(n1262) );
  ND2 U533 ( .A(n2602), .B(n2601), .Z(n1254) );
  MUX21L U534 ( .A(n2599), .B(n2600), .S(n4948), .Z(n2601) );
  MUX21L U535 ( .A(n2597), .B(n2598), .S(n4611), .Z(n2602) );
  NR2 U536 ( .A(n4611), .B(n4210), .Z(n2599) );
  ND2 U537 ( .A(n2770), .B(n4244), .Z(n1257) );
  EO U538 ( .A(n4886), .B(n4602), .Z(n2770) );
  ND2 U539 ( .A(n3207), .B(n3206), .Z(n1264) );
  MUX21L U540 ( .A(n3205), .B(n4236), .S(n4586), .Z(n3206) );
  AO2 U541 ( .A(n4910), .B(n4236), .C(n4910), .D(n4586), .Z(n3207) );
  NR2 U542 ( .A(n4910), .B(n4236), .Z(n3205) );
  OR2 U543 ( .A(n4635), .B(n4285), .Z(n413) );
  NR3 U544 ( .A(n4247), .B(n4898), .C(n4620), .Z(n774) );
  ND2 U545 ( .A(n4945), .B(n4228), .Z(n2516) );
  ND2 U546 ( .A(n4240), .B(n3262), .Z(n1265) );
  ND2 U547 ( .A(n4912), .B(n4589), .Z(n3262) );
  ND2 U548 ( .A(n4913), .B(n4616), .Z(n2882) );
  IVP U549 ( .A(n1241), .Z(n3849) );
  AO7 U550 ( .A(n4936), .B(n4576), .C(n4263), .Z(n1241) );
  ND2 U551 ( .A(n4904), .B(n4216), .Z(n2692) );
  ND2 U552 ( .A(n4606), .B(n4217), .Z(n2691) );
  ND2 U553 ( .A(n2686), .B(n2685), .Z(n1229) );
  ND2 U554 ( .A(n4904), .B(n4216), .Z(n2685) );
  EN U555 ( .A(n4892), .B(n4607), .Z(n2686) );
  NR3 U556 ( .A(n4222), .B(n4941), .C(n4568), .Z(n1224) );
  NR2 U557 ( .A(n4905), .B(n4252), .Z(n3085) );
  NR2 U558 ( .A(n415), .B(n416), .Z(n414) );
  EN U559 ( .A(n4562), .B(n4231), .Z(n415) );
  AN2P U560 ( .A(n4907), .B(n4231), .Z(n416) );
  ND2 U561 ( .A(n3153), .B(n3152), .Z(n1218) );
  EN U562 ( .A(n4563), .B(n4233), .Z(n3153) );
  EN U563 ( .A(n4893), .B(n4233), .Z(n3152) );
  OR3 U564 ( .A(n4257), .B(n4939), .C(n4628), .Z(n417) );
  ND2 U565 ( .A(n4590), .B(n4242), .Z(n3295) );
  EO U566 ( .A(n4890), .B(n4242), .Z(n3296) );
  ND2 U567 ( .A(n3291), .B(n3290), .Z(n1202) );
  ND2 U568 ( .A(n4590), .B(n4241), .Z(n3290) );
  EO U569 ( .A(n4890), .B(n4241), .Z(n3291) );
  ND2 U570 ( .A(n3155), .B(n3154), .Z(n1201) );
  EN U571 ( .A(n4563), .B(n4233), .Z(n3155) );
  EN U572 ( .A(n4893), .B(n4233), .Z(n3154) );
  NR2 U573 ( .A(n4906), .B(n4253), .Z(n3105) );
  ND3 U574 ( .A(n3060), .B(n3059), .C(n3058), .Z(n1199) );
  ND2 U575 ( .A(n4600), .B(n4922), .Z(n3060) );
  ND2 U576 ( .A(n4922), .B(n4266), .Z(n3059) );
  ND2 U577 ( .A(n4600), .B(n4266), .Z(n3058) );
  NR2 U578 ( .A(n4917), .B(n4273), .Z(n2957) );
  NR2 U579 ( .A(n4584), .B(n4233), .Z(n3157) );
  ND2 U580 ( .A(n2937), .B(n2936), .Z(n1184) );
  EO U581 ( .A(n4888), .B(n4274), .Z(n2937) );
  EO U582 ( .A(n4566), .B(n4274), .Z(n2936) );
  IVP U583 ( .A(n756), .Z(n3859) );
  AO4 U584 ( .A(n4585), .B(n4234), .C(n4909), .D(n4234), .Z(n756) );
  NR2 U585 ( .A(n4606), .B(n4217), .Z(n1181) );
  ND2 U586 ( .A(n2993), .B(n2992), .Z(n1176) );
  ND2 U587 ( .A(n4919), .B(n4270), .Z(n2992) );
  EO U588 ( .A(n4560), .B(n4270), .Z(n2993) );
  EO U589 ( .A(n4561), .B(n4252), .Z(n1178) );
  AO4 U590 ( .A(n4610), .B(n4212), .C(n4948), .D(n4210), .Z(n1173) );
  EN U591 ( .A(n4891), .B(n4237), .Z(n3223) );
  NR2 U592 ( .A(n4582), .B(n4253), .Z(n3109) );
  NR2 U593 ( .A(n4906), .B(n4253), .Z(n3110) );
  ND2 U594 ( .A(n4613), .B(n4274), .Z(n2940) );
  ND2 U595 ( .A(n4916), .B(n4274), .Z(n2941) );
  MUX21H U596 ( .A(n4911), .B(n4587), .S(n4237), .Z(n418) );
  ND2 U597 ( .A(n4907), .B(n4253), .Z(n3113) );
  NR2 U598 ( .A(n4590), .B(n4240), .Z(n3264) );
  ND3 U599 ( .A(n4581), .B(n4252), .C(n4905), .Z(n1160) );
  NR2 U600 ( .A(n4925), .B(n4296), .Z(n1996) );
  NR2 U601 ( .A(n4912), .B(n4239), .Z(n3252) );
  AO4 U602 ( .A(n4612), .B(n4271), .C(n4918), .D(n4271), .Z(n506) );
  ND2 U603 ( .A(n4583), .B(n4232), .Z(n3136) );
  MUX21L U604 ( .A(n1995), .B(n1996), .S(n4623), .Z(n1997) );
  MUX21L U605 ( .A(n1993), .B(n1994), .S(n4925), .Z(n1998) );
  AO4 U606 ( .A(n4637), .B(n4283), .C(n4952), .D(n4283), .Z(n491) );
  NR2 U607 ( .A(n4629), .B(n4259), .Z(n1875) );
  NR2 U608 ( .A(n4926), .B(n4298), .Z(n2030) );
  NR2 U609 ( .A(n4590), .B(n4241), .Z(n3276) );
  NR2 U610 ( .A(n4913), .B(n4241), .Z(n3277) );
  NR2 U611 ( .A(n4921), .B(n4268), .Z(n3026) );
  NR2 U612 ( .A(n4292), .B(n4625), .Z(n1946) );
  NR2 U613 ( .A(n4578), .B(n4280), .Z(n2123) );
  ND2 U614 ( .A(n2016), .B(n2015), .Z(n665) );
  EN U615 ( .A(n4885), .B(n4296), .Z(n2016) );
  EO U616 ( .A(n4561), .B(n4296), .Z(n2015) );
  ND2 U617 ( .A(n4629), .B(n4938), .Z(n1882) );
  ND2 U618 ( .A(n2874), .B(n2873), .Z(n683) );
  ND2 U619 ( .A(n2870), .B(n4617), .Z(n2873) );
  MUX21L U620 ( .A(n2871), .B(n2872), .S(n4894), .Z(n2874) );
  NR2 U621 ( .A(n4893), .B(n4251), .Z(n2870) );
  ND2 U622 ( .A(n2574), .B(n2573), .Z(n646) );
  ND2 U623 ( .A(n4632), .B(n4230), .Z(n2573) );
  EN U624 ( .A(n4891), .B(n4230), .Z(n2574) );
  ND2 U625 ( .A(n2744), .B(n2743), .Z(n649) );
  ND2 U626 ( .A(n4899), .B(n4243), .Z(n2743) );
  EO U627 ( .A(n4561), .B(n4243), .Z(n2744) );
  ND2 U628 ( .A(n2048), .B(n2047), .Z(n636) );
  EN U629 ( .A(n4886), .B(n4299), .Z(n2048) );
  EO U630 ( .A(n4560), .B(n4299), .Z(n2047) );
  ND2 U631 ( .A(n2185), .B(n2184), .Z(n607) );
  EO U632 ( .A(n4888), .B(n4277), .Z(n2185) );
  EO U633 ( .A(n4562), .B(n4277), .Z(n2184) );
  ND2 U634 ( .A(n2630), .B(n2629), .Z(n617) );
  ND2 U635 ( .A(n4609), .B(n4213), .Z(n2629) );
  EN U636 ( .A(n4890), .B(n4212), .Z(n2630) );
  ND2 U637 ( .A(n2515), .B(n2514), .Z(n615) );
  ND2 U638 ( .A(n4227), .B(n4595), .Z(n2514) );
  MUX21L U639 ( .A(n2513), .B(n4595), .S(n4945), .Z(n2515) );
  NR2 U640 ( .A(n4595), .B(n4227), .Z(n2513) );
  ND2 U641 ( .A(n3131), .B(n3130), .Z(n536) );
  EO U642 ( .A(n4893), .B(n4231), .Z(n3131) );
  EO U643 ( .A(n4562), .B(n4231), .Z(n3130) );
  EN U644 ( .A(n4565), .B(n4261), .Z(n693) );
  EN U645 ( .A(n4885), .B(n4625), .Z(n696) );
  ND3 U646 ( .A(n4561), .B(n4207), .C(n4885), .Z(n419) );
  IVP U647 ( .A(n526), .Z(n3855) );
  AO4 U648 ( .A(n4594), .B(n4226), .C(n4945), .D(n4226), .Z(n526) );
  ND2 U649 ( .A(n2180), .B(n2179), .Z(n700) );
  ND2 U650 ( .A(n4254), .B(n4951), .Z(n2179) );
  MUX21L U651 ( .A(n2178), .B(n4567), .S(n4951), .Z(n2180) );
  NR2 U652 ( .A(n4567), .B(n4254), .Z(n2178) );
  ND2 U653 ( .A(n2126), .B(n2125), .Z(n638) );
  MUX21L U654 ( .A(n2121), .B(n2122), .S(n4578), .Z(n2126) );
  MUX21L U655 ( .A(n2123), .B(n2124), .S(n4930), .Z(n2125) );
  NR3 U656 ( .A(n4244), .B(n4904), .C(n4602), .Z(n529) );
  NR3 U657 ( .A(n4222), .B(n4941), .C(n4568), .Z(n673) );
  AO7 U658 ( .A(n4950), .B(n4580), .C(n4255), .Z(n544) );
  AO4 U659 ( .A(n4620), .B(n4247), .C(n4898), .D(n4620), .Z(n742) );
  AO4 U660 ( .A(n4620), .B(n4247), .C(n4897), .D(n4247), .Z(n651) );
  AO4 U661 ( .A(n4579), .B(n4280), .C(n4930), .D(n4280), .Z(n572) );
  NR2 U662 ( .A(n4912), .B(n4588), .Z(n719) );
  NR2 U663 ( .A(n4912), .B(n4589), .Z(n658) );
  NR2 U664 ( .A(n4592), .B(n4224), .Z(n549) );
  NR2 U665 ( .A(n4618), .B(n4249), .Z(n532) );
  AN3 U666 ( .A(n4561), .B(n4208), .C(n4888), .Z(n728) );
  EN U667 ( .A(n4892), .B(n4229), .Z(n706) );
  EO U668 ( .A(n4893), .B(n4257), .Z(n663) );
  EO U669 ( .A(n4891), .B(n4575), .Z(n629) );
  EN U670 ( .A(n4893), .B(n4629), .Z(n631) );
  EO U671 ( .A(n4889), .B(n4283), .Z(n640) );
  EO U672 ( .A(n4563), .B(n4262), .Z(n598) );
  EO U673 ( .A(n4888), .B(n4571), .Z(n611) );
  EO U674 ( .A(n4886), .B(n4568), .Z(n613) );
  EO U675 ( .A(n4886), .B(n4602), .Z(n586) );
  EN U676 ( .A(n4888), .B(n4274), .Z(n590) );
  EO U677 ( .A(n4888), .B(n4620), .Z(n588) );
  EO U678 ( .A(n4564), .B(n4249), .Z(n557) );
  EN U679 ( .A(n4885), .B(n4599), .Z(n560) );
  EN U680 ( .A(n4887), .B(n4611), .Z(n559) );
  ND2 U681 ( .A(n4583), .B(n4232), .Z(n3138) );
  ND2 U682 ( .A(n4907), .B(n4232), .Z(n3139) );
  ND2 U683 ( .A(n4622), .B(n4925), .Z(n2009) );
  ND2 U684 ( .A(n3133), .B(n3132), .Z(n518) );
  ND2 U685 ( .A(n4907), .B(n4232), .Z(n3133) );
  ND2 U686 ( .A(n4583), .B(n4232), .Z(n3132) );
  ND2 U687 ( .A(n4603), .B(n4244), .Z(n680) );
  ND2 U688 ( .A(n2935), .B(n2934), .Z(n622) );
  ND2 U689 ( .A(n4916), .B(n4614), .Z(n2935) );
  ND2 U690 ( .A(n4613), .B(n4274), .Z(n2934) );
  ND2 U691 ( .A(n2187), .B(n2186), .Z(n573) );
  ND2 U692 ( .A(n4639), .B(n4277), .Z(n2186) );
  ND2 U693 ( .A(n4951), .B(n4277), .Z(n2187) );
  ND2 U694 ( .A(n2943), .B(n2942), .Z(n533) );
  ND2 U695 ( .A(n4916), .B(n4274), .Z(n2943) );
  ND2 U696 ( .A(n4613), .B(n4273), .Z(n2942) );
  AN2P U697 ( .A(n4597), .B(n4270), .Z(n420) );
  MUX21L U698 ( .A(n2033), .B(n4641), .S(n4298), .Z(n604) );
  ND2 U699 ( .A(n4926), .B(n4641), .Z(n2033) );
  MUX21L U700 ( .A(n2498), .B(n4594), .S(n4226), .Z(n581) );
  ND2 U701 ( .A(n4944), .B(n4594), .Z(n2498) );
  MUX21L U702 ( .A(n4239), .B(n4912), .S(n4589), .Z(n538) );
  ND2 U703 ( .A(n4639), .B(n4300), .Z(n571) );
  MUX21L U704 ( .A(n4582), .B(n4906), .S(n4252), .Z(n624) );
  IVP U705 ( .A(n4031), .Z(n4211) );
  IVP U706 ( .A(n4033), .Z(n4225) );
  IVP U707 ( .A(n4387), .Z(n4619) );
  IVP U708 ( .A(n4025), .Z(n4284) );
  IVP U709 ( .A(n4025), .Z(n4281) );
  IVP U710 ( .A(n4385), .Z(n4634) );
  IVP U711 ( .A(n4027), .Z(n4273) );
  IVP U712 ( .A(n4396), .Z(n4569) );
  IVP U713 ( .A(n4031), .Z(n4214) );
  IVP U714 ( .A(n4732), .Z(n4891) );
  IVP U715 ( .A(n4033), .Z(n4223) );
  IVP U716 ( .A(n4397), .Z(n4562) );
  IVP U717 ( .A(n4036), .Z(n4241) );
  IVP U718 ( .A(n4730), .Z(n4903) );
  IVP U719 ( .A(n4396), .Z(n4566) );
  IVP U720 ( .A(n4028), .Z(n4264) );
  IVP U721 ( .A(n4024), .Z(n4289) );
  IVP U722 ( .A(n4732), .Z(n4892) );
  IVP U723 ( .A(n4024), .Z(n4290) );
  IVP U724 ( .A(n4722), .Z(n4949) );
  IVP U725 ( .A(n4397), .Z(n4563) );
  IVP U726 ( .A(n4031), .Z(n4213) );
  IVP U727 ( .A(n4730), .Z(n4904) );
  IVP U728 ( .A(n4390), .Z(n4602) );
  IVP U729 ( .A(n4390), .Z(n4560) );
  IVP U730 ( .A(n4024), .Z(n4291) );
  IVP U731 ( .A(n4387), .Z(n4624) );
  IVP U732 ( .A(n4037), .Z(n4250) );
  IVP U733 ( .A(n4032), .Z(n4222) );
  IVP U734 ( .A(n4386), .Z(n4630) );
  IVP U735 ( .A(n4033), .Z(n4228) );
  IVP U736 ( .A(n4723), .Z(n4946) );
  IVP U737 ( .A(n4390), .Z(n4606) );
  IVP U738 ( .A(n4724), .Z(n4941) );
  IVP U739 ( .A(n4392), .Z(n4595) );
  NR2 U740 ( .A(n4630), .B(n4824), .Z(n1853) );
  NR2 U741 ( .A(n4630), .B(n4127), .Z(n1854) );
  NR2 U742 ( .A(n4250), .B(n4748), .Z(n2848) );
  NR2 U743 ( .A(n4250), .B(n4497), .Z(n2849) );
  ND2 U744 ( .A(n1786), .B(n1785), .Z(n1657) );
  ND2 U745 ( .A(n4935), .B(n4120), .Z(n1785) );
  EO U746 ( .A(n4564), .B(n4264), .Z(n1786) );
  ND2 U747 ( .A(n1856), .B(n1855), .Z(n1659) );
  MUX21L U748 ( .A(n1852), .B(n4260), .S(n4938), .Z(n1855) );
  NR2 U749 ( .A(n1854), .B(n1853), .Z(n1856) );
  NR2 U750 ( .A(n4259), .B(n4526), .Z(n1852) );
  ND2 U751 ( .A(n2581), .B(n2580), .Z(n1677) );
  ND2 U752 ( .A(n4060), .B(n4848), .Z(n2580) );
  EN U753 ( .A(n4564), .B(n4213), .Z(n2581) );
  ND2 U754 ( .A(n2417), .B(n2416), .Z(n1673) );
  ND2 U755 ( .A(n4567), .B(n4163), .Z(n2416) );
  EO U756 ( .A(n4886), .B(n4222), .Z(n2417) );
  ND2 U757 ( .A(n2135), .B(n2134), .Z(n1666) );
  ND2 U758 ( .A(n4281), .B(n4798), .Z(n2134) );
  EO U759 ( .A(n4561), .B(n4281), .Z(n2135) );
  ND2 U760 ( .A(n2345), .B(n4868), .Z(n1670) );
  EO U761 ( .A(n4560), .B(n4289), .Z(n2345) );
  ND2 U762 ( .A(n2851), .B(n2850), .Z(n1682) );
  MUX21L U763 ( .A(n2847), .B(n4617), .S(n4894), .Z(n2850) );
  NR2 U764 ( .A(n2849), .B(n2848), .Z(n2851) );
  NR2 U765 ( .A(n4617), .B(n4098), .Z(n2847) );
  ND2 U766 ( .A(n2828), .B(n2827), .Z(n1681) );
  ND2 U767 ( .A(n4248), .B(n4753), .Z(n2827) );
  EO U768 ( .A(n4889), .B(n4619), .Z(n2828) );
  ND2 U769 ( .A(n4214), .B(n4842), .Z(n2647) );
  ND2 U770 ( .A(n1774), .B(n1773), .Z(n1624) );
  ND2 U771 ( .A(n4515), .B(n4831), .Z(n1773) );
  MUX21L U772 ( .A(n4515), .B(n1772), .S(n4264), .Z(n1774) );
  ND2 U773 ( .A(n1701), .B(n1700), .Z(n1623) );
  ND2 U774 ( .A(n4290), .B(n4837), .Z(n1700) );
  EN U775 ( .A(n4564), .B(n4290), .Z(n1701) );
  ND2 U776 ( .A(n1971), .B(n1970), .Z(n1629) );
  ND2 U777 ( .A(n4923), .B(n4202), .Z(n1970) );
  EN U778 ( .A(n4885), .B(n4624), .Z(n1971) );
  ND2 U779 ( .A(n2255), .B(n2254), .Z(n1636) );
  ND2 U780 ( .A(n4636), .B(n4183), .Z(n2254) );
  EN U781 ( .A(n4889), .B(n4284), .Z(n2255) );
  ND2 U782 ( .A(n2351), .B(n2350), .Z(n1638) );
  ND2 U783 ( .A(n4171), .B(n4419), .Z(n2350) );
  EN U784 ( .A(n4888), .B(n4569), .Z(n2351) );
  ND2 U785 ( .A(n2051), .B(n2050), .Z(n1632) );
  ND2 U786 ( .A(n4193), .B(n4805), .Z(n2050) );
  EN U787 ( .A(n4560), .B(n4299), .Z(n2051) );
  ND2 U788 ( .A(n3281), .B(n3280), .Z(n1653) );
  ND2 U789 ( .A(n4913), .B(n4074), .Z(n3280) );
  EO U790 ( .A(n4565), .B(n4241), .Z(n3281) );
  ND2 U791 ( .A(n2853), .B(n2852), .Z(n1647) );
  ND2 U792 ( .A(n4250), .B(n4497), .Z(n2852) );
  EO U793 ( .A(n4889), .B(n4250), .Z(n2853) );
  MUX21L U794 ( .A(n2519), .B(n4853), .S(n4228), .Z(n2521) );
  ND2 U795 ( .A(n2303), .B(n2302), .Z(n1128) );
  ND2 U796 ( .A(n4634), .B(n4287), .Z(n2302) );
  MUX21L U797 ( .A(n2301), .B(n4872), .S(n4287), .Z(n2303) );
  NR2 U798 ( .A(n4634), .B(n4872), .Z(n2301) );
  IVP U799 ( .A(n4730), .Z(n4901) );
  IVP U800 ( .A(n4028), .Z(n4266) );
  IVP U801 ( .A(n4037), .Z(n4248) );
  IVP U802 ( .A(n4035), .Z(n4236) );
  IVP U803 ( .A(n4029), .Z(n4258) );
  IVP U804 ( .A(n4395), .Z(n4573) );
  IVP U805 ( .A(n4724), .Z(n4936) );
  IVP U806 ( .A(n4386), .Z(n4628) );
  IVP U807 ( .A(n4391), .Z(n4596) );
  IVP U808 ( .A(n4032), .Z(n4220) );
  IVP U809 ( .A(n4384), .Z(n4640) );
  IVP U810 ( .A(n4029), .Z(n4259) );
  IVP U811 ( .A(n4027), .Z(n4271) );
  IVP U812 ( .A(n4729), .Z(n4908) );
  IVP U813 ( .A(n4730), .Z(n4902) );
  IVP U814 ( .A(n4392), .Z(n4590) );
  IVP U815 ( .A(n4036), .Z(n4240) );
  IVP U816 ( .A(n4386), .Z(n4626) );
  IVP U817 ( .A(n4387), .Z(n4621) );
  IVP U818 ( .A(n4028), .Z(n4265) );
  IVP U819 ( .A(n4390), .Z(n4604) );
  IVP U820 ( .A(n4032), .Z(n4217) );
  IVP U821 ( .A(n4392), .Z(n4593) );
  IVP U822 ( .A(n4037), .Z(n4247) );
  IVP U823 ( .A(n4388), .Z(n4615) );
  IVP U824 ( .A(n4732), .Z(n4890) );
  IVP U825 ( .A(n4729), .Z(n4907) );
  IVP U826 ( .A(n4038), .Z(n4254) );
  IVP U827 ( .A(n4384), .Z(n4637) );
  IVP U828 ( .A(n4034), .Z(n4232) );
  IVP U829 ( .A(n4732), .Z(n4889) );
  IVP U830 ( .A(n4030), .Z(n4209) );
  IVP U831 ( .A(n4722), .Z(n4951) );
  IVP U832 ( .A(n4396), .Z(n4567) );
  IVP U833 ( .A(n4733), .Z(n4885) );
  IVP U834 ( .A(n4024), .Z(n4288) );
  IVP U835 ( .A(n4030), .Z(n4208) );
  IVP U836 ( .A(n4733), .Z(n4888) );
  IVP U837 ( .A(n4030), .Z(n4210) );
  IVP U838 ( .A(n4384), .Z(n4639) );
  IVP U839 ( .A(n4395), .Z(n4575) );
  IVP U840 ( .A(n4396), .Z(n4568) );
  IVP U841 ( .A(n4385), .Z(n4633) );
  IVP U842 ( .A(n4728), .Z(n4915) );
  IVP U843 ( .A(n4389), .Z(n4608) );
  IVP U844 ( .A(n4390), .Z(n4603) );
  IVP U845 ( .A(n4728), .Z(n4913) );
  IVP U846 ( .A(n4391), .Z(n4599) );
  IVP U847 ( .A(n4034), .Z(n4231) );
  IVP U848 ( .A(n4397), .Z(n4561) );
  IVP U849 ( .A(n4032), .Z(n4219) );
  IVP U850 ( .A(n4036), .Z(n4243) );
  IVP U851 ( .A(n4392), .Z(n4592) );
  IVP U852 ( .A(n4725), .Z(n4930) );
  IVP U853 ( .A(n4394), .Z(n4580) );
  IVP U854 ( .A(n4722), .Z(n4950) );
  IVP U855 ( .A(n4024), .Z(n4287) );
  IVP U856 ( .A(n4388), .Z(n4614) );
  IVP U857 ( .A(n4724), .Z(n4938) );
  IVP U858 ( .A(n4029), .Z(n4260) );
  IVP U859 ( .A(n4394), .Z(n4579) );
  IVP U860 ( .A(n4393), .Z(n4586) );
  IVP U861 ( .A(n4034), .Z(n4229) );
  IVP U862 ( .A(n4397), .Z(n4564) );
  IVP U863 ( .A(n4028), .Z(n4267) );
  IVP U864 ( .A(n4727), .Z(n4921) );
  IVP U865 ( .A(n4027), .Z(n4272) );
  IVP U866 ( .A(n4025), .Z(n4283) );
  IVP U867 ( .A(n4386), .Z(n4627) );
  IVP U868 ( .A(n4036), .Z(n4242) );
  IVP U869 ( .A(n4727), .Z(n4922) );
  IVP U870 ( .A(n4727), .Z(n4884) );
  IVP U871 ( .A(n4032), .Z(n4221) );
  IVP U872 ( .A(n4029), .Z(n4263) );
  IVP U873 ( .A(n4395), .Z(n4576) );
  IVP U874 ( .A(n4391), .Z(n4600) );
  IVP U875 ( .A(n4036), .Z(n4244) );
  IVP U876 ( .A(n4395), .Z(n4577) );
  IVP U877 ( .A(n4726), .Z(n4929) );
  IVP U878 ( .A(n4036), .Z(n4245) );
  IVP U879 ( .A(n4389), .Z(n4611) );
  IVP U880 ( .A(n4394), .Z(n4583) );
  IVP U881 ( .A(n4387), .Z(n4623) );
  IVP U882 ( .A(n4023), .Z(n4298) );
  IVP U883 ( .A(n4035), .Z(n4239) );
  IVP U884 ( .A(n4023), .Z(n4297) );
  IVP U885 ( .A(n4385), .Z(n4636) );
  IVP U886 ( .A(n4722), .Z(n4953) );
  IVP U887 ( .A(n4732), .Z(n4893) );
  IVP U888 ( .A(n4727), .Z(n4923) );
  IVP U889 ( .A(n4034), .Z(n4255) );
  IVP U890 ( .A(n4397), .Z(n4565) );
  IVP U891 ( .A(n4031), .Z(n4215) );
  IVP U892 ( .A(n4029), .Z(n4262) );
  IVP U893 ( .A(n4732), .Z(n4894) );
  IVP U894 ( .A(n4388), .Z(n4617) );
  IVP U895 ( .A(n4394), .Z(n4582) );
  IVP U896 ( .A(n4725), .Z(n4935) );
  IVP U897 ( .A(n4722), .Z(n4952) );
  IVP U898 ( .A(n4027), .Z(n4275) );
  IVP U899 ( .A(n4728), .Z(n4918) );
  IVP U900 ( .A(n4724), .Z(n4940) );
  IVP U901 ( .A(n4392), .Z(n4594) );
  IVP U902 ( .A(n4393), .Z(n4589) );
  AO7 U903 ( .A(n4938), .B(n4130), .C(n1886), .Z(n1085) );
  ND2 U904 ( .A(n4628), .B(n4258), .Z(n1886) );
  AO7 U905 ( .A(n4934), .B(n4115), .C(n1741), .Z(n1082) );
  ND2 U906 ( .A(n4573), .B(n4289), .Z(n1741) );
  AO7 U907 ( .A(n4571), .B(n4169), .C(n2373), .Z(n1097) );
  ND2 U908 ( .A(n4958), .B(n4220), .Z(n2373) );
  AO7 U909 ( .A(n4280), .B(n4800), .C(n2129), .Z(n1633) );
  ND2 U910 ( .A(n4930), .B(n4579), .Z(n2129) );
  AO7 U911 ( .A(n4896), .B(n4494), .C(n2829), .Z(n1646) );
  ND2 U912 ( .A(n4619), .B(n4248), .Z(n2829) );
  AO7 U913 ( .A(n4271), .B(n4735), .C(n2975), .Z(n1649) );
  ND2 U914 ( .A(n4918), .B(n4611), .Z(n2975) );
  NR2 U915 ( .A(n4283), .B(n4549), .Z(n2220) );
  NR2 U916 ( .A(n4637), .B(n4879), .Z(n2221) );
  NR2 U917 ( .A(n4575), .B(n4120), .Z(n1777) );
  NR2 U918 ( .A(n4936), .B(n4430), .Z(n1805) );
  NR2 U919 ( .A(n4936), .B(n4533), .Z(n1927) );
  ND2 U920 ( .A(n4929), .B(n4577), .Z(n2092) );
  ND3 U921 ( .A(n2780), .B(n2779), .C(n2778), .Z(n1679) );
  ND2 U922 ( .A(n4245), .B(n4756), .Z(n2779) );
  ND2 U923 ( .A(n4602), .B(n4756), .Z(n2780) );
  ND2 U924 ( .A(n4602), .B(n4245), .Z(n2778) );
  ND3 U925 ( .A(n2646), .B(n2645), .C(n2644), .Z(n1678) );
  ND2 U926 ( .A(n4054), .B(n4843), .Z(n2645) );
  ND2 U927 ( .A(n4608), .B(n4843), .Z(n2646) );
  ND2 U928 ( .A(n4608), .B(n4054), .Z(n2644) );
  ND2 U929 ( .A(n2224), .B(n2223), .Z(n1668) );
  NR2 U930 ( .A(n2222), .B(n2221), .Z(n2224) );
  MUX21L U931 ( .A(n2220), .B(n4283), .S(n4952), .Z(n2223) );
  NR2 U932 ( .A(n4637), .B(n4187), .Z(n2222) );
  ND2 U933 ( .A(n3050), .B(n3049), .Z(n1685) );
  ND2 U934 ( .A(n4266), .B(n4600), .Z(n3049) );
  MUX21L U935 ( .A(n3048), .B(n4771), .S(n4600), .Z(n3050) );
  NR2 U936 ( .A(n4266), .B(n4771), .Z(n3048) );
  ND2 U937 ( .A(n3142), .B(n3141), .Z(n1687) );
  ND2 U938 ( .A(n4232), .B(n4444), .Z(n3141) );
  MUX21L U939 ( .A(n4907), .B(n3140), .S(n4583), .Z(n3142) );
  NR2 U940 ( .A(n4908), .B(n4232), .Z(n3140) );
  ND2 U941 ( .A(n2751), .B(n2750), .Z(n1139) );
  MUX21L U942 ( .A(n2748), .B(n4757), .S(n4603), .Z(n2750) );
  AO6 U943 ( .A(n4603), .B(n4043), .C(n2749), .Z(n2751) );
  ND2 U944 ( .A(n2420), .B(n4162), .Z(n1132) );
  EN U945 ( .A(n4886), .B(n4566), .Z(n2420) );
  ND2 U946 ( .A(n2465), .B(n2464), .Z(n1133) );
  ND2 U947 ( .A(n4225), .B(n4857), .Z(n2464) );
  EO U948 ( .A(n4885), .B(n4592), .Z(n2465) );
  ND2 U949 ( .A(n2675), .B(n2674), .Z(n1137) );
  ND2 U950 ( .A(n4215), .B(n4476), .Z(n2674) );
  MUX21L U951 ( .A(n2673), .B(n4901), .S(n4215), .Z(n2675) );
  NR2 U952 ( .A(n4902), .B(n4476), .Z(n2673) );
  ND2 U953 ( .A(n2558), .B(n2557), .Z(n1135) );
  ND2 U954 ( .A(n4462), .B(n4850), .Z(n2557) );
  MUX21L U955 ( .A(n4463), .B(n2556), .S(n4229), .Z(n2558) );
  ND2 U956 ( .A(n2962), .B(n2961), .Z(n1144) );
  ND2 U957 ( .A(n4272), .B(n4737), .Z(n2961) );
  MUX21L U958 ( .A(n4509), .B(n2960), .S(n4917), .Z(n2962) );
  NR2 U959 ( .A(n4272), .B(n4509), .Z(n2960) );
  ND2 U960 ( .A(n3047), .B(n3046), .Z(n1145) );
  ND2 U961 ( .A(n4267), .B(n4452), .Z(n3046) );
  EO U962 ( .A(n4886), .B(n4266), .Z(n3047) );
  ND2 U963 ( .A(n2826), .B(n2825), .Z(n1141) );
  ND2 U964 ( .A(n4248), .B(n4494), .Z(n2825) );
  EO U965 ( .A(n4889), .B(n4248), .Z(n2826) );
  ND2 U966 ( .A(n3269), .B(n3268), .Z(n1148) );
  ND2 U967 ( .A(n4074), .B(n4431), .Z(n3268) );
  EO U968 ( .A(n4890), .B(n4590), .Z(n3269) );
  ND2 U969 ( .A(n1697), .B(n1696), .Z(n1116) );
  ND2 U970 ( .A(n4107), .B(n4523), .Z(n1696) );
  EN U971 ( .A(n4890), .B(n4291), .Z(n1697) );
  ND2 U972 ( .A(n1807), .B(n1806), .Z(n1119) );
  ND2 U973 ( .A(n1803), .B(n4829), .Z(n1806) );
  MUX21L U974 ( .A(n1804), .B(n1805), .S(n4263), .Z(n1807) );
  NR2 U975 ( .A(n4263), .B(n4576), .Z(n1803) );
  ND2 U976 ( .A(n1755), .B(n1754), .Z(n1083) );
  ND2 U977 ( .A(n4574), .B(n4118), .Z(n1754) );
  EN U978 ( .A(n4891), .B(n4265), .Z(n1755) );
  ND2 U979 ( .A(n2537), .B(n2536), .Z(n1102) );
  ND2 U980 ( .A(n4596), .B(n4063), .Z(n2536) );
  MUX21L U981 ( .A(n2535), .B(n4063), .S(n4947), .Z(n2537) );
  NR2 U982 ( .A(n4596), .B(n4062), .Z(n2535) );
  ND2 U983 ( .A(n3055), .B(n3054), .Z(n1111) );
  ND2 U984 ( .A(n4266), .B(n4772), .Z(n3054) );
  EO U985 ( .A(n4561), .B(n4266), .Z(n3055) );
  ND2 U986 ( .A(n3292), .B(n4796), .Z(n1114) );
  EO U987 ( .A(n4564), .B(n4242), .Z(n3292) );
  ND2 U988 ( .A(n2982), .B(n2981), .Z(n1110) );
  ND2 U989 ( .A(n4271), .B(n4488), .Z(n2981) );
  MUX21L U990 ( .A(n2980), .B(n4918), .S(n4271), .Z(n2982) );
  NR2 U991 ( .A(n4918), .B(n4512), .Z(n2980) );
  ND2 U992 ( .A(n2034), .B(n4807), .Z(n1090) );
  EN U993 ( .A(n4560), .B(n4298), .Z(n2034) );
  ND2 U994 ( .A(n2311), .B(n2310), .Z(n1096) );
  ND3 U995 ( .A(n4634), .B(n4178), .C(n4955), .Z(n2310) );
  MUX21L U996 ( .A(n2308), .B(n2309), .S(n4634), .Z(n2311) );
  NR2 U997 ( .A(n4955), .B(n4178), .Z(n2309) );
  ND2 U998 ( .A(n3063), .B(n3062), .Z(n1651) );
  ND2 U999 ( .A(n4600), .B(n4095), .Z(n3062) );
  MUX21L U1000 ( .A(n3061), .B(n4095), .S(n4918), .Z(n3063) );
  NR2 U1001 ( .A(n4600), .B(n4095), .Z(n3061) );
  ND2 U1002 ( .A(n3202), .B(n4788), .Z(n1652) );
  ND2 U1003 ( .A(n4586), .B(n4236), .Z(n3202) );
  ND2 U1004 ( .A(n2472), .B(n2471), .Z(n1609) );
  ND2 U1005 ( .A(n4071), .B(n4404), .Z(n2471) );
  EN U1006 ( .A(n4885), .B(n4225), .Z(n2472) );
  ND2 U1007 ( .A(n2377), .B(n4866), .Z(n1606) );
  EO U1008 ( .A(n4564), .B(n4221), .Z(n2377) );
  ND2 U1009 ( .A(n2098), .B(n2097), .Z(n1601) );
  MUX21L U1010 ( .A(n2095), .B(n2096), .S(n4929), .Z(n2097) );
  MUX21L U1011 ( .A(n2093), .B(n2094), .S(n4577), .Z(n2098) );
  NR2 U1012 ( .A(n4279), .B(n4428), .Z(n2096) );
  AN3 U1013 ( .A(n4478), .B(n4764), .C(n4217), .Z(n421) );
  MUX21L U1014 ( .A(n1925), .B(n1924), .S(n4627), .Z(n1661) );
  ND2 U1015 ( .A(n4940), .B(n4205), .Z(n1925) );
  ND2 U1016 ( .A(n4291), .B(n4816), .Z(n1924) );
  MUX21L U1017 ( .A(n4524), .B(n4932), .S(n4291), .Z(n1655) );
  MUX21L U1018 ( .A(n1819), .B(n4123), .S(n4577), .Z(n1658) );
  ND2 U1019 ( .A(n4123), .B(n4827), .Z(n1819) );
  MUX21L U1020 ( .A(n4957), .B(n4569), .S(n4219), .Z(n1671) );
  MUX21L U1021 ( .A(n4927), .B(n4544), .S(n4298), .Z(n1664) );
  MUX21L U1022 ( .A(n4552), .B(n4284), .S(n4953), .Z(n1669) );
  MUX21L U1023 ( .A(n2916), .B(n2915), .S(n4915), .Z(n1683) );
  ND2 U1024 ( .A(n4615), .B(n4144), .Z(n2916) );
  ND2 U1025 ( .A(n4615), .B(n4275), .Z(n2915) );
  MUX21L U1026 ( .A(n4570), .B(n4957), .S(n4220), .Z(n1130) );
  MUX21L U1027 ( .A(n2189), .B(n2188), .S(n4639), .Z(n1635) );
  ND2 U1028 ( .A(n4951), .B(n4281), .Z(n2189) );
  ND2 U1029 ( .A(n4281), .B(n4882), .Z(n2188) );
  MUX21L U1030 ( .A(n2166), .B(n2165), .S(n4580), .Z(n1634) );
  ND2 U1031 ( .A(n4950), .B(n4139), .Z(n2166) );
  ND2 U1032 ( .A(n4950), .B(n4255), .Z(n2165) );
  MUX21L U1033 ( .A(n4867), .B(n4172), .S(n4568), .Z(n1637) );
  MUX21L U1034 ( .A(n3038), .B(n3037), .S(n4921), .Z(n1650) );
  ND2 U1035 ( .A(n4156), .B(n4453), .Z(n3038) );
  ND2 U1036 ( .A(n4599), .B(n4267), .Z(n3037) );
  MUX21L U1037 ( .A(n2918), .B(n2917), .S(n4915), .Z(n1648) );
  ND2 U1038 ( .A(n4275), .B(n4505), .Z(n2918) );
  ND2 U1039 ( .A(n4614), .B(n4275), .Z(n2917) );
  IVP U1040 ( .A(n4027), .Z(n4270) );
  IVP U1041 ( .A(n4726), .Z(n4927) );
  IVP U1042 ( .A(n4723), .Z(n4943) );
  IVP U1043 ( .A(n4037), .Z(n4246) );
  IVP U1044 ( .A(n4727), .Z(n4919) );
  IVP U1045 ( .A(n4026), .Z(n4279) );
  IVP U1046 ( .A(n4385), .Z(n4631) );
  IVP U1047 ( .A(n4025), .Z(n4282) );
  IVP U1048 ( .A(n4395), .Z(n4574) );
  IVP U1049 ( .A(n4385), .Z(n4632) );
  IVP U1050 ( .A(n4026), .Z(n4278) );
  IVP U1051 ( .A(n4726), .Z(n4924) );
  IVP U1052 ( .A(n4731), .Z(n4896) );
  IVP U1053 ( .A(n4023), .Z(n4294) );
  IVP U1054 ( .A(n4035), .Z(n4234) );
  IVP U1055 ( .A(n4030), .Z(n4256) );
  IVP U1056 ( .A(n4728), .Z(n4914) );
  IVP U1057 ( .A(n4723), .Z(n4944) );
  IVP U1058 ( .A(n4393), .Z(n4587) );
  IVP U1059 ( .A(n4026), .Z(n4276) );
  IVP U1060 ( .A(n4726), .Z(n4926) );
  IVP U1061 ( .A(n4733), .Z(n4886) );
  IVP U1062 ( .A(n4386), .Z(n4625) );
  IVP U1063 ( .A(n4733), .Z(n4887) );
  IVP U1064 ( .A(n4391), .Z(n4597) );
  IVP U1065 ( .A(n4384), .Z(n4638) );
  IVP U1066 ( .A(n4723), .Z(n4942) );
  IVP U1067 ( .A(n4023), .Z(n4293) );
  IVP U1068 ( .A(n4724), .Z(n4937) );
  IVP U1069 ( .A(n4389), .Z(n4607) );
  IVP U1070 ( .A(n4389), .Z(n4610) );
  IVP U1071 ( .A(n4726), .Z(n4925) );
  IVP U1072 ( .A(n4394), .Z(n4578) );
  IVP U1073 ( .A(n4022), .Z(n4299) );
  IVP U1074 ( .A(n4722), .Z(n4948) );
  IVP U1075 ( .A(n4031), .Z(n4212) );
  IVP U1076 ( .A(n4033), .Z(n4224) );
  IVP U1077 ( .A(n4731), .Z(n4898) );
  IVP U1078 ( .A(n4725), .Z(n4931) );
  IVP U1079 ( .A(n4725), .Z(n4932) );
  IVP U1080 ( .A(n4391), .Z(n4601) );
  IVP U1081 ( .A(n4725), .Z(n4934) );
  IVP U1082 ( .A(n4396), .Z(n4570) );
  IVP U1083 ( .A(n4726), .Z(n4928) );
  IVP U1084 ( .A(n4723), .Z(n4947) );
  IVP U1085 ( .A(n4025), .Z(n4285) );
  IVP U1086 ( .A(n4031), .Z(n4216) );
  IVP U1087 ( .A(n4728), .Z(n4917) );
  IVP U1088 ( .A(n4026), .Z(n4280) );
  IVP U1089 ( .A(n4028), .Z(n4269) );
  IVP U1090 ( .A(n4035), .Z(n4238) );
  IVP U1091 ( .A(n4384), .Z(n4641) );
  IVP U1092 ( .A(n4025), .Z(n4286) );
  IVP U1093 ( .A(n4033), .Z(n4227) );
  IVP U1094 ( .A(n4731), .Z(n4900) );
  IVP U1095 ( .A(n4024), .Z(n4292) );
  IVP U1096 ( .A(n4037), .Z(n4251) );
  IVP U1097 ( .A(n4396), .Z(n4571) );
  AO7 U1098 ( .A(n4931), .B(n4424), .C(n4256), .Z(n1667) );
  AO7 U1099 ( .A(n4922), .B(n4533), .C(n4292), .Z(n1122) );
  AO7 U1100 ( .A(n4579), .B(n4189), .C(n2130), .Z(n1092) );
  ND2 U1101 ( .A(n4930), .B(n4280), .Z(n2130) );
  AO7 U1102 ( .A(n4927), .B(n4641), .C(n4194), .Z(n1631) );
  AO7 U1103 ( .A(n4633), .B(n4174), .C(n2330), .Z(n1605) );
  ND2 U1104 ( .A(n4956), .B(n4288), .Z(n2330) );
  AO7 U1105 ( .A(n4259), .B(n4527), .C(n1857), .Z(n1594) );
  ND2 U1106 ( .A(n4938), .B(n4630), .Z(n1857) );
  NR2 U1107 ( .A(n4948), .B(n4059), .Z(n2583) );
  NR2 U1108 ( .A(n4212), .B(n4466), .Z(n2585) );
  NR2 U1109 ( .A(n4929), .B(n4191), .Z(n2094) );
  NR2 U1110 ( .A(n4291), .B(n4523), .Z(n1590) );
  NR2 U1111 ( .A(n4956), .B(n4288), .Z(n2335) );
  ND3 U1112 ( .A(n2273), .B(n2272), .C(n2271), .Z(n1604) );
  ND2 U1113 ( .A(n4953), .B(n4555), .Z(n2272) );
  ND2 U1114 ( .A(n4286), .B(n4953), .Z(n2273) );
  ND2 U1115 ( .A(n4286), .B(n4555), .Z(n2271) );
  ND2 U1116 ( .A(n1747), .B(n4115), .Z(n1117) );
  ND2 U1117 ( .A(n4934), .B(n4573), .Z(n1747) );
  ND2 U1118 ( .A(n3166), .B(n3165), .Z(n1113) );
  ND2 U1119 ( .A(n4442), .B(n4782), .Z(n3166) );
  ND2 U1120 ( .A(n4234), .B(n4782), .Z(n3165) );
  ND2 U1121 ( .A(n4619), .B(n4099), .Z(n2836) );
  ND2 U1122 ( .A(n2054), .B(n2053), .Z(n1600) );
  ND2 U1123 ( .A(n4640), .B(n4804), .Z(n2053) );
  MUX21L U1124 ( .A(n4804), .B(n2052), .S(n4299), .Z(n2054) );
  NR2 U1125 ( .A(n4640), .B(n4804), .Z(n2052) );
  ND2 U1126 ( .A(n4255), .B(n4883), .Z(n1602) );
  ND2 U1127 ( .A(n2363), .B(n2362), .Z(n1068) );
  ND2 U1128 ( .A(n2359), .B(n4957), .Z(n2362) );
  MUX21L U1129 ( .A(n2360), .B(n2361), .S(n4220), .Z(n2363) );
  NR2 U1130 ( .A(n4570), .B(n4220), .Z(n2359) );
  ND2 U1131 ( .A(n2339), .B(n2338), .Z(n1067) );
  MUX21L U1132 ( .A(n2336), .B(n2337), .S(n4956), .Z(n2339) );
  ND2 U1133 ( .A(n2335), .B(n4632), .Z(n2338) );
  NR2 U1134 ( .A(n4632), .B(n4174), .Z(n2336) );
  ND2 U1135 ( .A(n2119), .B(n2118), .Z(n1063) );
  ND2 U1136 ( .A(n2115), .B(n4801), .Z(n2118) );
  MUX21L U1137 ( .A(n2116), .B(n2117), .S(n4578), .Z(n2119) );
  NR2 U1138 ( .A(n4279), .B(n4578), .Z(n2115) );
  ND2 U1139 ( .A(n2150), .B(n2149), .Z(n1064) );
  MUX21L U1140 ( .A(n2147), .B(n2148), .S(n4926), .Z(n2149) );
  MUX21L U1141 ( .A(n2145), .B(n2146), .S(n4580), .Z(n2150) );
  NR2 U1142 ( .A(n4256), .B(n4423), .Z(n2148) );
  ND2 U1143 ( .A(n1955), .B(n1954), .Z(n1058) );
  ND2 U1144 ( .A(n4293), .B(n4815), .Z(n1954) );
  EO U1145 ( .A(n4563), .B(n4293), .Z(n1955) );
  ND2 U1146 ( .A(n3231), .B(n3230), .Z(n1080) );
  ND2 U1147 ( .A(n4911), .B(n4436), .Z(n3230) );
  MUX21L U1148 ( .A(n4436), .B(n3229), .S(n4238), .Z(n3231) );
  NR2 U1149 ( .A(n4911), .B(n4435), .Z(n3229) );
  MUX21L U1150 ( .A(n2606), .B(n2605), .S(n4610), .Z(n1136) );
  ND2 U1151 ( .A(n4210), .B(n4846), .Z(n2605) );
  ND2 U1152 ( .A(n4948), .B(n4211), .Z(n2606) );
  MUX21L U1153 ( .A(n2904), .B(n2903), .S(n4276), .Z(n1143) );
  ND2 U1154 ( .A(n4914), .B(n4615), .Z(n2904) );
  ND2 U1155 ( .A(n4615), .B(n4742), .Z(n2903) );
  MUX21L U1156 ( .A(n3197), .B(n4082), .S(n4586), .Z(n1147) );
  ND2 U1157 ( .A(n4082), .B(n4787), .Z(n3197) );
  MUX21L U1158 ( .A(n2863), .B(n4498), .S(n4893), .Z(n1142) );
  ND2 U1159 ( .A(n4097), .B(n4499), .Z(n2863) );
  MUX21L U1160 ( .A(n1836), .B(n1835), .S(n4630), .Z(n1120) );
  ND2 U1161 ( .A(n4125), .B(n4826), .Z(n1836) );
  ND2 U1162 ( .A(n4260), .B(n4825), .Z(n1835) );
  MUX21L U1163 ( .A(n1978), .B(n1977), .S(n4294), .Z(n1088) );
  ND2 U1164 ( .A(n4624), .B(n4811), .Z(n1977) );
  ND2 U1165 ( .A(n4924), .B(n4624), .Z(n1978) );
  MUX21L U1166 ( .A(n4760), .B(n4484), .S(n4242), .Z(n1104) );
  MUX21L U1167 ( .A(n4212), .B(n2607), .S(n4948), .Z(n1103) );
  ND2 U1168 ( .A(n4211), .B(n4468), .Z(n2607) );
  MUX21L U1169 ( .A(n2196), .B(n2195), .S(n4638), .Z(n1094) );
  ND2 U1170 ( .A(n4951), .B(n4282), .Z(n2196) );
  ND2 U1171 ( .A(n4282), .B(n4880), .Z(n2195) );
  MUX21L U1172 ( .A(n4545), .B(n4300), .S(n4928), .Z(n1091) );
  MUX21L U1173 ( .A(n2996), .B(n2995), .S(n4270), .Z(n1617) );
  ND2 U1174 ( .A(n4459), .B(n4766), .Z(n2995) );
  ND2 U1175 ( .A(n4919), .B(n4597), .Z(n2996) );
  MUX21L U1176 ( .A(n4739), .B(n2946), .S(n4273), .Z(n1616) );
  ND2 U1177 ( .A(n4506), .B(n4739), .Z(n2946) );
  MUX21L U1178 ( .A(n4429), .B(n4828), .S(n4262), .Z(n1593) );
  MUX21L U1179 ( .A(n4541), .B(n4198), .S(n4925), .Z(n1597) );
  MUX21L U1180 ( .A(n4625), .B(n4203), .S(n4923), .Z(n1596) );
  MUX21L U1181 ( .A(n2559), .B(n4947), .S(n4229), .Z(n2561) );
  NR2 U1182 ( .A(n4947), .B(n4462), .Z(n2559) );
  IVP U1183 ( .A(n4023), .Z(n4295) );
  IVP U1184 ( .A(n4724), .Z(n4939) );
  IVP U1185 ( .A(n4391), .Z(n4598) );
  IVP U1186 ( .A(n4727), .Z(n4920) );
  IVP U1187 ( .A(n4394), .Z(n4581) );
  IVP U1188 ( .A(n4729), .Z(n4910) );
  IVP U1189 ( .A(n4725), .Z(n4933) );
  IVP U1190 ( .A(n4395), .Z(n4572) );
  IVP U1191 ( .A(n4728), .Z(n4916) );
  IVP U1192 ( .A(n4386), .Z(n4629) );
  IVP U1193 ( .A(n4729), .Z(n4911) );
  IVP U1194 ( .A(n4028), .Z(n4268) );
  NR2 U1195 ( .A(n4957), .B(n4570), .Z(n2361) );
  NR2 U1196 ( .A(n4930), .B(n4190), .Z(n2117) );
  NR2 U1197 ( .A(n4949), .B(n4137), .Z(n2146) );
  NR2 U1198 ( .A(n4920), .B(n4456), .Z(n3008) );
  NR2 U1199 ( .A(n4234), .B(n4783), .Z(n1079) );
  NR2 U1200 ( .A(n4581), .B(n4093), .Z(n1078) );
  ND2 U1201 ( .A(n4131), .B(n4822), .Z(n1893) );
  ND2 U1202 ( .A(n4131), .B(n4528), .Z(n1894) );
  ND2 U1203 ( .A(n4529), .B(n4822), .Z(n1895) );
  ND2 U1204 ( .A(n4256), .B(n4819), .Z(n1121) );
  ND2 U1205 ( .A(n2924), .B(n2923), .Z(n1583) );
  MUX21L U1206 ( .A(n2921), .B(n2922), .S(n4614), .Z(n2923) );
  MUX21L U1207 ( .A(n2919), .B(n2920), .S(n4915), .Z(n2924) );
  NR2 U1208 ( .A(n4275), .B(n4741), .Z(n2921) );
  ND2 U1209 ( .A(n3044), .B(n3043), .Z(n1585) );
  MUX21L U1210 ( .A(n3041), .B(n3042), .S(n4599), .Z(n3043) );
  MUX21L U1211 ( .A(n3039), .B(n3040), .S(n4921), .Z(n3044) );
  NR2 U1212 ( .A(n4267), .B(n4770), .Z(n3041) );
  ND2 U1213 ( .A(n4135), .B(n4818), .Z(n1920) );
  ND2 U1214 ( .A(n4927), .B(n4544), .Z(n1599) );
  ND2 U1215 ( .A(n2198), .B(n2197), .Z(n1065) );
  ND2 U1216 ( .A(n4951), .B(n4188), .Z(n2197) );
  EN U1217 ( .A(n4889), .B(n4638), .Z(n2198) );
  AN3 U1218 ( .A(n4143), .B(n4741), .C(n4615), .Z(n422) );
  MUX21L U1219 ( .A(n1715), .B(n1714), .S(n4572), .Z(n1053) );
  ND2 U1220 ( .A(n4933), .B(n4290), .Z(n1715) );
  ND2 U1221 ( .A(n4290), .B(n4837), .Z(n1714) );
  MUX21L U1222 ( .A(n1756), .B(n4574), .S(n4265), .Z(n1054) );
  ND2 U1223 ( .A(n4574), .B(n4832), .Z(n1756) );
  MUX21L U1224 ( .A(n1699), .B(n1698), .S(n4932), .Z(n1052) );
  ND2 U1225 ( .A(n4108), .B(n4522), .Z(n1699) );
  ND2 U1226 ( .A(n4621), .B(n4108), .Z(n1698) );
  MUX21L U1227 ( .A(n2864), .B(n4746), .S(n4617), .Z(n1075) );
  ND2 U1228 ( .A(n4250), .B(n4746), .Z(n2864) );
  IVP U1229 ( .A(n4388), .Z(n4613) );
  IVP U1230 ( .A(n4393), .Z(n4584) );
  IVP U1231 ( .A(n4032), .Z(n4218) );
  IVP U1232 ( .A(n4022), .Z(n4300) );
  IVP U1233 ( .A(n4731), .Z(n4895) );
  IVP U1234 ( .A(n4035), .Z(n4235) );
  NR2 U1235 ( .A(n4614), .B(n4145), .Z(n2919) );
  NR2 U1236 ( .A(n4599), .B(n4131), .Z(n3039) );
  NR2 U1237 ( .A(n4932), .B(n4109), .Z(n1703) );
  NR2 U1238 ( .A(n4290), .B(n4521), .Z(n1705) );
  NR2 U1239 ( .A(n4221), .B(n4417), .Z(n2383) );
  NR2 U1240 ( .A(n4908), .B(n4085), .Z(n3168) );
  NR2 U1241 ( .A(n4621), .B(n4754), .Z(n2805) );
  NR2 U1242 ( .A(n4957), .B(n4418), .Z(n2360) );
  ND2 U1243 ( .A(n4613), .B(n4739), .Z(n2947) );
  ND2 U1244 ( .A(n4613), .B(n4149), .Z(n2948) );
  ND2 U1245 ( .A(n4292), .B(n4816), .Z(n1931) );
  ND2 U1246 ( .A(n3260), .B(n3259), .Z(n1588) );
  ND2 U1247 ( .A(n4074), .B(n4432), .Z(n3259) );
  EO U1248 ( .A(n4890), .B(n4589), .Z(n3260) );
  ND2 U1249 ( .A(n1694), .B(n1693), .Z(n1554) );
  ND2 U1250 ( .A(n4631), .B(n4206), .Z(n1693) );
  MUX21L U1251 ( .A(n4838), .B(n1692), .S(n4291), .Z(n1694) );
  NR2 U1252 ( .A(n4631), .B(n4838), .Z(n1692) );
  ND2 U1253 ( .A(n1859), .B(n1858), .Z(n1558) );
  ND2 U1254 ( .A(n4259), .B(n4527), .Z(n1858) );
  EO U1255 ( .A(n4893), .B(n4630), .Z(n1859) );
  ND2 U1256 ( .A(n2449), .B(n2448), .Z(n1573) );
  ND2 U1257 ( .A(n4158), .B(n4406), .Z(n2448) );
  EO U1258 ( .A(n4886), .B(n4224), .Z(n2449) );
  ND2 U1259 ( .A(n2718), .B(n2717), .Z(n1578) );
  ND2 U1260 ( .A(n4218), .B(n4481), .Z(n2717) );
  MUX21L U1261 ( .A(n2716), .B(n4895), .S(n4218), .Z(n2718) );
  NR2 U1262 ( .A(n4894), .B(n4481), .Z(n2716) );
  ND2 U1263 ( .A(n2555), .B(n2554), .Z(n1575) );
  MUX21L U1264 ( .A(n2552), .B(n2553), .S(n4947), .Z(n2555) );
  ND2 U1265 ( .A(n2551), .B(n4596), .Z(n2554) );
  NR2 U1266 ( .A(n4596), .B(n4062), .Z(n2552) );
  ND2 U1267 ( .A(n2385), .B(n2384), .Z(n1572) );
  MUX21L U1268 ( .A(n2382), .B(n2383), .S(n4958), .Z(n2384) );
  MUX21L U1269 ( .A(n2380), .B(n2381), .S(n4570), .Z(n2385) );
  NR2 U1270 ( .A(n4570), .B(n4221), .Z(n2382) );
  ND2 U1271 ( .A(n2787), .B(n4039), .Z(n1579) );
  EO U1272 ( .A(n4887), .B(n4601), .Z(n2787) );
  ND2 U1273 ( .A(n2300), .B(n2299), .Z(n1568) );
  ND2 U1274 ( .A(n4287), .B(n4634), .Z(n2299) );
  MUX21L U1275 ( .A(n2298), .B(n4873), .S(n4634), .Z(n2300) );
  NR2 U1276 ( .A(n4287), .B(n4872), .Z(n2298) );
  ND2 U1277 ( .A(n2246), .B(n4552), .Z(n1567) );
  ND2 U1278 ( .A(n4953), .B(n4284), .Z(n2246) );
  ND2 U1279 ( .A(n4100), .B(n4751), .Z(n2837) );
  ND2 U1280 ( .A(n2038), .B(n2037), .Z(n1027) );
  ND2 U1281 ( .A(n4543), .B(n4806), .Z(n2037) );
  MUX21L U1282 ( .A(n4807), .B(n2036), .S(n4298), .Z(n2038) );
  MUX21L U1283 ( .A(n2830), .B(n4102), .S(n4619), .Z(n1581) );
  ND2 U1284 ( .A(n4896), .B(n4102), .Z(n2830) );
  MUX21L U1285 ( .A(n3064), .B(n4904), .S(n4251), .Z(n1586) );
  ND2 U1286 ( .A(n4904), .B(n4452), .Z(n3064) );
  MUX21L U1287 ( .A(n1897), .B(n1896), .S(n4258), .Z(n1559) );
  ND2 U1288 ( .A(n4939), .B(n4529), .Z(n1896) );
  ND2 U1289 ( .A(n4628), .B(n4939), .Z(n1897) );
  MUX21L U1290 ( .A(n1793), .B(n1792), .S(n4263), .Z(n1557) );
  ND2 U1291 ( .A(n4513), .B(n4830), .Z(n1792) );
  ND2 U1292 ( .A(n4936), .B(n4514), .Z(n1793) );
  MUX21L U1293 ( .A(n4051), .B(n4749), .S(n4608), .Z(n1577) );
  MUX21L U1294 ( .A(n2353), .B(n2352), .S(n4219), .Z(n1570) );
  ND2 U1295 ( .A(n4957), .B(n4419), .Z(n2352) );
  ND2 U1296 ( .A(n4569), .B(n4957), .Z(n2353) );
  MUX21L U1297 ( .A(n2341), .B(n4173), .S(n4632), .Z(n1569) );
  ND2 U1298 ( .A(n4173), .B(n4869), .Z(n2341) );
  ND2 U1299 ( .A(n2908), .B(n2907), .Z(n1046) );
  ND3 U1300 ( .A(n4615), .B(n4143), .C(n4914), .Z(n2907) );
  MUX21L U1301 ( .A(n2905), .B(n2906), .S(n4615), .Z(n2908) );
  NR2 U1302 ( .A(n4915), .B(n4143), .Z(n2906) );
  IVP U1303 ( .A(n4026), .Z(n4277) );
  IVP U1304 ( .A(n4034), .Z(n4230) );
  IVP U1305 ( .A(n4388), .Z(n4618) );
  AO7 U1306 ( .A(n4579), .B(n4798), .C(n4189), .Z(n1565) );
  NR2 U1307 ( .A(n4954), .B(n4167), .Z(n2381) );
  NR2 U1308 ( .A(n4277), .B(n4546), .Z(n2071) );
  ND3 U1309 ( .A(n4280), .B(n4799), .C(n4579), .Z(n1029) );
  ND3 U1310 ( .A(n2458), .B(n2457), .C(n2456), .Z(n1037) );
  ND2 U1311 ( .A(n4943), .B(n4157), .Z(n2457) );
  ND2 U1312 ( .A(n4592), .B(n4942), .Z(n2458) );
  ND2 U1313 ( .A(n4592), .B(n4158), .Z(n2456) );
  ND2 U1314 ( .A(n4088), .B(n4444), .Z(n1146) );
  ND2 U1315 ( .A(n4895), .B(n4056), .Z(n1576) );
  ND2 U1316 ( .A(n4298), .B(n4808), .Z(n1563) );
  MUX21L U1317 ( .A(n2227), .B(n2226), .S(n4952), .Z(n1532) );
  ND2 U1318 ( .A(n4187), .B(n4550), .Z(n2227) );
  ND2 U1319 ( .A(n4637), .B(n4283), .Z(n2226) );
  ND2 U1320 ( .A(n4195), .B(n4543), .Z(n2035) );
  ND2 U1321 ( .A(n1869), .B(n1868), .Z(n1022) );
  ND2 U1322 ( .A(n4259), .B(n4528), .Z(n1868) );
  EO U1323 ( .A(n4893), .B(n4259), .Z(n1869) );
  ND2 U1324 ( .A(n1782), .B(n1781), .Z(n1020) );
  ND2 U1325 ( .A(n4120), .B(n4514), .Z(n1781) );
  EO U1326 ( .A(n4892), .B(n4264), .Z(n1782) );
  ND2 U1327 ( .A(n1942), .B(n1941), .Z(n1024) );
  ND2 U1328 ( .A(n4292), .B(n4534), .Z(n1941) );
  MUX21L U1329 ( .A(n4922), .B(n1940), .S(n4626), .Z(n1942) );
  NR2 U1330 ( .A(n4922), .B(n4292), .Z(n1940) );
  ND2 U1331 ( .A(n1717), .B(n1716), .Z(n1019) );
  ND2 U1332 ( .A(n4933), .B(n4111), .Z(n1717) );
  ND2 U1333 ( .A(n4933), .B(n4520), .Z(n1716) );
  ND2 U1334 ( .A(n2575), .B(n4848), .Z(n1039) );
  EO U1335 ( .A(n4564), .B(n4230), .Z(n2575) );
  ND2 U1336 ( .A(n2491), .B(n2490), .Z(n1038) );
  ND2 U1337 ( .A(n4068), .B(n4401), .Z(n2491) );
  ND2 U1338 ( .A(n4944), .B(n4067), .Z(n2490) );
  MUX21L U1339 ( .A(n4875), .B(n2262), .S(n4636), .Z(n1032) );
  ND2 U1340 ( .A(n4285), .B(n4876), .Z(n2262) );
  MUX21L U1341 ( .A(n4417), .B(n4866), .S(n4220), .Z(n1034) );
  MUX21L U1342 ( .A(n2609), .B(n2608), .S(n4949), .Z(n1040) );
  ND2 U1343 ( .A(n4610), .B(n4058), .Z(n2609) );
  ND2 U1344 ( .A(n4211), .B(n4469), .Z(n2608) );
  MUX21L U1345 ( .A(n2753), .B(n2752), .S(n4243), .Z(n1043) );
  ND2 U1346 ( .A(n4901), .B(n4486), .Z(n2752) );
  ND2 U1347 ( .A(n4603), .B(n4901), .Z(n2753) );
  IVP U1348 ( .A(n4035), .Z(n4237) );
  IVP U1349 ( .A(n4390), .Z(n4605) );
  AO7 U1350 ( .A(n4254), .B(n4882), .C(n4421), .Z(n1566) );
  ND2 U1351 ( .A(n2389), .B(n2388), .Z(n1536) );
  MUX21L U1352 ( .A(n2386), .B(n4865), .S(n4221), .Z(n2388) );
  AO6 U1353 ( .A(n4221), .B(n4416), .C(n2387), .Z(n2389) );
  AO7 U1354 ( .A(n4583), .B(n4779), .C(n4089), .Z(n1049) );
  ND2 U1355 ( .A(n2355), .B(n2354), .Z(n1534) );
  ND2 U1356 ( .A(n4569), .B(n4171), .Z(n2354) );
  EN U1357 ( .A(n4888), .B(n4219), .Z(n2355) );
  ND2 U1358 ( .A(n3144), .B(n3143), .Z(n1551) );
  ND2 U1359 ( .A(n4087), .B(n4780), .Z(n3143) );
  EN U1360 ( .A(n4563), .B(n4232), .Z(n3144) );
  ND2 U1361 ( .A(n2926), .B(n2925), .Z(n1547) );
  ND2 U1362 ( .A(n4275), .B(n4505), .Z(n2925) );
  EO U1363 ( .A(n4888), .B(n4275), .Z(n2926) );
  ND2 U1364 ( .A(n2977), .B(n2976), .Z(n1548) );
  ND2 U1365 ( .A(n4271), .B(n4511), .Z(n2976) );
  EO U1366 ( .A(n4887), .B(n4611), .Z(n2977) );
  ND2 U1367 ( .A(n1953), .B(n4535), .Z(n1526) );
  EN U1368 ( .A(n4885), .B(n4293), .Z(n1953) );
  ND3 U1369 ( .A(n4459), .B(n4765), .C(n4153), .Z(n1076) );
  MUX21L U1370 ( .A(n4217), .B(n2699), .S(n4606), .Z(n1542) );
  ND2 U1371 ( .A(n4217), .B(n4764), .Z(n2699) );
  MUX21L U1372 ( .A(n2474), .B(n2473), .S(n4225), .Z(n1538) );
  ND2 U1373 ( .A(n4403), .B(n4856), .Z(n2473) );
  ND2 U1374 ( .A(n4593), .B(n4856), .Z(n2474) );
  MUX21L U1375 ( .A(n2650), .B(n2649), .S(n4214), .Z(n1541) );
  ND2 U1376 ( .A(n4472), .B(n4842), .Z(n2649) );
  ND2 U1377 ( .A(n4896), .B(n4472), .Z(n2650) );
  MUX21L U1378 ( .A(n2789), .B(n2788), .S(n4245), .Z(n1545) );
  ND2 U1379 ( .A(n4601), .B(n4901), .Z(n2789) );
  ND2 U1380 ( .A(n4901), .B(n4489), .Z(n2788) );
  MUX21L U1381 ( .A(n4631), .B(n1695), .S(n4932), .Z(n1520) );
  ND2 U1382 ( .A(n4631), .B(n4181), .Z(n1695) );
  ND2 U1383 ( .A(n1899), .B(n1898), .Z(n1525) );
  ND2 U1384 ( .A(n4132), .B(n4821), .Z(n1899) );
  ND2 U1385 ( .A(n4628), .B(n4821), .Z(n1898) );
  ND2 U1386 ( .A(n4216), .B(n4478), .Z(n1041) );
  ND2 U1387 ( .A(n1732), .B(n1731), .Z(n1521) );
  ND2 U1388 ( .A(n4573), .B(n4934), .Z(n1731) );
  MUX21L U1389 ( .A(n1730), .B(n4114), .S(n4934), .Z(n1732) );
  NR2 U1390 ( .A(n4573), .B(n4114), .Z(n1730) );
  ND2 U1391 ( .A(n1760), .B(n1759), .Z(n988) );
  MUX21L U1392 ( .A(n1757), .B(n4832), .S(n4574), .Z(n1759) );
  AO6 U1393 ( .A(n4574), .B(n4118), .C(n1758), .Z(n1760) );
  IVP U1394 ( .A(n4029), .Z(n4261) );
  AO7 U1395 ( .A(n4576), .B(n4830), .C(n4121), .Z(n1522) );
  NR2 U1396 ( .A(n4294), .B(n4536), .Z(n1527) );
  ND3 U1397 ( .A(n4251), .B(n4500), .C(n4913), .Z(n1546) );
  ND2 U1398 ( .A(n4631), .B(n4847), .Z(n2588) );
  ND2 U1399 ( .A(n4631), .B(n4059), .Z(n2589) );
  ND2 U1400 ( .A(n4583), .B(n4090), .Z(n1550) );
  ND2 U1401 ( .A(n1795), .B(n1794), .Z(n1523) );
  ND2 U1402 ( .A(n4122), .B(n4513), .Z(n1795) );
  ND2 U1403 ( .A(n4936), .B(n4122), .Z(n1794) );
  ND2 U1404 ( .A(n3079), .B(n3078), .Z(n1015) );
  MUX21L U1405 ( .A(n3076), .B(n3077), .S(n4252), .Z(n3079) );
  ND2 U1406 ( .A(n3075), .B(n4905), .Z(n3078) );
  NR2 U1407 ( .A(n4905), .B(n4451), .Z(n3076) );
  MUX21L U1408 ( .A(n2964), .B(n2963), .S(n4612), .Z(n1013) );
  ND2 U1409 ( .A(n4918), .B(n4151), .Z(n2964) );
  ND2 U1410 ( .A(n4272), .B(n4737), .Z(n2963) );
  MUX21L U1411 ( .A(n2312), .B(n4955), .S(n4287), .Z(n999) );
  ND2 U1412 ( .A(n4955), .B(n4634), .Z(n2312) );
  AO7 U1413 ( .A(n4215), .B(n4477), .C(n2678), .Z(n1006) );
  ND2 U1414 ( .A(n4902), .B(n4607), .Z(n2678) );
  MUX21L U1415 ( .A(n2502), .B(n2501), .S(n4945), .Z(n1004) );
  ND2 U1416 ( .A(n4594), .B(n4067), .Z(n2502) );
  ND2 U1417 ( .A(n4594), .B(n4227), .Z(n2501) );
  ND2 U1418 ( .A(n4295), .B(n4538), .Z(n1979) );
  AN3 U1419 ( .A(n4234), .B(n4783), .C(n4584), .Z(n423) );
  ND2 U1420 ( .A(n2867), .B(n2866), .Z(n1011) );
  ND2 U1421 ( .A(n4499), .B(n4745), .Z(n2866) );
  MUX21L U1422 ( .A(n4746), .B(n2865), .S(n4250), .Z(n2867) );
  ND2 U1423 ( .A(n2133), .B(n2132), .Z(n995) );
  ND2 U1424 ( .A(n4424), .B(n4799), .Z(n2132) );
  MUX21L U1425 ( .A(n4799), .B(n2131), .S(n4281), .Z(n2133) );
  ND2 U1426 ( .A(n2367), .B(n2366), .Z(n1000) );
  ND3 U1427 ( .A(n4570), .B(n4171), .C(n4958), .Z(n2366) );
  MUX21L U1428 ( .A(n2364), .B(n2365), .S(n4570), .Z(n2367) );
  NR2 U1429 ( .A(n4958), .B(n4170), .Z(n2365) );
  IVP U1430 ( .A(n4723), .Z(n4945) );
  IVP U1431 ( .A(n4038), .Z(n4252) );
  IVP U1432 ( .A(n4730), .Z(n4905) );
  IVP U1433 ( .A(n4030), .Z(n4257) );
  IVP U1434 ( .A(n4389), .Z(n4612) );
  IVP U1435 ( .A(n4731), .Z(n4899) );
  AO6 U1436 ( .A(n4630), .B(n4126), .C(n1839), .Z(n1841) );
  NR2 U1437 ( .A(n4937), .B(n4260), .Z(n1839) );
  AO7 U1438 ( .A(n4224), .B(n4405), .C(n4857), .Z(n1003) );
  NR2 U1439 ( .A(n4947), .B(n4398), .Z(n1005) );
  ND2 U1440 ( .A(n2701), .B(n2700), .Z(n1508) );
  ND2 U1441 ( .A(n4048), .B(n4764), .Z(n2700) );
  EN U1442 ( .A(n4560), .B(n4217), .Z(n2701) );
  ND2 U1443 ( .A(n2766), .B(n2765), .Z(n1509) );
  ND2 U1444 ( .A(n4602), .B(n4040), .Z(n2765) );
  EO U1445 ( .A(n4886), .B(n4244), .Z(n2766) );
  ND2 U1446 ( .A(n2247), .B(n4552), .Z(n1498) );
  EO U1447 ( .A(n4889), .B(n4284), .Z(n2247) );
  ND2 U1448 ( .A(n1936), .B(n1935), .Z(n1491) );
  ND2 U1449 ( .A(n1932), .B(n4816), .Z(n1935) );
  MUX21L U1450 ( .A(n1933), .B(n1934), .S(n4626), .Z(n1936) );
  NR2 U1451 ( .A(n4292), .B(n4626), .Z(n1932) );
  ND2 U1452 ( .A(n2278), .B(n2277), .Z(n1499) );
  ND2 U1453 ( .A(n2274), .B(n4954), .Z(n2277) );
  MUX21L U1454 ( .A(n2275), .B(n2276), .S(n4954), .Z(n2278) );
  NR2 U1455 ( .A(n4635), .B(n4286), .Z(n2274) );
  ND2 U1456 ( .A(n3147), .B(n3146), .Z(n1517) );
  ND2 U1457 ( .A(n4583), .B(n4780), .Z(n3146) );
  MUX21L U1458 ( .A(n4780), .B(n3145), .S(n4232), .Z(n3147) );
  NR2 U1459 ( .A(n4583), .B(n4781), .Z(n3145) );
  MUX21L U1460 ( .A(n1838), .B(n4824), .S(n4630), .Z(n1840) );
  MUX21L U1461 ( .A(n2739), .B(n4044), .S(n4604), .Z(n1007) );
  ND2 U1462 ( .A(n4045), .B(n4760), .Z(n2739) );
  ND2 U1463 ( .A(n2230), .B(n2229), .Z(n967) );
  ND2 U1464 ( .A(n4550), .B(n4878), .Z(n2229) );
  MUX21L U1465 ( .A(n4550), .B(n2228), .S(n4283), .Z(n2230) );
  IVP U1466 ( .A(n4387), .Z(n4620) );
  IVP U1467 ( .A(n4023), .Z(n4296) );
  IVP U1468 ( .A(n4731), .Z(n4897) );
  IVP U1469 ( .A(n4385), .Z(n4635) );
  AO7 U1470 ( .A(n4250), .B(n4498), .C(n4748), .Z(n1512) );
  NR2 U1471 ( .A(n4922), .B(n4205), .Z(n1934) );
  NR2 U1472 ( .A(n4635), .B(n4181), .Z(n2275) );
  NR2 U1473 ( .A(n4623), .B(n4810), .Z(n1989) );
  NR2 U1474 ( .A(n4623), .B(n4200), .Z(n1990) );
  MUX21L U1475 ( .A(n1988), .B(n4295), .S(n4924), .Z(n1991) );
  NR2 U1476 ( .A(n4296), .B(n4539), .Z(n1988) );
  ND3 U1477 ( .A(n1974), .B(n1973), .C(n1972), .Z(n1492) );
  ND2 U1478 ( .A(n4201), .B(n4812), .Z(n1973) );
  ND2 U1479 ( .A(n4624), .B(n4812), .Z(n1974) );
  ND2 U1480 ( .A(n4624), .B(n4201), .Z(n1972) );
  ND3 U1481 ( .A(n2477), .B(n2476), .C(n2475), .Z(n1504) );
  ND2 U1482 ( .A(n4070), .B(n4403), .Z(n2476) );
  ND2 U1483 ( .A(n4943), .B(n4403), .Z(n2477) );
  ND2 U1484 ( .A(n4943), .B(n4070), .Z(n2475) );
  ND2 U1485 ( .A(n4228), .B(n4852), .Z(n2523) );
  ND2 U1486 ( .A(n4946), .B(n4065), .Z(n2524) );
  MUX21L U1487 ( .A(n2463), .B(n4072), .S(n4592), .Z(n1503) );
  ND2 U1488 ( .A(n4943), .B(n4156), .Z(n2463) );
  AO7 U1489 ( .A(n4639), .B(n4193), .C(n2069), .Z(n1495) );
  ND2 U1490 ( .A(n4928), .B(n4300), .Z(n2069) );
  MUX21L U1491 ( .A(n4273), .B(n2949), .S(n4917), .Z(n1514) );
  ND2 U1492 ( .A(n4273), .B(n4506), .Z(n2949) );
  MUX21L U1493 ( .A(n4501), .B(n2883), .S(n4277), .Z(n1513) );
  ND2 U1494 ( .A(n4914), .B(n4501), .Z(n2883) );
  MUX21L U1495 ( .A(n3066), .B(n3065), .S(n4600), .Z(n1516) );
  ND2 U1496 ( .A(n4094), .B(n4773), .Z(n3065) );
  ND2 U1497 ( .A(n4905), .B(n4094), .Z(n3066) );
  ND2 U1498 ( .A(n4043), .B(n4758), .Z(n2745) );
  AO7 U1499 ( .A(n4568), .B(n4168), .C(n2374), .Z(n970) );
  ND2 U1500 ( .A(n4958), .B(n4220), .Z(n2374) );
  AN3 U1501 ( .A(n4107), .B(n4837), .C(n4631), .Z(n424) );
  MUX21L U1502 ( .A(n4519), .B(n4834), .S(n4289), .Z(n1486) );
  ND2 U1503 ( .A(n2392), .B(n2391), .Z(n1502) );
  ND2 U1504 ( .A(n4221), .B(n4865), .Z(n2391) );
  MUX21L U1505 ( .A(n4416), .B(n2390), .S(n4940), .Z(n2392) );
  NR2 U1506 ( .A(n4221), .B(n4416), .Z(n2390) );
  MUX21L U1507 ( .A(n4866), .B(n4168), .S(n4570), .Z(n1500) );
  MUX21L U1508 ( .A(n4927), .B(n4545), .S(n4298), .Z(n1494) );
  MUX21L U1509 ( .A(n4620), .B(n4103), .S(n4897), .Z(n1511) );
  ND2 U1510 ( .A(n2810), .B(n2809), .Z(n981) );
  ND2 U1511 ( .A(n4899), .B(n4492), .Z(n2809) );
  MUX21L U1512 ( .A(n4492), .B(n2808), .S(n4247), .Z(n2810) );
  NR2 U1513 ( .A(n4899), .B(n4491), .Z(n2808) );
  IVP U1514 ( .A(n4027), .Z(n4274) );
  ND2 U1515 ( .A(n2528), .B(n2527), .Z(n1472) );
  MUX21L U1516 ( .A(n4946), .B(n2525), .S(n4595), .Z(n2527) );
  AO6 U1517 ( .A(n4946), .B(n4064), .C(n2526), .Z(n2528) );
  NR2 U1518 ( .A(n4946), .B(n4064), .Z(n2525) );
  ND3 U1519 ( .A(n2408), .B(n2407), .C(n2406), .Z(n1002) );
  ND2 U1520 ( .A(n4413), .B(n4862), .Z(n2408) );
  ND2 U1521 ( .A(n4166), .B(n4413), .Z(n2407) );
  ND2 U1522 ( .A(n4166), .B(n4863), .Z(n2406) );
  ND3 U1523 ( .A(n2612), .B(n2611), .C(n2610), .Z(n976) );
  ND2 U1524 ( .A(n4469), .B(n4846), .Z(n2611) );
  ND2 U1525 ( .A(n4210), .B(n4469), .Z(n2610) );
  ND2 U1526 ( .A(n4211), .B(n4846), .Z(n2612) );
  ND2 U1527 ( .A(n4196), .B(n4809), .Z(n2022) );
  MUX21L U1528 ( .A(n2293), .B(n2292), .S(n4954), .Z(n968) );
  ND2 U1529 ( .A(n4180), .B(n4556), .Z(n2293) );
  ND2 U1530 ( .A(n4634), .B(n4286), .Z(n2292) );
  ND2 U1531 ( .A(n4274), .B(n4740), .Z(n2927) );
  ND2 U1532 ( .A(n4905), .B(n4451), .Z(n3080) );
  ND2 U1533 ( .A(n4905), .B(n4092), .Z(n3081) );
  MUX21L U1534 ( .A(n2539), .B(n2538), .S(n4228), .Z(n975) );
  ND2 U1535 ( .A(n4947), .B(n4448), .Z(n2538) );
  ND2 U1536 ( .A(n4596), .B(n4947), .Z(n2539) );
  ND2 U1537 ( .A(n2434), .B(n2433), .Z(n973) );
  ND2 U1538 ( .A(n4410), .B(n4858), .Z(n2434) );
  ND2 U1539 ( .A(n4223), .B(n4410), .Z(n2433) );
  ND2 U1540 ( .A(n2410), .B(n2409), .Z(n972) );
  ND2 U1541 ( .A(n4165), .B(n4862), .Z(n2410) );
  ND2 U1542 ( .A(n4568), .B(n4165), .Z(n2409) );
  ND2 U1543 ( .A(n2693), .B(n4050), .Z(n977) );
  ND2 U1544 ( .A(n4903), .B(n4606), .Z(n2693) );
  IVP U1545 ( .A(n4729), .Z(n4909) );
  IVP U1546 ( .A(n4387), .Z(n4622) );
  IVP U1547 ( .A(n4389), .Z(n4609) );
  IVP U1548 ( .A(n4393), .Z(n4585) );
  NR2 U1549 ( .A(n4951), .B(n4547), .Z(n2201) );
  ND2 U1550 ( .A(n2013), .B(n2012), .Z(n1459) );
  ND2 U1551 ( .A(n4296), .B(n4809), .Z(n2012) );
  EO U1552 ( .A(n4885), .B(n4622), .Z(n2013) );
  ND2 U1553 ( .A(n2137), .B(n2136), .Z(n1463) );
  ND2 U1554 ( .A(n4281), .B(n4798), .Z(n2136) );
  EO U1555 ( .A(n4561), .B(n4281), .Z(n2137) );
  ND2 U1556 ( .A(n3214), .B(n3213), .Z(n1484) );
  ND2 U1557 ( .A(n4079), .B(n4788), .Z(n3213) );
  EN U1558 ( .A(n4565), .B(n4237), .Z(n3214) );
  ND2 U1559 ( .A(n2881), .B(n4500), .Z(n1479) );
  EO U1560 ( .A(n4892), .B(n4251), .Z(n2881) );
  ND2 U1561 ( .A(n4467), .B(n4847), .Z(n2590) );
  MUX21L U1562 ( .A(n2652), .B(n2651), .S(n4214), .Z(n1474) );
  ND2 U1563 ( .A(n4472), .B(n4841), .Z(n2651) );
  ND2 U1564 ( .A(n4897), .B(n4473), .Z(n2652) );
  MUX21L U1565 ( .A(n2372), .B(n2371), .S(n4958), .Z(n1468) );
  ND2 U1566 ( .A(n4220), .B(n4418), .Z(n2372) );
  ND2 U1567 ( .A(n4571), .B(n4220), .Z(n2371) );
  MUX21L U1568 ( .A(n2998), .B(n2997), .S(n4270), .Z(n1481) );
  ND2 U1569 ( .A(n4459), .B(n4766), .Z(n2997) );
  ND2 U1570 ( .A(n4919), .B(n4597), .Z(n2998) );
  MUX21L U1571 ( .A(n1733), .B(n4115), .S(n4934), .Z(n1735) );
  NR2 U1572 ( .A(n4573), .B(n4114), .Z(n1733) );
  ND2 U1573 ( .A(n1798), .B(n1797), .Z(n1456) );
  ND2 U1574 ( .A(n4936), .B(n4512), .Z(n1797) );
  MUX21L U1575 ( .A(n4513), .B(n1796), .S(n4263), .Z(n1798) );
  NR2 U1576 ( .A(n4936), .B(n4512), .Z(n1796) );
  ND2 U1577 ( .A(n2333), .B(n2332), .Z(n1467) );
  ND2 U1578 ( .A(n4288), .B(n4466), .Z(n2332) );
  MUX21L U1579 ( .A(n2331), .B(n4956), .S(n4288), .Z(n2333) );
  NR2 U1580 ( .A(n4956), .B(n4465), .Z(n2331) );
  ND2 U1581 ( .A(n3099), .B(n3098), .Z(n1482) );
  ND2 U1582 ( .A(n4091), .B(n4776), .Z(n3098) );
  MUX21L U1583 ( .A(n4448), .B(n3097), .S(n4253), .Z(n3099) );
  ND2 U1584 ( .A(n2437), .B(n2436), .Z(n942) );
  ND2 U1585 ( .A(n4942), .B(n4409), .Z(n2436) );
  MUX21L U1586 ( .A(n2435), .B(n4160), .S(n4942), .Z(n2437) );
  ND2 U1587 ( .A(n2203), .B(n2202), .Z(n938) );
  ND2 U1588 ( .A(n2199), .B(n4880), .Z(n2202) );
  MUX21L U1589 ( .A(n2200), .B(n2201), .S(n4282), .Z(n2203) );
  NR2 U1590 ( .A(n4282), .B(n4638), .Z(n2199) );
  IVP U1591 ( .A(n4037), .Z(n4249) );
  IVP U1592 ( .A(n4038), .Z(n4253) );
  IVP U1593 ( .A(n4393), .Z(n4588) );
  NR2 U1594 ( .A(n4289), .B(n4519), .Z(n1737) );
  NR2 U1595 ( .A(n4629), .B(n4823), .Z(n1871) );
  NR2 U1596 ( .A(n4629), .B(n4129), .Z(n1872) );
  ND2 U1597 ( .A(n1874), .B(n1873), .Z(n932) );
  MUX21L U1598 ( .A(n1870), .B(n4259), .S(n4938), .Z(n1873) );
  NR2 U1599 ( .A(n1872), .B(n1871), .Z(n1874) );
  NR2 U1600 ( .A(n4259), .B(n4528), .Z(n1870) );
  ND2 U1601 ( .A(n1784), .B(n1783), .Z(n930) );
  ND2 U1602 ( .A(n4264), .B(n4514), .Z(n1783) );
  EO U1603 ( .A(n4892), .B(n4264), .Z(n1784) );
  ND2 U1604 ( .A(n3014), .B(n3013), .Z(n953) );
  ND2 U1605 ( .A(n4154), .B(n4768), .Z(n3013) );
  EN U1606 ( .A(n4560), .B(n4268), .Z(n3014) );
  ND3 U1607 ( .A(n4231), .B(n4445), .C(n4907), .Z(n954) );
  ND2 U1608 ( .A(n2191), .B(n2190), .Z(n1465) );
  ND2 U1609 ( .A(n4638), .B(n4188), .Z(n2191) );
  ND2 U1610 ( .A(n4638), .B(n4882), .Z(n2190) );
  ND2 U1611 ( .A(n4572), .B(n4836), .Z(n1718) );
  ND2 U1612 ( .A(n4627), .B(n4820), .Z(n1909) );
  ND2 U1613 ( .A(n4627), .B(n4134), .Z(n1910) );
  MUX21L U1614 ( .A(n4249), .B(n2838), .S(n4895), .Z(n950) );
  ND2 U1615 ( .A(n4249), .B(n4496), .Z(n2838) );
  AO7 U1616 ( .A(n4910), .B(n4081), .C(n3198), .Z(n955) );
  ND2 U1617 ( .A(n4586), .B(n4236), .Z(n3198) );
  MUX21L U1618 ( .A(n2933), .B(n4147), .S(n4614), .Z(n951) );
  ND2 U1619 ( .A(n4916), .B(n4147), .Z(n2933) );
  MUX21L U1620 ( .A(n3233), .B(n3232), .S(n4588), .Z(n956) );
  ND2 U1621 ( .A(n4077), .B(n4791), .Z(n3233) );
  ND2 U1622 ( .A(n4238), .B(n4791), .Z(n3232) );
  AN3 U1623 ( .A(n4211), .B(n4845), .C(n4610), .Z(n425) );
  MUX21L U1624 ( .A(n4501), .B(n4914), .S(n4277), .Z(n1480) );
  ND2 U1625 ( .A(n1958), .B(n1957), .Z(n934) );
  ND2 U1626 ( .A(n4293), .B(n4625), .Z(n1957) );
  MUX21L U1627 ( .A(n1956), .B(n4815), .S(n4625), .Z(n1958) );
  NR2 U1628 ( .A(n4293), .B(n4814), .Z(n1956) );
  ND2 U1629 ( .A(n2985), .B(n2984), .Z(n952) );
  ND2 U1630 ( .A(n4271), .B(n4431), .Z(n2984) );
  MUX21L U1631 ( .A(n2983), .B(n4918), .S(n4271), .Z(n2985) );
  NR2 U1632 ( .A(n4919), .B(n4559), .Z(n2983) );
  IVP U1633 ( .A(n4392), .Z(n4591) );
  ND2 U1634 ( .A(n2793), .B(n2792), .Z(n1444) );
  MUX21L U1635 ( .A(n2790), .B(n4755), .S(n4246), .Z(n2792) );
  AO6 U1636 ( .A(n4246), .B(n4489), .C(n2791), .Z(n2793) );
  AO7 U1637 ( .A(n4247), .B(n4753), .C(n4621), .Z(n949) );
  NR2 U1638 ( .A(n4937), .B(n4428), .Z(n1822) );
  NR2 U1639 ( .A(n4937), .B(n4124), .Z(n1823) );
  NR2 U1640 ( .A(n4569), .B(n4864), .Z(n2395) );
  ND2 U1641 ( .A(n2991), .B(n4734), .Z(n1447) );
  EO U1642 ( .A(n4560), .B(n4270), .Z(n2991) );
  ND2 U1643 ( .A(n2499), .B(n4854), .Z(n1437) );
  EN U1644 ( .A(n4563), .B(n4227), .Z(n2499) );
  ND2 U1645 ( .A(n2240), .B(n2239), .Z(n1430) );
  ND2 U1646 ( .A(n4284), .B(n4878), .Z(n2239) );
  EO U1647 ( .A(n4889), .B(n4637), .Z(n2240) );
  ND3 U1648 ( .A(n2704), .B(n2703), .C(n2702), .Z(n1441) );
  ND2 U1649 ( .A(n4047), .B(n4479), .Z(n2703) );
  ND2 U1650 ( .A(n4902), .B(n4479), .Z(n2704) );
  ND2 U1651 ( .A(n4902), .B(n4048), .Z(n2702) );
  ND3 U1652 ( .A(n4489), .B(n4755), .C(n4039), .Z(n979) );
  ND2 U1653 ( .A(n2305), .B(n2304), .Z(n1432) );
  ND2 U1654 ( .A(n4955), .B(n4559), .Z(n2305) );
  ND2 U1655 ( .A(n4287), .B(n4558), .Z(n2304) );
  ND2 U1656 ( .A(n4954), .B(n4179), .Z(n1466) );
  ND2 U1657 ( .A(n4227), .B(n4400), .Z(n943) );
  MUX21L U1658 ( .A(n1821), .B(n4261), .S(n4577), .Z(n1824) );
  NR2 U1659 ( .A(n4261), .B(n4826), .Z(n1821) );
  ND2 U1660 ( .A(n2423), .B(n2422), .Z(n1436) );
  ND2 U1661 ( .A(n4591), .B(n4161), .Z(n2422) );
  MUX21L U1662 ( .A(n4860), .B(n2421), .S(n4223), .Z(n2423) );
  NR2 U1663 ( .A(n4591), .B(n4860), .Z(n2421) );
  ND2 U1664 ( .A(n2397), .B(n2396), .Z(n1435) );
  ND2 U1665 ( .A(n2393), .B(n4415), .Z(n2396) );
  MUX21L U1666 ( .A(n2394), .B(n2395), .S(n4221), .Z(n2397) );
  NR2 U1667 ( .A(n4940), .B(n4221), .Z(n2393) );
  ND2 U1668 ( .A(n2102), .B(n2101), .Z(n1428) );
  ND2 U1669 ( .A(n4279), .B(n4427), .Z(n2101) );
  MUX21L U1670 ( .A(n4929), .B(n2100), .S(n4578), .Z(n2102) );
  NR2 U1671 ( .A(n4929), .B(n4279), .Z(n2100) );
  MUX21L U1672 ( .A(n2232), .B(n2233), .S(n4952), .Z(n2235) );
  NR2 U1673 ( .A(n4637), .B(n4186), .Z(n2232) );
  ND2 U1674 ( .A(n2544), .B(n2543), .Z(n916) );
  ND2 U1675 ( .A(n2540), .B(n4852), .Z(n2543) );
  MUX21L U1676 ( .A(n2541), .B(n2542), .S(n4229), .Z(n2544) );
  NR2 U1677 ( .A(n4229), .B(n4596), .Z(n2540) );
  ND2 U1678 ( .A(n2041), .B(n2040), .Z(n909) );
  ND2 U1679 ( .A(n4543), .B(n4806), .Z(n2040) );
  MUX21L U1680 ( .A(n4806), .B(n2039), .S(n4298), .Z(n2041) );
  IVP U1681 ( .A(n4388), .Z(n4616) );
  IVP U1682 ( .A(n4729), .Z(n4912) );
  AO7 U1683 ( .A(n4901), .B(n4488), .C(n4041), .Z(n1442) );
  ND2 U1684 ( .A(n1845), .B(n1844), .Z(n904) );
  MUX21L U1685 ( .A(n1842), .B(n4824), .S(n4630), .Z(n1844) );
  AO6 U1686 ( .A(n4630), .B(n4126), .C(n1843), .Z(n1845) );
  NR2 U1687 ( .A(n4947), .B(n4464), .Z(n2542) );
  ND2 U1688 ( .A(n4277), .B(n4744), .Z(n2884) );
  ND2 U1689 ( .A(n2257), .B(n2256), .Z(n1431) );
  ND2 U1690 ( .A(n4182), .B(n4877), .Z(n2257) );
  ND2 U1691 ( .A(n4636), .B(n4182), .Z(n2256) );
  ND2 U1692 ( .A(n4288), .B(n4871), .Z(n2316) );
  ND2 U1693 ( .A(n2172), .B(n2171), .Z(n911) );
  ND2 U1694 ( .A(n4254), .B(n4421), .Z(n2171) );
  MUX21L U1695 ( .A(n2170), .B(n4950), .S(n4255), .Z(n2172) );
  NR2 U1696 ( .A(n4950), .B(n4421), .Z(n2170) );
  ND2 U1697 ( .A(n1763), .B(n1762), .Z(n902) );
  ND2 U1698 ( .A(n4574), .B(n4832), .Z(n1762) );
  MUX21L U1699 ( .A(n1761), .B(n4118), .S(n4574), .Z(n1763) );
  ND2 U1700 ( .A(n1815), .B(n1814), .Z(n903) );
  ND2 U1701 ( .A(n4429), .B(n4828), .Z(n1814) );
  MUX21L U1702 ( .A(n4429), .B(n1813), .S(n4262), .Z(n1815) );
  ND2 U1703 ( .A(n1952), .B(n1951), .Z(n906) );
  ND2 U1704 ( .A(n4625), .B(n4203), .Z(n1951) );
  EO U1705 ( .A(n4885), .B(n4293), .Z(n1952) );
  MUX21L U1706 ( .A(n2840), .B(n2839), .S(n4618), .Z(n922) );
  ND2 U1707 ( .A(n4099), .B(n4750), .Z(n2840) );
  ND2 U1708 ( .A(n4249), .B(n4750), .Z(n2839) );
  AN3 U1709 ( .A(n4092), .B(n4774), .C(n4581), .Z(n426) );
  MUX21L U1710 ( .A(n2058), .B(n2057), .S(n4640), .Z(n1427) );
  ND2 U1711 ( .A(n4299), .B(n4803), .Z(n2057) );
  ND2 U1712 ( .A(n4928), .B(n4299), .Z(n2058) );
  MUX21L U1713 ( .A(n1981), .B(n4201), .S(n4924), .Z(n1983) );
  ND2 U1714 ( .A(n1752), .B(n1751), .Z(n1391) );
  ND2 U1715 ( .A(n4117), .B(n4516), .Z(n1751) );
  EN U1716 ( .A(n4891), .B(n4265), .Z(n1752) );
  AO7 U1717 ( .A(n4958), .B(n4417), .C(n4168), .Z(n1433) );
  NR2 U1718 ( .A(n4258), .B(n4823), .Z(n1883) );
  ND2 U1719 ( .A(n4254), .B(n4420), .Z(n1429) );
  ND2 U1720 ( .A(n4263), .B(n4414), .Z(n1799) );
  ND2 U1721 ( .A(n4933), .B(n4110), .Z(n1708) );
  ND2 U1722 ( .A(n2635), .B(n4843), .Z(n1407) );
  EO U1723 ( .A(n4562), .B(n4213), .Z(n2635) );
  ND2 U1724 ( .A(n2479), .B(n2478), .Z(n1406) );
  ND2 U1725 ( .A(n4943), .B(n4070), .Z(n2478) );
  EN U1726 ( .A(n4885), .B(n4593), .Z(n2479) );
  ND2 U1727 ( .A(n4924), .B(n4538), .Z(n1982) );
  ND2 U1728 ( .A(n4257), .B(n4530), .Z(n1911) );
  ND2 U1729 ( .A(n3172), .B(n3171), .Z(n926) );
  ND2 U1730 ( .A(n4085), .B(n4783), .Z(n3172) );
  ND2 U1731 ( .A(n4584), .B(n4085), .Z(n3171) );
  ND2 U1732 ( .A(n1902), .B(n1901), .Z(n1394) );
  ND2 U1733 ( .A(n4628), .B(n4132), .Z(n1901) );
  MUX21L U1734 ( .A(n1900), .B(n4133), .S(n4939), .Z(n1902) );
  NR2 U1735 ( .A(n4628), .B(n4132), .Z(n1900) );
  ND2 U1736 ( .A(n2859), .B(n2858), .Z(n1413) );
  MUX21L U1737 ( .A(n2856), .B(n2857), .S(n4617), .Z(n2858) );
  MUX21L U1738 ( .A(n2854), .B(n2855), .S(n4894), .Z(n2859) );
  NR2 U1739 ( .A(n4250), .B(n4748), .Z(n2856) );
  ND2 U1740 ( .A(n3069), .B(n3068), .Z(n1417) );
  ND2 U1741 ( .A(n4600), .B(n4773), .Z(n3068) );
  MUX21L U1742 ( .A(n3067), .B(n4094), .S(n4600), .Z(n3069) );
  ND2 U1743 ( .A(n2460), .B(n2459), .Z(n887) );
  ND2 U1744 ( .A(n4592), .B(n4157), .Z(n2459) );
  EO U1745 ( .A(n4885), .B(n4224), .Z(n2460) );
  IVP U1746 ( .A(n4033), .Z(n4226) );
  AO7 U1747 ( .A(n4235), .B(n4439), .C(n4785), .Z(n1418) );
  AO7 U1748 ( .A(n4952), .B(n4551), .C(n2241), .Z(n1399) );
  ND2 U1749 ( .A(n4637), .B(n4284), .Z(n2241) );
  AO7 U1750 ( .A(n4288), .B(n4869), .C(n4466), .Z(n1401) );
  NR2 U1751 ( .A(n4617), .B(n4097), .Z(n2854) );
  ND2 U1752 ( .A(n4141), .B(n4744), .Z(n2885) );
  ND2 U1753 ( .A(n4229), .B(n4464), .Z(n2545) );
  ND2 U1754 ( .A(n4229), .B(n4851), .Z(n2547) );
  ND2 U1755 ( .A(n3216), .B(n3215), .Z(n1419) );
  ND2 U1756 ( .A(n4438), .B(n4789), .Z(n3216) );
  ND2 U1757 ( .A(n4237), .B(n4438), .Z(n3215) );
  ND2 U1758 ( .A(n2281), .B(n2280), .Z(n1400) );
  ND2 U1759 ( .A(n4286), .B(n4954), .Z(n2280) );
  MUX21L U1760 ( .A(n2279), .B(n4635), .S(n4954), .Z(n2281) );
  NR2 U1761 ( .A(n4635), .B(n4286), .Z(n2279) );
  ND2 U1762 ( .A(n2104), .B(n2103), .Z(n1398) );
  ND2 U1763 ( .A(n4191), .B(n4427), .Z(n2103) );
  EN U1764 ( .A(n4887), .B(n4279), .Z(n2104) );
  ND2 U1765 ( .A(n4605), .B(n4047), .Z(n2709) );
  ND2 U1766 ( .A(n2208), .B(n2207), .Z(n883) );
  ND2 U1767 ( .A(n2204), .B(n4880), .Z(n2207) );
  MUX21L U1768 ( .A(n2205), .B(n2206), .S(n4282), .Z(n2208) );
  NR2 U1769 ( .A(n4282), .B(n4638), .Z(n2204) );
  ND2 U1770 ( .A(n2267), .B(n2266), .Z(n884) );
  ND2 U1771 ( .A(n4635), .B(n4182), .Z(n2266) );
  MUX21L U1772 ( .A(n4875), .B(n2265), .S(n4285), .Z(n2267) );
  NR2 U1773 ( .A(n4635), .B(n4875), .Z(n2265) );
  ND2 U1774 ( .A(n1945), .B(n1944), .Z(n877) );
  ND2 U1775 ( .A(n4923), .B(n4534), .Z(n1944) );
  MUX21L U1776 ( .A(n4535), .B(n1943), .S(n4292), .Z(n1945) );
  NR2 U1777 ( .A(n4923), .B(n4534), .Z(n1943) );
  ND2 U1778 ( .A(n3116), .B(n3115), .Z(n897) );
  ND2 U1779 ( .A(n4446), .B(n4777), .Z(n3115) );
  MUX21L U1780 ( .A(n4777), .B(n3114), .S(n4254), .Z(n3116) );
  ND2 U1781 ( .A(n3193), .B(n3192), .Z(n898) );
  ND2 U1782 ( .A(n4082), .B(n4786), .Z(n3192) );
  EO U1783 ( .A(n4892), .B(n4586), .Z(n3193) );
  MUX21L U1784 ( .A(n4743), .B(n2886), .S(n4276), .Z(n1414) );
  ND2 U1785 ( .A(n4616), .B(n4744), .Z(n2886) );
  MUX21L U1786 ( .A(n4267), .B(n4453), .S(n4921), .Z(n1416) );
  MUX21L U1787 ( .A(n4149), .B(n4613), .S(n4917), .Z(n1415) );
  MUX21L U1788 ( .A(n2356), .B(n4957), .S(n4219), .Z(n1402) );
  ND2 U1789 ( .A(n4957), .B(n4569), .Z(n2356) );
  MUX21L U1790 ( .A(n4763), .B(n2708), .S(n4218), .Z(n2710) );
  NR2 U1791 ( .A(n4605), .B(n4763), .Z(n2708) );
  ND2 U1792 ( .A(n3018), .B(n3017), .Z(n896) );
  ND3 U1793 ( .A(n4598), .B(n4154), .C(n4920), .Z(n3017) );
  MUX21L U1794 ( .A(n3015), .B(n3016), .S(n4598), .Z(n3018) );
  NR2 U1795 ( .A(n4920), .B(n4154), .Z(n3016) );
  NR2 U1796 ( .A(n4951), .B(n4548), .Z(n2206) );
  NR2 U1797 ( .A(n4567), .B(n4140), .Z(n2174) );
  ND2 U1798 ( .A(n4111), .B(n4836), .Z(n1719) );
  ND2 U1799 ( .A(n4623), .B(n4200), .Z(n1984) );
  ND2 U1800 ( .A(n4262), .B(n4829), .Z(n1808) );
  ND2 U1801 ( .A(n4262), .B(n4430), .Z(n1809) );
  ND2 U1802 ( .A(n1722), .B(n1721), .Z(n872) );
  ND2 U1803 ( .A(n4572), .B(n4112), .Z(n1721) );
  MUX21L U1804 ( .A(n1720), .B(n4112), .S(n4933), .Z(n1722) );
  NR2 U1805 ( .A(n4572), .B(n4112), .Z(n1720) );
  AN3 U1806 ( .A(n4144), .B(n4741), .C(n4615), .Z(n427) );
  ND2 U1807 ( .A(n3220), .B(n3219), .Z(n1388) );
  AO6 U1808 ( .A(n4237), .B(n4437), .C(n3218), .Z(n3220) );
  MUX21L U1809 ( .A(n3217), .B(n4789), .S(n4237), .Z(n3219) );
  NR2 U1810 ( .A(n4911), .B(n4587), .Z(n3218) );
  MUX21L U1811 ( .A(n4516), .B(n1764), .S(n4265), .Z(n873) );
  ND2 U1812 ( .A(n4516), .B(n4831), .Z(n1764) );
  MUX21L U1813 ( .A(n2812), .B(n2811), .S(n4899), .Z(n893) );
  ND2 U1814 ( .A(n4106), .B(n4492), .Z(n2812) );
  ND2 U1815 ( .A(n4621), .B(n4105), .Z(n2811) );
  MUX21L U1816 ( .A(n4736), .B(n2965), .S(n4272), .Z(n895) );
  ND2 U1817 ( .A(n4612), .B(n4736), .Z(n2965) );
  AO7 U1818 ( .A(n4633), .B(n4288), .C(n4870), .Z(n1371) );
  ND2 U1819 ( .A(n1863), .B(n1862), .Z(n1362) );
  ND2 U1820 ( .A(n4629), .B(n4128), .Z(n1862) );
  EO U1821 ( .A(n4893), .B(n4259), .Z(n1863) );
  ND2 U1822 ( .A(n4273), .B(n4738), .Z(n2950) );
  ND2 U1823 ( .A(n4628), .B(n4821), .Z(n1903) );
  ND2 U1824 ( .A(n3053), .B(n3052), .Z(n1385) );
  ND2 U1825 ( .A(n4266), .B(n4600), .Z(n3052) );
  MUX21L U1826 ( .A(n3051), .B(n4772), .S(n4600), .Z(n3053) );
  NR2 U1827 ( .A(n4266), .B(n4772), .Z(n3051) );
  MUX21L U1828 ( .A(n4553), .B(n2258), .S(n4953), .Z(n1370) );
  ND2 U1829 ( .A(n4285), .B(n4553), .Z(n2258) );
  ND2 U1830 ( .A(n4153), .B(n4460), .Z(n924) );
  ND2 U1831 ( .A(n4955), .B(n4536), .Z(n2318) );
  ND2 U1832 ( .A(n4955), .B(n4177), .Z(n2319) );
  AN3 U1833 ( .A(n4167), .B(n4864), .C(n4569), .Z(n428) );
  ND2 U1834 ( .A(n1802), .B(n1801), .Z(n1361) );
  ND2 U1835 ( .A(n4576), .B(n4122), .Z(n1801) );
  MUX21L U1836 ( .A(n4830), .B(n1800), .S(n4263), .Z(n1802) );
  NR2 U1837 ( .A(n4576), .B(n4829), .Z(n1800) );
  MUX21L U1838 ( .A(n2746), .B(n4900), .S(n4243), .Z(n1380) );
  ND2 U1839 ( .A(n4900), .B(n4485), .Z(n2746) );
  MUX21L U1840 ( .A(n4399), .B(n4066), .S(n4945), .Z(n1375) );
  MUX21L U1841 ( .A(n4218), .B(n4482), .S(n4894), .Z(n1379) );
  ND2 U1842 ( .A(n2020), .B(n2019), .Z(n1366) );
  ND2 U1843 ( .A(n4925), .B(n4197), .Z(n2019) );
  MUX21L U1844 ( .A(n4542), .B(n2018), .S(n4297), .Z(n2020) );
  NR2 U1845 ( .A(n4926), .B(n4541), .Z(n2018) );
  MUX21L U1846 ( .A(n2358), .B(n2357), .S(n4570), .Z(n1372) );
  ND2 U1847 ( .A(n4957), .B(n4219), .Z(n2358) );
  ND2 U1848 ( .A(n4219), .B(n4867), .Z(n2357) );
  ND2 U1849 ( .A(n2107), .B(n2106), .Z(n1368) );
  ND2 U1850 ( .A(n4929), .B(n4426), .Z(n2106) );
  MUX21L U1851 ( .A(n4427), .B(n2105), .S(n4279), .Z(n2107) );
  NR2 U1852 ( .A(n4929), .B(n4426), .Z(n2105) );
  NR2 U1853 ( .A(n4604), .B(n4046), .Z(n2723) );
  NR2 U1854 ( .A(n4605), .B(n4761), .Z(n2722) );
  NR2 U1855 ( .A(n4594), .B(n4066), .Z(n2506) );
  ND2 U1856 ( .A(n2725), .B(n2724), .Z(n862) );
  MUX21L U1857 ( .A(n2721), .B(n4219), .S(n4894), .Z(n2724) );
  NR2 U1858 ( .A(n2723), .B(n2722), .Z(n2725) );
  NR2 U1859 ( .A(n4219), .B(n4482), .Z(n2721) );
  ND2 U1860 ( .A(n2025), .B(n2024), .Z(n850) );
  ND2 U1861 ( .A(n4297), .B(n4808), .Z(n2024) );
  EN U1862 ( .A(n4560), .B(n4297), .Z(n2025) );
  ND3 U1863 ( .A(n2572), .B(n2571), .C(n2570), .Z(n860) );
  ND2 U1864 ( .A(n4597), .B(n4849), .Z(n2572) );
  ND2 U1865 ( .A(n4230), .B(n4849), .Z(n2571) );
  ND2 U1866 ( .A(n4597), .B(n4230), .Z(n2570) );
  ND2 U1867 ( .A(n4607), .B(n4840), .Z(n1378) );
  ND2 U1868 ( .A(n4530), .B(n4820), .Z(n1912) );
  ND2 U1869 ( .A(n4256), .B(n4423), .Z(n2154) );
  ND2 U1870 ( .A(n4256), .B(n4797), .Z(n2156) );
  ND2 U1871 ( .A(n3020), .B(n3019), .Z(n867) );
  ND2 U1872 ( .A(n4920), .B(n4155), .Z(n3019) );
  EN U1873 ( .A(n4560), .B(n4268), .Z(n3020) );
  MUX21L U1874 ( .A(n2987), .B(n2986), .S(n4919), .Z(n866) );
  ND2 U1875 ( .A(n4611), .B(n4152), .Z(n2987) );
  ND2 U1876 ( .A(n4611), .B(n4271), .Z(n2986) );
  ND2 U1877 ( .A(n2245), .B(n2244), .Z(n854) );
  ND2 U1878 ( .A(n4185), .B(n4877), .Z(n2244) );
  EO U1879 ( .A(n4566), .B(n4284), .Z(n2245) );
  ND2 U1880 ( .A(n2347), .B(n2346), .Z(n856) );
  ND2 U1881 ( .A(n4956), .B(n4283), .Z(n2346) );
  EN U1882 ( .A(n4888), .B(n4568), .Z(n2347) );
  MUX21L U1883 ( .A(n4409), .B(n2439), .S(n4942), .Z(n858) );
  ND2 U1884 ( .A(n4223), .B(n4409), .Z(n2439) );
  ND2 U1885 ( .A(n4925), .B(n4622), .Z(n2017) );
  AN3 U1886 ( .A(n4144), .B(n4502), .C(n4915), .Z(n429) );
  ND2 U1887 ( .A(n2944), .B(n4148), .Z(n1354) );
  EN U1888 ( .A(n4888), .B(n4613), .Z(n2944) );
  IVP U1889 ( .A(n4034), .Z(n4233) );
  NR2 U1890 ( .A(n4578), .B(n4801), .Z(n2110) );
  NR2 U1891 ( .A(n4635), .B(n4874), .Z(n2283) );
  NR2 U1892 ( .A(n4635), .B(n4181), .Z(n2284) );
  ND2 U1893 ( .A(n4079), .B(n4789), .Z(n3222) );
  ND2 U1894 ( .A(n4587), .B(n4790), .Z(n3221) );
  ND2 U1895 ( .A(n4233), .B(n4444), .Z(n3148) );
  ND2 U1896 ( .A(n4233), .B(n4781), .Z(n3150) );
  ND2 U1897 ( .A(n2427), .B(n2426), .Z(n1346) );
  MUX21L U1898 ( .A(n2424), .B(n4859), .S(n4591), .Z(n2426) );
  AO6 U1899 ( .A(n4591), .B(n4160), .C(n2425), .Z(n2427) );
  ND2 U1900 ( .A(n2578), .B(n4060), .Z(n1348) );
  EO U1901 ( .A(n4891), .B(n4632), .Z(n2578) );
  MUX21L U1902 ( .A(n2481), .B(n2480), .S(n4226), .Z(n1347) );
  ND2 U1903 ( .A(n4943), .B(n4593), .Z(n2481) );
  ND2 U1904 ( .A(n4593), .B(n4855), .Z(n2480) );
  MUX21L U1905 ( .A(n4536), .B(n1975), .S(n4923), .Z(n1336) );
  ND2 U1906 ( .A(n4294), .B(n4537), .Z(n1975) );
  ND2 U1907 ( .A(n2194), .B(n2193), .Z(n1341) );
  ND2 U1908 ( .A(n4281), .B(n4881), .Z(n2193) );
  MUX21L U1909 ( .A(n2192), .B(n4881), .S(n4638), .Z(n2194) );
  NR2 U1910 ( .A(n4282), .B(n4881), .Z(n2192) );
  ND2 U1911 ( .A(n2286), .B(n2285), .Z(n1342) );
  MUX21L U1912 ( .A(n2282), .B(n4286), .S(n4954), .Z(n2285) );
  NR2 U1913 ( .A(n2284), .B(n2283), .Z(n2286) );
  NR2 U1914 ( .A(n4286), .B(n4555), .Z(n2282) );
  AN3 U1915 ( .A(n4243), .B(n4758), .C(n4604), .Z(n430) );
  MUX21L U1916 ( .A(n4093), .B(n4905), .S(n4596), .Z(n1357) );
  ND2 U1917 ( .A(n2672), .B(n2671), .Z(n1350) );
  ND2 U1918 ( .A(n4475), .B(n4765), .Z(n2671) );
  MUX21L U1919 ( .A(n4476), .B(n2670), .S(n4215), .Z(n2672) );
  ND2 U1920 ( .A(n1923), .B(n1922), .Z(n1334) );
  ND2 U1921 ( .A(n4256), .B(n4627), .Z(n1922) );
  MUX21L U1922 ( .A(n1921), .B(n4818), .S(n4627), .Z(n1923) );
  NR2 U1923 ( .A(n4256), .B(n4817), .Z(n1921) );
  ND2 U1924 ( .A(n1866), .B(n1865), .Z(n1333) );
  ND2 U1925 ( .A(n4938), .B(n4629), .Z(n1865) );
  MUX21L U1926 ( .A(n1864), .B(n4128), .S(n4629), .Z(n1866) );
  NR2 U1927 ( .A(n4938), .B(n4128), .Z(n1864) );
  ND2 U1928 ( .A(n1713), .B(n1712), .Z(n1330) );
  ND2 U1929 ( .A(n4572), .B(n4110), .Z(n1712) );
  MUX21L U1930 ( .A(n1711), .B(n4111), .S(n4933), .Z(n1713) );
  NR2 U1931 ( .A(n4572), .B(n4110), .Z(n1711) );
  ND2 U1932 ( .A(n2112), .B(n2111), .Z(n1340) );
  ND2 U1933 ( .A(n2108), .B(n4426), .Z(n2111) );
  MUX21L U1934 ( .A(n2109), .B(n2110), .S(n4279), .Z(n2112) );
  NR2 U1935 ( .A(n4929), .B(n4279), .Z(n2108) );
  NR2 U1936 ( .A(n4604), .B(n4046), .Z(n2727) );
  ND2 U1937 ( .A(n2044), .B(n2043), .Z(n1338) );
  ND2 U1938 ( .A(n4298), .B(n4805), .Z(n2043) );
  EO U1939 ( .A(n4886), .B(n4641), .Z(n2044) );
  ND3 U1940 ( .A(n4570), .B(n4220), .C(n4957), .Z(n1343) );
  ND2 U1941 ( .A(n4226), .B(n4401), .Z(n2495) );
  ND2 U1942 ( .A(n4226), .B(n4855), .Z(n2497) );
  ND2 U1943 ( .A(n2663), .B(n2662), .Z(n833) );
  ND2 U1944 ( .A(n4608), .B(n4841), .Z(n2662) );
  MUX21L U1945 ( .A(n2661), .B(n4052), .S(n4608), .Z(n2663) );
  ND2 U1946 ( .A(n2776), .B(n2775), .Z(n835) );
  ND2 U1947 ( .A(n4488), .B(n4756), .Z(n2775) );
  MUX21L U1948 ( .A(n4757), .B(n2774), .S(n4245), .Z(n2776) );
  ND2 U1949 ( .A(n3174), .B(n3173), .Z(n842) );
  ND2 U1950 ( .A(n4909), .B(n4442), .Z(n3174) );
  ND2 U1951 ( .A(n4234), .B(n4441), .Z(n3173) );
  ND2 U1952 ( .A(n2322), .B(n2321), .Z(n828) );
  ND2 U1953 ( .A(n4633), .B(n4176), .Z(n2321) );
  MUX21L U1954 ( .A(n2320), .B(n4177), .S(n4955), .Z(n2322) );
  NR2 U1955 ( .A(n4633), .B(n4176), .Z(n2320) );
  ND2 U1956 ( .A(n2061), .B(n2060), .Z(n1339) );
  ND2 U1957 ( .A(n4640), .B(n4193), .Z(n2060) );
  MUX21L U1958 ( .A(n4803), .B(n2059), .S(n4299), .Z(n2061) );
  NR2 U1959 ( .A(n4640), .B(n4803), .Z(n2059) );
  MUX21L U1960 ( .A(n3083), .B(n3082), .S(n4252), .Z(n841) );
  ND2 U1961 ( .A(n4450), .B(n4775), .Z(n3082) );
  ND2 U1962 ( .A(n4581), .B(n4774), .Z(n3083) );
  MUX21L U1963 ( .A(n2813), .B(n4899), .S(n4247), .Z(n837) );
  ND2 U1964 ( .A(n4899), .B(n4493), .Z(n2813) );
  ND2 U1965 ( .A(n1834), .B(n1833), .Z(n1301) );
  ND2 U1966 ( .A(n4261), .B(n4826), .Z(n1833) );
  EN U1967 ( .A(n4566), .B(n4261), .Z(n1834) );
  NR2 U1968 ( .A(n4211), .B(n4467), .Z(n2594) );
  NR2 U1969 ( .A(n4592), .B(n4857), .Z(n2452) );
  NR2 U1970 ( .A(n4592), .B(n4158), .Z(n2453) );
  ND2 U1971 ( .A(n1905), .B(n1904), .Z(n1302) );
  ND2 U1972 ( .A(n4939), .B(n4133), .Z(n1904) );
  EN U1973 ( .A(n4565), .B(n4258), .Z(n1905) );
  ND2 U1974 ( .A(n4061), .B(n4848), .Z(n1376) );
  ND2 U1975 ( .A(n2455), .B(n2454), .Z(n1313) );
  MUX21L U1976 ( .A(n2451), .B(n4224), .S(n4942), .Z(n2454) );
  NR2 U1977 ( .A(n2453), .B(n2452), .Z(n2455) );
  NR2 U1978 ( .A(n4224), .B(n4406), .Z(n2451) );
  ND2 U1979 ( .A(n2769), .B(n2768), .Z(n1319) );
  ND2 U1980 ( .A(n4244), .B(n4487), .Z(n2768) );
  MUX21L U1981 ( .A(n2767), .B(n4904), .S(n4244), .Z(n2769) );
  NR2 U1982 ( .A(n4903), .B(n4487), .Z(n2767) );
  ND2 U1983 ( .A(n2400), .B(n2399), .Z(n1312) );
  ND2 U1984 ( .A(n4222), .B(n4863), .Z(n2399) );
  MUX21L U1985 ( .A(n2398), .B(n4864), .S(n4569), .Z(n2400) );
  NR2 U1986 ( .A(n4222), .B(n4863), .Z(n2398) );
  ND2 U1987 ( .A(n3123), .B(n3122), .Z(n1326) );
  ND2 U1988 ( .A(n4231), .B(n4778), .Z(n3122) );
  EO U1989 ( .A(n4562), .B(n4231), .Z(n3123) );
  ND2 U1990 ( .A(n2291), .B(n2290), .Z(n1308) );
  ND2 U1991 ( .A(n2287), .B(n4954), .Z(n2290) );
  MUX21L U1992 ( .A(n2288), .B(n2289), .S(n4954), .Z(n2291) );
  NR2 U1993 ( .A(n4635), .B(n4286), .Z(n2287) );
  ND2 U1994 ( .A(n4554), .B(n4874), .Z(n2268) );
  ND2 U1995 ( .A(n4422), .B(n4797), .Z(n2155) );
  ND2 U1996 ( .A(n2142), .B(n4136), .Z(n826) );
  ND2 U1997 ( .A(n4931), .B(n4579), .Z(n2142) );
  MUX21L U1998 ( .A(n1937), .B(n4204), .S(n4922), .Z(n1939) );
  NR2 U1999 ( .A(n4626), .B(n4204), .Z(n1937) );
  AO7 U2000 ( .A(n4896), .B(n4495), .C(n4248), .Z(n1322) );
  AO7 U2001 ( .A(n4598), .B(n4153), .C(n4919), .Z(n1325) );
  AO7 U2002 ( .A(n4952), .B(n4284), .C(n4551), .Z(n1307) );
  NR2 U2003 ( .A(n4948), .B(n4059), .Z(n2592) );
  NR2 U2004 ( .A(n4635), .B(n4180), .Z(n2288) );
  NR2 U2005 ( .A(n4601), .B(n4755), .Z(n1321) );
  ND2 U2006 ( .A(n4895), .B(n4045), .Z(n2732) );
  ND2 U2007 ( .A(n4604), .B(n4895), .Z(n2733) );
  ND2 U2008 ( .A(n4604), .B(n4045), .Z(n2731) );
  ND2 U2009 ( .A(n4226), .B(n4855), .Z(n2482) );
  ND2 U2010 ( .A(n4226), .B(n4402), .Z(n2483) );
  ND2 U2011 ( .A(n4896), .B(n4473), .Z(n2653) );
  ND2 U2012 ( .A(n4958), .B(n2375), .Z(n1310) );
  ND2 U2013 ( .A(n4571), .B(n4220), .Z(n2375) );
  ND2 U2014 ( .A(n2816), .B(n2815), .Z(n813) );
  ND2 U2015 ( .A(n4247), .B(n4493), .Z(n2815) );
  MUX21L U2016 ( .A(n4898), .B(n2814), .S(n4620), .Z(n2816) );
  NR2 U2017 ( .A(n4898), .B(n4247), .Z(n2814) );
  MUX21L U2018 ( .A(n4150), .B(n4917), .S(n4613), .Z(n1324) );
  MUX21L U2019 ( .A(n2114), .B(n2113), .S(n4279), .Z(n1306) );
  ND2 U2020 ( .A(n4425), .B(n4801), .Z(n2113) );
  ND2 U2021 ( .A(n4930), .B(n4578), .Z(n2114) );
  ND2 U2022 ( .A(n2431), .B(n2430), .Z(n1281) );
  MUX21L U2023 ( .A(n2428), .B(n4859), .S(n4591), .Z(n2430) );
  AO6 U2024 ( .A(n4591), .B(n4160), .C(n2429), .Z(n2431) );
  ND2 U2025 ( .A(n2891), .B(n2890), .Z(n1291) );
  ND2 U2026 ( .A(n2887), .B(n4502), .Z(n2890) );
  MUX21L U2027 ( .A(n2888), .B(n2889), .S(n4276), .Z(n2891) );
  NR2 U2028 ( .A(n4914), .B(n4276), .Z(n2887) );
  ND2 U2029 ( .A(n4400), .B(n4854), .Z(n2496) );
  ND2 U2030 ( .A(n4408), .B(n4858), .Z(n2440) );
  ND2 U2031 ( .A(n4270), .B(n4460), .Z(n815) );
  NR2 U2032 ( .A(n4616), .B(n4743), .Z(n2889) );
  ND3 U2033 ( .A(n2626), .B(n2625), .C(n2624), .Z(n1284) );
  ND2 U2034 ( .A(n4945), .B(n4471), .Z(n2625) );
  ND2 U2035 ( .A(n4211), .B(n4949), .Z(n2626) );
  ND2 U2036 ( .A(n4213), .B(n4471), .Z(n2624) );
  ND3 U2037 ( .A(n2261), .B(n2260), .C(n2259), .Z(n1277) );
  ND2 U2038 ( .A(n4553), .B(n4876), .Z(n2260) );
  ND2 U2039 ( .A(n4285), .B(n4876), .Z(n2261) );
  ND2 U2040 ( .A(n4285), .B(n4554), .Z(n2259) );
  ND2 U2041 ( .A(n4054), .B(n4473), .Z(n2654) );
  ND2 U2042 ( .A(n4944), .B(n4402), .Z(n2484) );
  ND2 U2043 ( .A(n4944), .B(n4069), .Z(n2485) );
  ND2 U2044 ( .A(n4946), .B(n4398), .Z(n2529) );
  ND2 U2045 ( .A(n4222), .B(n4415), .Z(n2401) );
  ND2 U2046 ( .A(n4941), .B(n4415), .Z(n2402) );
  ND2 U2047 ( .A(n3002), .B(n3001), .Z(n1293) );
  ND2 U2048 ( .A(n4269), .B(n4766), .Z(n3001) );
  MUX21L U2049 ( .A(n4458), .B(n3000), .S(n4920), .Z(n3002) );
  NR2 U2050 ( .A(n4269), .B(n4458), .Z(n3000) );
  ND2 U2051 ( .A(n2344), .B(n2343), .Z(n1278) );
  ND2 U2052 ( .A(n4289), .B(n4567), .Z(n2343) );
  MUX21L U2053 ( .A(n2342), .B(n4869), .S(n4567), .Z(n2344) );
  NR2 U2054 ( .A(n4289), .B(n4868), .Z(n2342) );
  ND2 U2055 ( .A(n2141), .B(n4136), .Z(n1274) );
  ND2 U2056 ( .A(n4931), .B(n4579), .Z(n2141) );
  ND2 U2057 ( .A(n4194), .B(n4545), .Z(n824) );
  ND2 U2058 ( .A(n4179), .B(n4557), .Z(n827) );
  MUX21L U2059 ( .A(n2795), .B(n2794), .S(n4246), .Z(n1289) );
  ND2 U2060 ( .A(n4490), .B(n4754), .Z(n2794) );
  ND2 U2061 ( .A(n4601), .B(n4754), .Z(n2795) );
  MUX21L U2062 ( .A(n2953), .B(n4917), .S(n4273), .Z(n1292) );
  ND2 U2063 ( .A(n4917), .B(n4507), .Z(n2953) );
  ND2 U2064 ( .A(n4238), .B(n4792), .Z(n3234) );
  ND2 U2065 ( .A(n4620), .B(n4105), .Z(n2817) );
  ND2 U2066 ( .A(n4898), .B(n4105), .Z(n2818) );
  ND2 U2067 ( .A(n3176), .B(n3175), .Z(n797) );
  ND2 U2068 ( .A(n4909), .B(n4084), .Z(n3175) );
  EN U2069 ( .A(n4563), .B(n4234), .Z(n3176) );
  ND2 U2070 ( .A(n2843), .B(n2842), .Z(n792) );
  ND2 U2071 ( .A(n4249), .B(n4496), .Z(n2842) );
  MUX21L U2072 ( .A(n4497), .B(n2841), .S(n4895), .Z(n2843) );
  NR2 U2073 ( .A(n4249), .B(n4496), .Z(n2841) );
  ND2 U2074 ( .A(n3023), .B(n3022), .Z(n795) );
  ND2 U2075 ( .A(n4268), .B(n4768), .Z(n3022) );
  MUX21L U2076 ( .A(n4455), .B(n3021), .S(n4921), .Z(n3023) );
  NR2 U2077 ( .A(n4268), .B(n4455), .Z(n3021) );
  ND2 U2078 ( .A(n2307), .B(n2306), .Z(n1248) );
  ND2 U2079 ( .A(n4955), .B(n4178), .Z(n2306) );
  EN U2080 ( .A(n4566), .B(n4287), .Z(n2307) );
  NR2 U2081 ( .A(n4211), .B(n4468), .Z(n2600) );
  ND2 U2082 ( .A(n4568), .B(n4166), .Z(n2403) );
  ND2 U2083 ( .A(n2720), .B(n2719), .Z(n1256) );
  ND2 U2084 ( .A(n4605), .B(n4046), .Z(n2719) );
  EO U2085 ( .A(n4884), .B(n4219), .Z(n2720) );
  ND2 U2086 ( .A(n2657), .B(n2656), .Z(n1255) );
  ND2 U2087 ( .A(n4897), .B(n4474), .Z(n2656) );
  MUX21L U2088 ( .A(n2655), .B(n4053), .S(n4897), .Z(n2657) );
  ND2 U2089 ( .A(n2532), .B(n2531), .Z(n1253) );
  ND2 U2090 ( .A(n4228), .B(n4398), .Z(n2531) );
  MUX21L U2091 ( .A(n4946), .B(n2530), .S(n4596), .Z(n2532) );
  NR2 U2092 ( .A(n4946), .B(n4228), .Z(n2530) );
  ND2 U2093 ( .A(n3074), .B(n3073), .Z(n1263) );
  MUX21L U2094 ( .A(n3071), .B(n4774), .S(n4251), .Z(n3073) );
  AO6 U2095 ( .A(n4252), .B(n4451), .C(n3072), .Z(n3074) );
  ND2 U2096 ( .A(n2893), .B(n2892), .Z(n1261) );
  ND2 U2097 ( .A(n4141), .B(n4743), .Z(n2893) );
  ND2 U2098 ( .A(n4616), .B(n4742), .Z(n2892) );
  ND2 U2099 ( .A(n4179), .B(n4558), .Z(n805) );
  ND2 U2100 ( .A(n3238), .B(n3237), .Z(n781) );
  ND2 U2101 ( .A(n4588), .B(n4076), .Z(n3237) );
  MUX21L U2102 ( .A(n4792), .B(n3236), .S(n4238), .Z(n3238) );
  NR2 U2103 ( .A(n4588), .B(n4792), .Z(n3236) );
  ND2 U2104 ( .A(n2968), .B(n2967), .Z(n777) );
  ND2 U2105 ( .A(n4918), .B(n4510), .Z(n2967) );
  MUX21L U2106 ( .A(n4510), .B(n2966), .S(n4272), .Z(n2968) );
  NR2 U2107 ( .A(n4918), .B(n4509), .Z(n2966) );
  ND2 U2108 ( .A(n3118), .B(n3117), .Z(n779) );
  ND2 U2109 ( .A(n4090), .B(n4446), .Z(n3117) );
  EO U2110 ( .A(n4884), .B(n4254), .Z(n3118) );
  ND2 U2111 ( .A(n2911), .B(n2910), .Z(n776) );
  ND2 U2112 ( .A(n4276), .B(n4503), .Z(n2910) );
  MUX21L U2113 ( .A(n4276), .B(n2909), .S(n4915), .Z(n2911) );
  NR2 U2114 ( .A(n4276), .B(n4503), .Z(n2909) );
  AO7 U2115 ( .A(n4619), .B(n4753), .C(n4102), .Z(n1259) );
  NR2 U2116 ( .A(n4948), .B(n4058), .Z(n2598) );
  ND2 U2117 ( .A(n4941), .B(n4167), .Z(n2404) );
  AN3 U2118 ( .A(n4150), .B(n4508), .C(n4917), .Z(n431) );
  MUX21L U2119 ( .A(n4617), .B(n4097), .S(n4894), .Z(n1260) );
  MUX21L U2120 ( .A(n3024), .B(n4598), .S(n4268), .Z(n778) );
  ND2 U2121 ( .A(n4598), .B(n4768), .Z(n3024) );
  ND2 U2122 ( .A(n2898), .B(n2897), .Z(n1235) );
  ND2 U2123 ( .A(n2894), .B(n4502), .Z(n2897) );
  MUX21L U2124 ( .A(n2895), .B(n2896), .S(n4276), .Z(n2898) );
  NR2 U2125 ( .A(n4914), .B(n4276), .Z(n2894) );
  ND2 U2126 ( .A(n2797), .B(n2796), .Z(n1233) );
  ND2 U2127 ( .A(n4038), .B(n4490), .Z(n2796) );
  EN U2128 ( .A(n4887), .B(n4246), .Z(n2797) );
  ND2 U2129 ( .A(n2772), .B(n2771), .Z(n1231) );
  ND2 U2130 ( .A(n4244), .B(n4487), .Z(n2771) );
  EO U2131 ( .A(n4886), .B(n4244), .Z(n2772) );
  ND2 U2132 ( .A(n4077), .B(n4791), .Z(n3235) );
  NR2 U2133 ( .A(n4616), .B(n4742), .Z(n2896) );
  ND2 U2134 ( .A(n4411), .B(n4859), .Z(n2432) );
  ND2 U2135 ( .A(n3101), .B(n3100), .Z(n1237) );
  ND2 U2136 ( .A(n4253), .B(n4447), .Z(n3100) );
  EO U2137 ( .A(n4884), .B(n4253), .Z(n3101) );
  ND2 U2138 ( .A(n3210), .B(n4080), .Z(n1238) );
  ND2 U2139 ( .A(n4910), .B(n4587), .Z(n3210) );
  ND2 U2140 ( .A(n2488), .B(n2487), .Z(n1226) );
  ND2 U2141 ( .A(n4593), .B(n4069), .Z(n2487) );
  MUX21L U2142 ( .A(n2486), .B(n4069), .S(n4944), .Z(n2488) );
  NR2 U2143 ( .A(n4593), .B(n4068), .Z(n2486) );
  ND2 U2144 ( .A(n2534), .B(n2533), .Z(n1227) );
  ND2 U2145 ( .A(n4947), .B(n4064), .Z(n2534) );
  ND2 U2146 ( .A(n4596), .B(n4063), .Z(n2533) );
  AN3 U2147 ( .A(n4273), .B(n4508), .C(n4917), .Z(n432) );
  MUX21L U2148 ( .A(n4479), .B(n2706), .S(n4900), .Z(n1230) );
  ND2 U2149 ( .A(n4217), .B(n4480), .Z(n2706) );
  MUX21L U2150 ( .A(n2604), .B(n2603), .S(n4211), .Z(n1228) );
  ND2 U2151 ( .A(n4468), .B(n4847), .Z(n2603) );
  ND2 U2152 ( .A(n4948), .B(n4611), .Z(n2604) );
  ND2 U2153 ( .A(n2945), .B(n4148), .Z(n767) );
  ND2 U2154 ( .A(n4917), .B(n4613), .Z(n2945) );
  ND2 U2155 ( .A(n2800), .B(n2799), .Z(n1212) );
  ND2 U2156 ( .A(n4246), .B(n4490), .Z(n2799) );
  MUX21L U2157 ( .A(n4901), .B(n2798), .S(n4601), .Z(n2800) );
  NR2 U2158 ( .A(n4900), .B(n4246), .Z(n2798) );
  ND2 U2159 ( .A(n3283), .B(n3282), .Z(n1219) );
  ND2 U2160 ( .A(n4241), .B(n4795), .Z(n3282) );
  EO U2161 ( .A(n4890), .B(n4590), .Z(n3283) );
  ND2 U2162 ( .A(n2862), .B(n2861), .Z(n1213) );
  ND2 U2163 ( .A(n4498), .B(n4747), .Z(n2861) );
  MUX21L U2164 ( .A(n4747), .B(n2860), .S(n4250), .Z(n2862) );
  ND2 U2165 ( .A(n3087), .B(n3086), .Z(n770) );
  MUX21L U2166 ( .A(n3084), .B(n4775), .S(n4581), .Z(n3086) );
  AO6 U2167 ( .A(n4581), .B(n4091), .C(n3085), .Z(n3087) );
  ND2 U2168 ( .A(n2641), .B(n4056), .Z(n1209) );
  ND2 U2169 ( .A(n4895), .B(n4609), .Z(n2641) );
  ND2 U2170 ( .A(n2660), .B(n2659), .Z(n1210) );
  ND2 U2171 ( .A(n4608), .B(n4053), .Z(n2659) );
  MUX21L U2172 ( .A(n2658), .B(n4053), .S(n4897), .Z(n2660) );
  NR2 U2173 ( .A(n4608), .B(n4052), .Z(n2658) );
  ND2 U2174 ( .A(n4458), .B(n4767), .Z(n3003) );
  ND2 U2175 ( .A(n4909), .B(n4084), .Z(n3178) );
  MUX21L U2176 ( .A(n2955), .B(n2954), .S(n4273), .Z(n1215) );
  ND2 U2177 ( .A(n4508), .B(n4738), .Z(n2954) );
  ND2 U2178 ( .A(n4612), .B(n4738), .Z(n2955) );
  MUX21L U2179 ( .A(n4093), .B(n4905), .S(n4581), .Z(n1217) );
  MUX21L U2180 ( .A(n4269), .B(n3004), .S(n4920), .Z(n1216) );
  ND2 U2181 ( .A(n4269), .B(n4457), .Z(n3004) );
  NR2 U2182 ( .A(n4914), .B(n4142), .Z(n2899) );
  ND2 U2183 ( .A(n2979), .B(n2978), .Z(n1198) );
  ND2 U2184 ( .A(n4151), .B(n4511), .Z(n2978) );
  EO U2185 ( .A(n4887), .B(n4271), .Z(n2979) );
  ND2 U2186 ( .A(n2902), .B(n2901), .Z(n1197) );
  AO6 U2187 ( .A(n4914), .B(n4142), .C(n2900), .Z(n2902) );
  MUX21L U2188 ( .A(n4914), .B(n2899), .S(n4616), .Z(n2901) );
  NR2 U2189 ( .A(n4616), .B(n4276), .Z(n2900) );
  ND2 U2190 ( .A(n4071), .B(n4404), .Z(n1225) );
  IVP U2191 ( .A(n4730), .Z(n4906) );
  NR2 U2192 ( .A(n4582), .B(n4091), .Z(n3102) );
  ND2 U2193 ( .A(n3107), .B(n3106), .Z(n1200) );
  MUX21L U2194 ( .A(n3104), .B(n3105), .S(n4582), .Z(n3106) );
  MUX21L U2195 ( .A(n3102), .B(n3103), .S(n4906), .Z(n3107) );
  NR2 U2196 ( .A(n4253), .B(n4776), .Z(n3104) );
  ND2 U2197 ( .A(n2802), .B(n2801), .Z(n1195) );
  ND2 U2198 ( .A(n4900), .B(n4089), .Z(n2802) );
  ND2 U2199 ( .A(n4601), .B(n4106), .Z(n2801) );
  MUX21L U2200 ( .A(n4793), .B(n3239), .S(n4238), .Z(n3241) );
  NR2 U2201 ( .A(n4588), .B(n4793), .Z(n3239) );
  ND2 U2202 ( .A(n2959), .B(n2958), .Z(n1185) );
  MUX21L U2203 ( .A(n2956), .B(n4737), .S(n4612), .Z(n2958) );
  AO6 U2204 ( .A(n4612), .B(n4150), .C(n2957), .Z(n2959) );
  ND2 U2205 ( .A(n3159), .B(n3158), .Z(n1188) );
  MUX21L U2206 ( .A(n4908), .B(n3156), .S(n4584), .Z(n3158) );
  AO6 U2207 ( .A(n4908), .B(n4087), .C(n3157), .Z(n3159) );
  NR2 U2208 ( .A(n4908), .B(n4087), .Z(n3156) );
  ND2 U2209 ( .A(n4588), .B(n4793), .Z(n3240) );
  MUX21L U2210 ( .A(n4434), .B(n3242), .S(n4912), .Z(n3244) );
  NR2 U2211 ( .A(n4239), .B(n4434), .Z(n3242) );
  ND3 U2212 ( .A(n4240), .B(n4795), .C(n4590), .Z(n1189) );
  ND2 U2213 ( .A(n4086), .B(n4443), .Z(n3161) );
  ND2 U2214 ( .A(n4584), .B(n4086), .Z(n3160) );
  ND2 U2215 ( .A(n3196), .B(n3195), .Z(n1171) );
  ND2 U2216 ( .A(n4235), .B(n4586), .Z(n3195) );
  MUX21L U2217 ( .A(n3194), .B(n4786), .S(n4586), .Z(n3196) );
  NR2 U2218 ( .A(n4236), .B(n4787), .Z(n3194) );
  ND2 U2219 ( .A(n3112), .B(n3111), .Z(n1170) );
  MUX21L U2220 ( .A(n4447), .B(n3108), .S(n4906), .Z(n3111) );
  NR2 U2221 ( .A(n3110), .B(n3109), .Z(n3112) );
  ND2 U2222 ( .A(n4456), .B(n4767), .Z(n3006) );
  ND2 U2223 ( .A(n3164), .B(n3163), .Z(n1166) );
  ND2 U2224 ( .A(n4233), .B(n4443), .Z(n3163) );
  MUX21L U2225 ( .A(n4233), .B(n3162), .S(n4908), .Z(n3164) );
  NR2 U2226 ( .A(n4233), .B(n4442), .Z(n3162) );
  ND2 U2227 ( .A(n4588), .B(n4076), .Z(n3245) );
  ND2 U2228 ( .A(n4078), .B(n4437), .Z(n3225) );
  ND2 U2229 ( .A(n4237), .B(n4437), .Z(n3224) );
  ND2 U2230 ( .A(n3267), .B(n3266), .Z(n1162) );
  NR2 U2231 ( .A(n3265), .B(n3264), .Z(n3267) );
  MUX21L U2232 ( .A(n4432), .B(n3263), .S(n4913), .Z(n3266) );
  NR2 U2233 ( .A(n4913), .B(n4240), .Z(n3265) );
  NR2 U2234 ( .A(n4623), .B(n4199), .Z(n1993) );
  NR2 U2235 ( .A(n4296), .B(n4810), .Z(n1995) );
  NR2 U2236 ( .A(n4589), .B(n4795), .Z(n3254) );
  OR3 U2237 ( .A(n4220), .B(n4958), .C(n4571), .Z(n433) );
  ND2 U2238 ( .A(n3252), .B(n4432), .Z(n3255) );
  MUX21L U2239 ( .A(n3253), .B(n3254), .S(n4239), .Z(n3256) );
  AO6 U2240 ( .A(n4264), .B(n4515), .C(n1766), .Z(n1768) );
  NR2 U2241 ( .A(n4935), .B(n4574), .Z(n1766) );
  ND2 U2242 ( .A(n3028), .B(n3027), .Z(n746) );
  MUX21L U2243 ( .A(n3025), .B(n4769), .S(n4599), .Z(n3027) );
  AO6 U2244 ( .A(n4599), .B(n4155), .C(n3026), .Z(n3028) );
  NR2 U2245 ( .A(n4629), .B(n4129), .Z(n1876) );
  NR2 U2246 ( .A(n4904), .B(n4042), .Z(n2758) );
  NR2 U2247 ( .A(n4617), .B(n4096), .Z(n2871) );
  NR2 U2248 ( .A(n4296), .B(n4540), .Z(n2002) );
  NR2 U2249 ( .A(n4622), .B(n4810), .Z(n2003) );
  NR2 U2250 ( .A(n4930), .B(n4190), .Z(n2122) );
  NR2 U2251 ( .A(n4950), .B(n4139), .Z(n2161) );
  NR2 U2252 ( .A(n4928), .B(n4546), .Z(n2066) );
  NR2 U2253 ( .A(n4230), .B(n4461), .Z(n2565) );
  NR2 U2254 ( .A(n4597), .B(n4849), .Z(n2566) );
  NR2 U2255 ( .A(n4251), .B(n4745), .Z(n2876) );
  NR2 U2256 ( .A(n4913), .B(n4500), .Z(n2877) );
  NR2 U2257 ( .A(n4582), .B(n4775), .Z(n3094) );
  ND2 U2258 ( .A(n4925), .B(n4539), .Z(n2000) );
  ND2 U2259 ( .A(n4296), .B(n4925), .Z(n2001) );
  ND2 U2260 ( .A(n4296), .B(n4539), .Z(n1999) );
  ND2 U2261 ( .A(n3185), .B(n3184), .Z(n688) );
  ND2 U2262 ( .A(n4235), .B(n4440), .Z(n3184) );
  EN U2263 ( .A(n4892), .B(n4585), .Z(n3185) );
  ND2 U2264 ( .A(n1963), .B(n1962), .Z(n601) );
  ND2 U2265 ( .A(n4203), .B(n4813), .Z(n1962) );
  EO U2266 ( .A(n4563), .B(n4293), .Z(n1963) );
  ND2 U2267 ( .A(n2349), .B(n2348), .Z(n610) );
  ND2 U2268 ( .A(n4956), .B(n4277), .Z(n2348) );
  EN U2269 ( .A(n4888), .B(n4569), .Z(n2349) );
  ND2 U2270 ( .A(n3297), .B(n4073), .Z(n594) );
  EO U2271 ( .A(n4890), .B(n4586), .Z(n3297) );
  ND2 U2272 ( .A(n4255), .B(n4422), .Z(n2159) );
  ND2 U2273 ( .A(n2212), .B(n4879), .Z(n2215) );
  NR2 U2274 ( .A(n4282), .B(n4638), .Z(n2212) );
  ND2 U2275 ( .A(n4938), .B(n4129), .Z(n1881) );
  ND2 U2276 ( .A(n4629), .B(n4130), .Z(n1880) );
  ND2 U2277 ( .A(n4952), .B(n4186), .Z(n2237) );
  ND2 U2278 ( .A(n2158), .B(n2157), .Z(n729) );
  ND2 U2279 ( .A(n4255), .B(n4797), .Z(n2157) );
  EN U2280 ( .A(n4560), .B(n4255), .Z(n2158) );
  ND2 U2281 ( .A(n2211), .B(n2210), .Z(n730) );
  ND2 U2282 ( .A(n4638), .B(n4879), .Z(n2210) );
  MUX21L U2283 ( .A(n2209), .B(n4187), .S(n4638), .Z(n2211) );
  ND2 U2284 ( .A(n2079), .B(n2078), .Z(n727) );
  ND2 U2285 ( .A(n4192), .B(n4802), .Z(n2078) );
  EO U2286 ( .A(n4563), .B(n4277), .Z(n2079) );
  ND2 U2287 ( .A(n2760), .B(n2759), .Z(n740) );
  ND3 U2288 ( .A(n4603), .B(n4042), .C(n4898), .Z(n2759) );
  MUX21L U2289 ( .A(n2757), .B(n2758), .S(n4603), .Z(n2760) );
  ND2 U2290 ( .A(n2694), .B(n4050), .Z(n739) );
  EO U2291 ( .A(n4893), .B(n4606), .Z(n2694) );
  ND2 U2292 ( .A(n3279), .B(n3278), .Z(n749) );
  MUX21L U2293 ( .A(n4431), .B(n3275), .S(n4913), .Z(n3278) );
  NR2 U2294 ( .A(n3277), .B(n3276), .Z(n3279) );
  ND2 U2295 ( .A(n3057), .B(n3056), .Z(n716) );
  ND2 U2296 ( .A(n4157), .B(n4773), .Z(n3056) );
  EO U2297 ( .A(n4561), .B(n4266), .Z(n3057) );
  ND2 U2298 ( .A(n2869), .B(n4745), .Z(n713) );
  EN U2299 ( .A(n4564), .B(n4251), .Z(n2869) );
  ND2 U2300 ( .A(n2512), .B(n2511), .Z(n705) );
  ND2 U2301 ( .A(n4227), .B(n4400), .Z(n2511) );
  EO U2302 ( .A(n4892), .B(n4227), .Z(n2512) );
  ND2 U2303 ( .A(n1818), .B(n1817), .Z(n661) );
  ND2 U2304 ( .A(n4428), .B(n4827), .Z(n1817) );
  MUX21L U2305 ( .A(n4827), .B(n1816), .S(n4262), .Z(n1818) );
  ND2 U2306 ( .A(n2971), .B(n2970), .Z(n685) );
  ND2 U2307 ( .A(n4612), .B(n4735), .Z(n2970) );
  MUX21L U2308 ( .A(n2969), .B(n4151), .S(n4612), .Z(n2971) );
  ND2 U2309 ( .A(n2564), .B(n2563), .Z(n676) );
  ND2 U2310 ( .A(n4461), .B(n4850), .Z(n2563) );
  MUX21L U2311 ( .A(n4461), .B(n2562), .S(n4230), .Z(n2564) );
  ND2 U2312 ( .A(n2736), .B(n2735), .Z(n679) );
  ND2 U2313 ( .A(n4483), .B(n4760), .Z(n2735) );
  MUX21L U2314 ( .A(n4483), .B(n2734), .S(n4219), .Z(n2736) );
  ND2 U2315 ( .A(n2616), .B(n2615), .Z(n677) );
  ND2 U2316 ( .A(n4949), .B(n4470), .Z(n2615) );
  MUX21L U2317 ( .A(n2614), .B(n4058), .S(n4949), .Z(n2616) );
  ND2 U2318 ( .A(n2462), .B(n2461), .Z(n644) );
  ND2 U2319 ( .A(n4592), .B(n4055), .Z(n2461) );
  EO U2320 ( .A(n4885), .B(n4224), .Z(n2462) );
  ND2 U2321 ( .A(n2681), .B(n2680), .Z(n648) );
  ND2 U2322 ( .A(n4903), .B(n4607), .Z(n2680) );
  MUX21L U2323 ( .A(n2679), .B(n4051), .S(n4607), .Z(n2681) );
  NR2 U2324 ( .A(n4903), .B(n4051), .Z(n2679) );
  ND2 U2325 ( .A(n1950), .B(n1949), .Z(n633) );
  MUX21L U2326 ( .A(n1947), .B(n1948), .S(n4292), .Z(n1950) );
  ND2 U2327 ( .A(n1946), .B(n4815), .Z(n1949) );
  NR2 U2328 ( .A(n4923), .B(n4535), .Z(n1948) );
  ND2 U2329 ( .A(n2164), .B(n2163), .Z(n639) );
  AO6 U2330 ( .A(n4950), .B(n4139), .C(n2162), .Z(n2164) );
  MUX21L U2331 ( .A(n4950), .B(n2161), .S(n4580), .Z(n2163) );
  NR2 U2332 ( .A(n4580), .B(n4255), .Z(n2162) );
  ND2 U2333 ( .A(n2296), .B(n2295), .Z(n641) );
  ND2 U2334 ( .A(n4556), .B(n4873), .Z(n2295) );
  MUX21L U2335 ( .A(n4873), .B(n2294), .S(n4287), .Z(n2296) );
  ND2 U2336 ( .A(n2081), .B(n2080), .Z(n605) );
  ND2 U2337 ( .A(n4192), .B(n4802), .Z(n2080) );
  EO U2338 ( .A(n4562), .B(n4278), .Z(n2081) );
  ND2 U2339 ( .A(n2880), .B(n2879), .Z(n621) );
  NR2 U2340 ( .A(n2878), .B(n2877), .Z(n2880) );
  MUX21L U2341 ( .A(n2876), .B(n4251), .S(n4616), .Z(n2879) );
  NR2 U2342 ( .A(n4913), .B(n4096), .Z(n2878) );
  ND2 U2343 ( .A(n2668), .B(n2667), .Z(n584) );
  ND2 U2344 ( .A(n4215), .B(n4475), .Z(n2667) );
  MUX21L U2345 ( .A(n4475), .B(n2666), .S(n4899), .Z(n2668) );
  NR2 U2346 ( .A(n4215), .B(n4474), .Z(n2666) );
  ND2 U2347 ( .A(n3201), .B(n3200), .Z(n593) );
  ND2 U2348 ( .A(n4910), .B(n4081), .Z(n3200) );
  EO U2349 ( .A(n4564), .B(n4236), .Z(n3201) );
  ND2 U2350 ( .A(n2270), .B(n2269), .Z(n575) );
  ND2 U2351 ( .A(n4286), .B(n4874), .Z(n2269) );
  EN U2352 ( .A(n4564), .B(n4286), .Z(n2270) );
  ND2 U2353 ( .A(n2329), .B(n2328), .Z(n576) );
  ND2 U2354 ( .A(n4633), .B(n4175), .Z(n2328) );
  MUX21L U2355 ( .A(n2327), .B(n4175), .S(n4956), .Z(n2329) );
  NR2 U2356 ( .A(n4633), .B(n4175), .Z(n2327) );
  ND2 U2357 ( .A(n2370), .B(n2369), .Z(n577) );
  ND2 U2358 ( .A(n4571), .B(n4169), .Z(n2369) );
  MUX21L U2359 ( .A(n2368), .B(n4170), .S(n4958), .Z(n2370) );
  NR2 U2360 ( .A(n4571), .B(n4169), .Z(n2368) );
  ND2 U2361 ( .A(n2914), .B(n2913), .Z(n558) );
  ND2 U2362 ( .A(n4915), .B(n4504), .Z(n2913) );
  MUX21L U2363 ( .A(n4504), .B(n2912), .S(n4275), .Z(n2914) );
  NR2 U2364 ( .A(n4915), .B(n4504), .Z(n2912) );
  ND2 U2365 ( .A(n3096), .B(n3095), .Z(n561) );
  ND2 U2366 ( .A(n3092), .B(n4448), .Z(n3095) );
  MUX21L U2367 ( .A(n3093), .B(n3094), .S(n4252), .Z(n3096) );
  NR2 U2368 ( .A(n4906), .B(n4253), .Z(n3092) );
  ND2 U2369 ( .A(n2715), .B(n2714), .Z(n553) );
  ND2 U2370 ( .A(n4895), .B(n4047), .Z(n2714) );
  EN U2371 ( .A(n4560), .B(n4218), .Z(n2715) );
  ND2 U2372 ( .A(n4198), .B(n4540), .Z(n2011) );
  ND2 U2373 ( .A(n4622), .B(n4296), .Z(n2010) );
  MUX21L U2374 ( .A(n1765), .B(n4831), .S(n4265), .Z(n1767) );
  MUX21L U2375 ( .A(n2213), .B(n2214), .S(n4282), .Z(n2216) );
  NR2 U2376 ( .A(n4952), .B(n4548), .Z(n2214) );
  ND2 U2377 ( .A(n2443), .B(n2442), .Z(n735) );
  ND2 U2378 ( .A(n4942), .B(n4408), .Z(n2442) );
  MUX21L U2379 ( .A(n2441), .B(n4159), .S(n4942), .Z(n2443) );
  ND2 U2380 ( .A(n1725), .B(n1724), .Z(n660) );
  ND2 U2381 ( .A(n4290), .B(n4835), .Z(n1724) );
  MUX21L U2382 ( .A(n1723), .B(n4835), .S(n4572), .Z(n1725) );
  NR2 U2383 ( .A(n4290), .B(n4834), .Z(n1723) );
  ND2 U2384 ( .A(n1961), .B(n1960), .Z(n664) );
  ND2 U2385 ( .A(n4625), .B(n4293), .Z(n1960) );
  MUX21L U2386 ( .A(n1959), .B(n4814), .S(n4293), .Z(n1961) );
  NR2 U2387 ( .A(n4625), .B(n4814), .Z(n1959) );
  ND2 U2388 ( .A(n2006), .B(n2005), .Z(n634) );
  NR2 U2389 ( .A(n2004), .B(n2003), .Z(n2006) );
  MUX21L U2390 ( .A(n2002), .B(n4296), .S(n4925), .Z(n2005) );
  NR2 U2391 ( .A(n4622), .B(n4199), .Z(n2004) );
  ND2 U2392 ( .A(n1918), .B(n1917), .Z(n632) );
  ND2 U2393 ( .A(n4257), .B(n4532), .Z(n1917) );
  MUX21L U2394 ( .A(n4940), .B(n1916), .S(n4627), .Z(n1918) );
  NR2 U2395 ( .A(n4940), .B(n4257), .Z(n1916) );
  ND2 U2396 ( .A(n2326), .B(n2325), .Z(n642) );
  ND2 U2397 ( .A(n4956), .B(n4465), .Z(n2325) );
  MUX21L U2398 ( .A(n2324), .B(n4176), .S(n4956), .Z(n2326) );
  ND2 U2399 ( .A(n2068), .B(n2067), .Z(n637) );
  ND2 U2400 ( .A(n2064), .B(n4802), .Z(n2067) );
  MUX21L U2401 ( .A(n2065), .B(n2066), .S(n4300), .Z(n2068) );
  NR2 U2402 ( .A(n4300), .B(n4639), .Z(n2064) );
  ND2 U2403 ( .A(n1851), .B(n1850), .Z(n599) );
  ND2 U2404 ( .A(n4260), .B(n4526), .Z(n1850) );
  MUX21L U2405 ( .A(n4260), .B(n1849), .S(n4938), .Z(n1851) );
  NR2 U2406 ( .A(n4260), .B(n4526), .Z(n1849) );
  ND2 U2407 ( .A(n1771), .B(n1770), .Z(n597) );
  ND2 U2408 ( .A(n4575), .B(n4119), .Z(n1770) );
  MUX21L U2409 ( .A(n1769), .B(n4119), .S(n4935), .Z(n1771) );
  NR2 U2410 ( .A(n4575), .B(n4119), .Z(n1769) );
  ND2 U2411 ( .A(n2219), .B(n2218), .Z(n608) );
  ND2 U2412 ( .A(n4283), .B(n4549), .Z(n2218) );
  MUX21L U2413 ( .A(n4549), .B(n2217), .S(n4952), .Z(n2219) );
  NR2 U2414 ( .A(n4283), .B(n4548), .Z(n2217) );
  ND2 U2415 ( .A(n2569), .B(n2568), .Z(n616) );
  NR2 U2416 ( .A(n2567), .B(n2566), .Z(n2569) );
  MUX21L U2417 ( .A(n2565), .B(n4230), .S(n4948), .Z(n2568) );
  NR2 U2418 ( .A(n4597), .B(n4061), .Z(n2567) );
  ND2 U2419 ( .A(n2713), .B(n2712), .Z(n619) );
  ND2 U2420 ( .A(n4218), .B(n4762), .Z(n2712) );
  MUX21L U2421 ( .A(n2711), .B(n4762), .S(n4605), .Z(n2713) );
  NR2 U2422 ( .A(n4218), .B(n4761), .Z(n2711) );
  ND2 U2423 ( .A(n2633), .B(n2632), .Z(n583) );
  ND2 U2424 ( .A(n4213), .B(n4609), .Z(n2632) );
  MUX21L U2425 ( .A(n2631), .B(n4844), .S(n4609), .Z(n2633) );
  NR2 U2426 ( .A(n4212), .B(n4844), .Z(n2631) );
  ND2 U2427 ( .A(n2415), .B(n2414), .Z(n579) );
  ND2 U2428 ( .A(n4567), .B(n4163), .Z(n2414) );
  MUX21L U2429 ( .A(n2413), .B(n4164), .S(n4941), .Z(n2415) );
  NR2 U2430 ( .A(n4568), .B(n4163), .Z(n2413) );
  ND2 U2431 ( .A(n3091), .B(n3090), .Z(n592) );
  ND2 U2432 ( .A(n4906), .B(n4449), .Z(n3090) );
  MUX21L U2433 ( .A(n4449), .B(n3089), .S(n4252), .Z(n3091) );
  NR2 U2434 ( .A(n4906), .B(n4449), .Z(n3089) );
  ND2 U2435 ( .A(n3188), .B(n3187), .Z(n562) );
  ND2 U2436 ( .A(n4585), .B(n4785), .Z(n3187) );
  MUX21L U2437 ( .A(n3186), .B(n4083), .S(n4585), .Z(n3188) );
  ND2 U2438 ( .A(n2823), .B(n2822), .Z(n556) );
  ND2 U2439 ( .A(n4620), .B(n4103), .Z(n2822) );
  MUX21L U2440 ( .A(n2821), .B(n4104), .S(n4897), .Z(n2823) );
  NR2 U2441 ( .A(n4620), .B(n4103), .Z(n2821) );
  ND2 U2442 ( .A(n2763), .B(n2762), .Z(n554) );
  ND2 U2443 ( .A(n4602), .B(n4041), .Z(n2762) );
  MUX21L U2444 ( .A(n2761), .B(n4041), .S(n4904), .Z(n2763) );
  NR2 U2445 ( .A(n4602), .B(n4040), .Z(n2761) );
  ND2 U2446 ( .A(n3036), .B(n3035), .Z(n535) );
  ND2 U2447 ( .A(n4267), .B(n4454), .Z(n3035) );
  MUX21L U2448 ( .A(n4267), .B(n3034), .S(n4921), .Z(n3036) );
  NR2 U2449 ( .A(n4267), .B(n4453), .Z(n3034) );
  ND2 U2450 ( .A(n2974), .B(n2973), .Z(n534) );
  ND2 U2451 ( .A(n4272), .B(n4511), .Z(n2973) );
  MUX21L U2452 ( .A(n4272), .B(n2972), .S(n4918), .Z(n2974) );
  NR2 U2453 ( .A(n4272), .B(n4510), .Z(n2972) );
  ND2 U2454 ( .A(n2028), .B(n2027), .Z(n698) );
  ND2 U2455 ( .A(n4926), .B(n4196), .Z(n2027) );
  MUX21L U2456 ( .A(n4542), .B(n2026), .S(n4297), .Z(n2028) );
  NR2 U2457 ( .A(n4926), .B(n4542), .Z(n2026) );
  ND2 U2458 ( .A(n2032), .B(n2031), .Z(n667) );
  MUX21L U2459 ( .A(n2029), .B(n4808), .S(n4641), .Z(n2031) );
  AO6 U2460 ( .A(n4641), .B(n4196), .C(n2030), .Z(n2032) );
  AO7 U2461 ( .A(n4602), .B(n4039), .C(n2777), .Z(n710) );
  ND2 U2462 ( .A(n4902), .B(n4245), .Z(n2777) );
  AO7 U2463 ( .A(n4254), .B(n4777), .C(n3119), .Z(n687) );
  ND2 U2464 ( .A(n4904), .B(n4582), .Z(n3119) );
  AO7 U2465 ( .A(n4239), .B(n4433), .C(n4912), .Z(n689) );
  AO7 U2466 ( .A(n4944), .B(n4067), .C(n4594), .Z(n675) );
  AO7 U2467 ( .A(n4611), .B(n4152), .C(n2990), .Z(n654) );
  ND2 U2468 ( .A(n4919), .B(n4270), .Z(n2990) );
  AO7 U2469 ( .A(n4287), .B(n4556), .C(n2297), .Z(n609) );
  ND2 U2470 ( .A(n4954), .B(n4634), .Z(n2297) );
  AO7 U2471 ( .A(n4910), .B(n4081), .C(n3199), .Z(n625) );
  ND2 U2472 ( .A(n4586), .B(n4236), .Z(n3199) );
  AO7 U2473 ( .A(n4243), .B(n4759), .C(n4484), .Z(n585) );
  AO7 U2474 ( .A(n4599), .B(n4266), .C(n4771), .Z(n591) );
  NR2 U2475 ( .A(n4280), .B(n4425), .Z(n2124) );
  NR2 U2476 ( .A(n4618), .B(n4750), .Z(n743) );
  ND2 U2477 ( .A(n2046), .B(n2045), .Z(n726) );
  ND2 U2478 ( .A(n4299), .B(n4805), .Z(n2045) );
  EO U2479 ( .A(n4886), .B(n4641), .Z(n2046) );
  ND3 U2480 ( .A(n3127), .B(n3126), .C(n3125), .Z(n717) );
  ND2 U2481 ( .A(n4582), .B(n4778), .Z(n3127) );
  ND2 U2482 ( .A(n4231), .B(n4778), .Z(n3126) );
  ND2 U2483 ( .A(n4582), .B(n4231), .Z(n3125) );
  ND3 U2484 ( .A(n4088), .B(n4779), .C(n4583), .Z(n656) );
  ND3 U2485 ( .A(n2550), .B(n2549), .C(n2548), .Z(n582) );
  ND2 U2486 ( .A(n4463), .B(n4850), .Z(n2549) );
  ND2 U2487 ( .A(n4229), .B(n4851), .Z(n2550) );
  ND2 U2488 ( .A(n4229), .B(n4463), .Z(n2548) );
  ND2 U2489 ( .A(n2076), .B(n2075), .Z(n668) );
  ND2 U2490 ( .A(n4192), .B(n4547), .Z(n2075) );
  EO U2491 ( .A(n4887), .B(n4639), .Z(n2076) );
  ND2 U2492 ( .A(n4610), .B(n4845), .Z(n2617) );
  ND2 U2493 ( .A(n4610), .B(n4057), .Z(n2618) );
  ND2 U2494 ( .A(n4622), .B(n4199), .Z(n2007) );
  ND2 U2495 ( .A(n4925), .B(n4198), .Z(n2008) );
  ND2 U2496 ( .A(n4572), .B(n4113), .Z(n1728) );
  ND2 U2497 ( .A(n4933), .B(n4113), .Z(n1729) );
  ND2 U2498 ( .A(n2379), .B(n2378), .Z(n732) );
  ND2 U2499 ( .A(n4958), .B(n4221), .Z(n2379) );
  ND2 U2500 ( .A(n4570), .B(n4221), .Z(n2378) );
  ND2 U2501 ( .A(n4632), .B(n4061), .Z(n737) );
  ND2 U2502 ( .A(n2695), .B(n4049), .Z(n708) );
  ND2 U2503 ( .A(n4903), .B(n4606), .Z(n2695) );
  ND3 U2504 ( .A(n1848), .B(n1847), .C(n1846), .Z(n662) );
  ND2 U2505 ( .A(n4127), .B(n4525), .Z(n1847) );
  ND2 U2506 ( .A(n4937), .B(n4525), .Z(n1848) );
  ND2 U2507 ( .A(n4937), .B(n4127), .Z(n1846) );
  ND3 U2508 ( .A(n2931), .B(n2930), .C(n2929), .Z(n684) );
  ND2 U2509 ( .A(n4916), .B(n4145), .Z(n2930) );
  ND2 U2510 ( .A(n4614), .B(n4916), .Z(n2931) );
  ND2 U2511 ( .A(n4614), .B(n4146), .Z(n2929) );
  ND2 U2512 ( .A(n2835), .B(n4101), .Z(n682) );
  ND2 U2513 ( .A(n4895), .B(n4619), .Z(n2835) );
  ND2 U2514 ( .A(n2470), .B(n4072), .Z(n674) );
  ND2 U2515 ( .A(n4943), .B(n4593), .Z(n2470) );
  ND2 U2516 ( .A(n1727), .B(n1726), .Z(n628) );
  ND2 U2517 ( .A(n4933), .B(n4520), .Z(n1727) );
  ND2 U2518 ( .A(n4290), .B(n4519), .Z(n1726) );
  ND2 U2519 ( .A(n1811), .B(n1810), .Z(n630) );
  ND2 U2520 ( .A(n4576), .B(n4123), .Z(n1811) );
  ND2 U2521 ( .A(n4576), .B(n4828), .Z(n1810) );
  ND3 U2522 ( .A(n3249), .B(n3248), .C(n3247), .Z(n626) );
  ND2 U2523 ( .A(n4075), .B(n4794), .Z(n3248) );
  ND2 U2524 ( .A(n4589), .B(n4794), .Z(n3249) );
  ND2 U2525 ( .A(n4589), .B(n4075), .Z(n3247) );
  ND3 U2526 ( .A(n2846), .B(n2845), .C(n2844), .Z(n589) );
  ND2 U2527 ( .A(n4098), .B(n4749), .Z(n2845) );
  ND2 U2528 ( .A(n4618), .B(n4749), .Z(n2846) );
  ND2 U2529 ( .A(n4618), .B(n4098), .Z(n2844) );
  ND2 U2530 ( .A(n2049), .B(n4194), .Z(n570) );
  ND2 U2531 ( .A(n4927), .B(n4640), .Z(n2049) );
  ND2 U2532 ( .A(n2248), .B(n4185), .Z(n574) );
  ND2 U2533 ( .A(n4953), .B(n4636), .Z(n2248) );
  ND2 U2534 ( .A(n3251), .B(n3250), .Z(n563) );
  ND2 U2535 ( .A(n4075), .B(n4433), .Z(n3251) );
  ND2 U2536 ( .A(n4912), .B(n4433), .Z(n3250) );
  ND2 U2537 ( .A(n2696), .B(n4049), .Z(n552) );
  ND2 U2538 ( .A(n4903), .B(n4606), .Z(n2696) );
  ND2 U2539 ( .A(n2518), .B(n4066), .Z(n550) );
  ND2 U2540 ( .A(n4945), .B(n4595), .Z(n2518) );
  AN3 U2541 ( .A(n4481), .B(n4762), .C(n4218), .Z(n434) );
  MUX21L U2542 ( .A(n1913), .B(n4940), .S(n4257), .Z(n724) );
  ND2 U2543 ( .A(n4939), .B(n4531), .Z(n1913) );
  MUX21L U2544 ( .A(n2340), .B(n4173), .S(n4956), .Z(n731) );
  ND2 U2545 ( .A(n4632), .B(n4174), .Z(n2340) );
  MUX21L U2546 ( .A(n4470), .B(n2613), .S(n4949), .Z(n738) );
  ND2 U2547 ( .A(n4212), .B(n4470), .Z(n2613) );
  MUX21L U2548 ( .A(n2412), .B(n2411), .S(n4568), .Z(n734) );
  ND2 U2549 ( .A(n4164), .B(n4861), .Z(n2411) );
  ND2 U2550 ( .A(n4941), .B(n4164), .Z(n2412) );
  MUX21L U2551 ( .A(n2510), .B(n4853), .S(n4594), .Z(n736) );
  ND2 U2552 ( .A(n4227), .B(n4854), .Z(n2510) );
  MUX21L U2553 ( .A(n4736), .B(n4612), .S(n4272), .Z(n745) );
  MUX21L U2554 ( .A(n3183), .B(n3182), .S(n4234), .Z(n748) );
  ND2 U2555 ( .A(n4440), .B(n4784), .Z(n3182) );
  ND2 U2556 ( .A(n4585), .B(n4784), .Z(n3183) );
  MUX21L U2557 ( .A(n4450), .B(n3088), .S(n4252), .Z(n747) );
  ND2 U2558 ( .A(n4906), .B(n4450), .Z(n3088) );
  MUX21L U2559 ( .A(n4785), .B(n4235), .S(n4585), .Z(n718) );
  MUX21L U2560 ( .A(n2820), .B(n2819), .S(n4898), .Z(n712) );
  ND2 U2561 ( .A(n4104), .B(n4493), .Z(n2820) );
  ND2 U2562 ( .A(n4620), .B(n4104), .Z(n2819) );
  MUX21L U2563 ( .A(n4503), .B(n4275), .S(n4915), .Z(n714) );
  MUX21L U2564 ( .A(n4759), .B(n4484), .S(n4242), .Z(n709) );
  MUX21L U2565 ( .A(n4057), .B(n4845), .S(n4610), .Z(n707) );
  MUX21L U2566 ( .A(n4591), .B(n2444), .S(n4942), .Z(n704) );
  ND2 U2567 ( .A(n4591), .B(n4159), .Z(n2444) );
  MUX21L U2568 ( .A(n3030), .B(n3029), .S(n4268), .Z(n686) );
  ND2 U2569 ( .A(n4921), .B(n4454), .Z(n3029) );
  ND2 U2570 ( .A(n4599), .B(n4921), .Z(n3030) );
  MUX21L U2571 ( .A(n2664), .B(n4899), .S(n4214), .Z(n678) );
  ND2 U2572 ( .A(n4899), .B(n4474), .Z(n2664) );
  MUX21L U2573 ( .A(n4769), .B(n3031), .S(n4267), .Z(n655) );
  ND2 U2574 ( .A(n4454), .B(n4769), .Z(n3031) );
  MUX21L U2575 ( .A(n4787), .B(n4438), .S(n4236), .Z(n657) );
  MUX21L U2576 ( .A(n2932), .B(n4146), .S(n4916), .Z(n653) );
  ND2 U2577 ( .A(n4614), .B(n4146), .Z(n2932) );
  MUX21L U2578 ( .A(n4251), .B(n4499), .S(n4895), .Z(n652) );
  MUX21L U2579 ( .A(n2128), .B(n2127), .S(n4280), .Z(n606) );
  ND2 U2580 ( .A(n4425), .B(n4800), .Z(n2127) );
  ND2 U2581 ( .A(n4930), .B(n4579), .Z(n2128) );
  MUX21L U2582 ( .A(n4840), .B(n2665), .S(n4214), .Z(n618) );
  ND2 U2583 ( .A(n4608), .B(n4841), .Z(n2665) );
  MUX21L U2584 ( .A(n4407), .B(n2445), .S(n4942), .Z(n614) );
  ND2 U2585 ( .A(n4224), .B(n4407), .Z(n2445) );
  MUX21L U2586 ( .A(n3033), .B(n3032), .S(n4599), .Z(n623) );
  ND2 U2587 ( .A(n4155), .B(n4770), .Z(n3032) );
  ND2 U2588 ( .A(n4921), .B(n4156), .Z(n3033) );
  MUX21L U2589 ( .A(n4406), .B(n2446), .S(n4224), .Z(n580) );
  ND2 U2590 ( .A(n4407), .B(n4858), .Z(n2446) );
  MUX21L U2591 ( .A(n2634), .B(n4056), .S(n4609), .Z(n551) );
  ND2 U2592 ( .A(n4057), .B(n4844), .Z(n2634) );
  MUX21L U2593 ( .A(n4235), .B(n3189), .S(n4909), .Z(n537) );
  ND2 U2594 ( .A(n4235), .B(n4440), .Z(n3189) );
  ND2 U2595 ( .A(n1915), .B(n1914), .Z(n695) );
  ND2 U2596 ( .A(n4531), .B(n4819), .Z(n1915) );
  ND2 U2597 ( .A(n4257), .B(n4531), .Z(n1914) );
  ND2 U2598 ( .A(n4611), .B(n4734), .Z(n715) );
  ND3 U2599 ( .A(n4495), .B(n4752), .C(n4100), .Z(n505) );
  ND3 U2600 ( .A(n4412), .B(n4861), .C(n4162), .Z(n703) );
  ND3 U2601 ( .A(n4411), .B(n4861), .C(n4161), .Z(n548) );
  ND3 U2602 ( .A(n4494), .B(n4752), .C(n4101), .Z(n531) );
  ND2 U2603 ( .A(n4506), .B(n4740), .Z(n744) );
  MUX41 U2604 ( .D0(n1654), .D1(n1639), .D2(n1645), .D3(n1630), .A(n3871), .B(
        n3884), .Z(N133) );
  ND4 U2605 ( .A(n3825), .B(n3824), .C(n3823), .D(n3822), .Z(n1645) );
  MUX21L U2606 ( .A(n3819), .B(n3818), .S(n3921), .Z(n3824) );
  AO2 U2607 ( .A(n3815), .B(n3958), .C(n3814), .D(n3958), .Z(n3823) );
  MUX21L U2608 ( .A(n3816), .B(n3817), .S(n3921), .Z(n3825) );
  MUX21L U2609 ( .A(n3821), .B(n3820), .S(n3923), .Z(n3822) );
  AN3 U2610 ( .A(n3996), .B(n1642), .C(n3953), .Z(n3821) );
  ND2 U2611 ( .A(n2419), .B(n2418), .Z(n1640) );
  NR3 U2612 ( .A(n3997), .B(n3857), .C(n3958), .Z(n3816) );
  IVP U2613 ( .A(n1644), .Z(n3857) );
  AO7 U2614 ( .A(n4244), .B(n4757), .C(n2764), .Z(n1644) );
  ND2 U2615 ( .A(n4904), .B(n4602), .Z(n2764) );
  MUX41 U2616 ( .D0(n1149), .D1(n1131), .D2(n1140), .D3(n1124), .A(n3872), .B(
        n3883), .Z(N186) );
  NR2 U2617 ( .A(n3998), .B(n37), .Z(n3815) );
  ND2 U2618 ( .A(n4471), .B(n4842), .Z(n2648) );
  MUX41 U2619 ( .D0(n1689), .D1(n1672), .D2(n1680), .D3(n1663), .A(n3871), .B(
        n3884), .Z(N134) );
  NR2 U2620 ( .A(n3998), .B(n38), .Z(n3817) );
  AO6 U2621 ( .A(n4228), .B(n4399), .C(n2520), .Z(n2522) );
  ND4 U2622 ( .A(n3765), .B(n3764), .C(n3763), .D(n3762), .Z(n1131) );
  AO2 U2623 ( .A(n3755), .B(n3923), .C(n3754), .D(n1130), .Z(n3763) );
  MUX21L U2624 ( .A(n3761), .B(n3760), .S(n3921), .Z(n3762) );
  MUX21L U2625 ( .A(n3759), .B(n3758), .S(n3921), .Z(n3764) );
  ND3 U2626 ( .A(n1895), .B(n1894), .C(n1893), .Z(n1660) );
  AO7 U2627 ( .A(n4623), .B(n4200), .C(n4811), .Z(n1662) );
  AO7 U2628 ( .A(n4573), .B(n4113), .C(n4834), .Z(n1656) );
  ND2 U2629 ( .A(n4943), .B(n4405), .Z(n1674) );
  AO7 U2630 ( .A(n4595), .B(n4228), .C(n4946), .Z(n1676) );
  AO7 U2631 ( .A(n4593), .B(n4225), .C(n4943), .Z(n1675) );
  MUX21L U2632 ( .A(n1920), .B(n4134), .S(n4627), .Z(n1627) );
  MUX21L U2633 ( .A(n4822), .B(n4130), .S(n4628), .Z(n1626) );
  AO7 U2634 ( .A(n4937), .B(n4124), .C(n1820), .Z(n1625) );
  MUX41 U2635 ( .D0(n1621), .D1(n1607), .D2(n1612), .D3(n1598), .A(n3871), .B(
        n3884), .Z(N132) );
  MUX41 U2636 ( .D0(n1115), .D1(n1098), .D2(n1106), .D3(n1089), .A(n3872), .B(
        n3883), .Z(N185) );
  NR2 U2637 ( .A(n3957), .B(n3853), .Z(n3758) );
  IVP U2638 ( .A(n1126), .Z(n3853) );
  AO7 U2639 ( .A(n4579), .B(n4189), .C(n4800), .Z(n1126) );
  ND3 U2640 ( .A(n4202), .B(n4813), .C(n4624), .Z(n1087) );
  MUX21L U2641 ( .A(n4135), .B(n4532), .S(n4940), .Z(n1086) );
  MUX21L U2642 ( .A(n4262), .B(n1812), .S(n4937), .Z(n1084) );
  NR2 U2643 ( .A(n4222), .B(n4414), .Z(n1099) );
  NR2 U2644 ( .A(n4944), .B(n4402), .Z(n1101) );
  MUX21L U2645 ( .A(n4491), .B(n4246), .S(n4900), .Z(n1107) );
  ND2 U2646 ( .A(n4913), .B(n2875), .Z(n1108) );
  MUX21L U2647 ( .A(n4142), .B(n4914), .S(n4615), .Z(n1109) );
  ND2 U2648 ( .A(n4606), .B(n4217), .Z(n1611) );
  AO7 U2649 ( .A(n4916), .B(n4147), .C(n4505), .Z(n1615) );
  AO7 U2650 ( .A(n4910), .B(n4587), .C(n4080), .Z(n1619) );
  ND2 U2651 ( .A(n2837), .B(n2836), .Z(n1614) );
  AN3 U2652 ( .A(n3996), .B(n3952), .C(n1125), .Z(n3760) );
  MUX21L U2653 ( .A(n4621), .B(n4926), .S(n4297), .Z(n1125) );
  IVP U2654 ( .A(n4721), .Z(n4957) );
  IVP U2655 ( .A(n4721), .Z(n4955) );
  IVP U2656 ( .A(n4721), .Z(n4956) );
  NR3 U2657 ( .A(n39), .B(n3999), .C(n3954), .Z(n3549) );
  ND2 U2658 ( .A(n4901), .B(n4245), .Z(n2785) );
  NR3 U2659 ( .A(n41), .B(n3999), .C(n3954), .Z(n3548) );
  ND2 U2660 ( .A(n4229), .B(n4462), .Z(n2560) );
  NR3 U2661 ( .A(n42), .B(n3998), .C(n3927), .Z(n3545) );
  ND2 U2662 ( .A(n4215), .B(n4477), .Z(n2677) );
  MUX41 U2663 ( .D0(n1081), .D1(n1069), .D2(n1073), .D3(n1060), .A(n3872), .B(
        n3883), .Z(N184) );
  AO7 U2664 ( .A(n4954), .B(n4180), .C(n4557), .Z(n1066) );
  ND2 U2665 ( .A(n2062), .B(n4640), .Z(n1062) );
  MUX21L U2666 ( .A(n2035), .B(n4195), .S(n4926), .Z(n1061) );
  ND2 U2667 ( .A(n4124), .B(n4524), .Z(n1055) );
  ND2 U2668 ( .A(n4256), .B(n4819), .Z(n1057) );
  AO7 U2669 ( .A(n4624), .B(n4811), .C(n4295), .Z(n1059) );
  AN3 U2670 ( .A(n1071), .B(n3914), .C(n3994), .Z(n3547) );
  MUX21L U2671 ( .A(n2489), .B(n4944), .S(n4593), .Z(n1071) );
  ND2 U2672 ( .A(n4944), .B(n4068), .Z(n2489) );
  AN3 U2673 ( .A(n1070), .B(n3914), .C(n3994), .Z(n3546) );
  MUX21L U2674 ( .A(n4413), .B(n2405), .S(n4941), .Z(n1070) );
  ND2 U2675 ( .A(n4222), .B(n4414), .Z(n2405) );
  ND3 U2676 ( .A(n3552), .B(n3551), .C(n3550), .Z(n1073) );
  MUX21L U2677 ( .A(n3544), .B(n3545), .S(n3955), .Z(n3552) );
  MUX21L U2678 ( .A(n3547), .B(n3546), .S(n3954), .Z(n3550) );
  MUX21L U2679 ( .A(n3549), .B(n3548), .S(n3927), .Z(n3551) );
  MUX41 U2680 ( .D0(n1589), .D1(n1571), .D2(n1580), .D3(n1562), .A(n3873), .B(
        n3884), .Z(N131) );
  IVP U2681 ( .A(n4721), .Z(n4958) );
  NR2 U2682 ( .A(n4002), .B(n3955), .Z(n3754) );
  NR2 U2683 ( .A(n4002), .B(n3957), .Z(n3755) );
  AO4 U2684 ( .A(n4618), .B(n4248), .C(n4896), .D(n4619), .Z(n1582) );
  ND2 U2685 ( .A(n2948), .B(n2947), .Z(n1584) );
  MUX21L U2686 ( .A(n4910), .B(n4439), .S(n4235), .Z(n1587) );
  ND3 U2687 ( .A(n4575), .B(n4121), .C(n4936), .Z(n1556) );
  MUX21L U2688 ( .A(n4813), .B(n4294), .S(n4624), .Z(n1561) );
  MUX21L U2689 ( .A(n4292), .B(n1931), .S(n4626), .Z(n1560) );
  AN3 U2690 ( .A(n3952), .B(n1127), .C(n3996), .Z(n3761) );
  ND2 U2691 ( .A(n4185), .B(n4877), .Z(n1127) );
  IVP U2692 ( .A(n4721), .Z(n4954) );
  MUX41 U2693 ( .D0(n1051), .D1(n1035), .D2(n1044), .D3(n1026), .A(n3872), .B(
        n3882), .Z(N183) );
  NR2 U2694 ( .A(n4580), .B(n4138), .Z(n1030) );
  AO7 U2695 ( .A(n4284), .B(n4878), .C(n4551), .Z(n1031) );
  ND3 U2696 ( .A(n4569), .B(n4172), .C(n4957), .Z(n1033) );
  AN3 U2697 ( .A(n1045), .B(n3995), .C(n3914), .Z(n3649) );
  ND2 U2698 ( .A(n2807), .B(n2806), .Z(n1045) );
  ND2 U2699 ( .A(n2803), .B(n4491), .Z(n2806) );
  MUX21L U2700 ( .A(n2804), .B(n2805), .S(n4246), .Z(n2807) );
  EO U2701 ( .A(n4890), .B(n4590), .Z(n435) );
  MUX41 U2702 ( .D0(n1553), .D1(n1535), .D2(n1544), .D3(n1528), .A(n3873), .B(
        n3884), .Z(N130) );
  ND4 U2703 ( .A(n3777), .B(n3776), .C(n3775), .D(n3774), .Z(n1535) );
  MUX21L U2704 ( .A(n3768), .B(n3769), .S(n3921), .Z(n3777) );
  AO2 U2705 ( .A(n3767), .B(n4001), .C(n3766), .D(n1534), .Z(n3775) );
  MUX21L U2706 ( .A(n3770), .B(n3771), .S(n3957), .Z(n3776) );
  NR2 U2707 ( .A(n4628), .B(n4133), .Z(n1023) );
  NR2 U2708 ( .A(n4576), .B(n4262), .Z(n1021) );
  AO7 U2709 ( .A(n4924), .B(n4538), .C(n4295), .Z(n1025) );
  MUX21L U2710 ( .A(n3773), .B(n3772), .S(n3923), .Z(n3774) );
  AN3 U2711 ( .A(n1529), .B(n3952), .C(n3996), .Z(n3772) );
  MUX21L U2712 ( .A(n4195), .B(n4807), .S(n4641), .Z(n1529) );
  MUX41 U2713 ( .D0(n1017), .D1(n1001), .D2(n1009), .D3(n992), .A(n3872), .B(
        n3882), .Z(N182) );
  ND2 U2714 ( .A(n4230), .B(n4460), .Z(n1539) );
  ND2 U2715 ( .A(n2589), .B(n2588), .Z(n1540) );
  MUX21L U2716 ( .A(n4758), .B(n2745), .S(n4604), .Z(n1543) );
  AN3 U2717 ( .A(n987), .B(n3916), .C(n3951), .Z(n3329) );
  ND2 U2718 ( .A(n1743), .B(n1742), .Z(n987) );
  ND2 U2719 ( .A(n4934), .B(n4289), .Z(n1742) );
  EN U2720 ( .A(n4891), .B(n4573), .Z(n1743) );
  NR3 U2721 ( .A(n3957), .B(n4000), .C(n43), .Z(n3769) );
  ND2 U2722 ( .A(n4951), .B(n4140), .Z(n2181) );
  ND2 U2723 ( .A(n4281), .B(n4424), .Z(n1531) );
  NR2 U2724 ( .A(n3957), .B(n3923), .Z(n3766) );
  NR2 U2725 ( .A(n3957), .B(n3921), .Z(n3767) );
  ND2 U2726 ( .A(n4613), .B(n4148), .Z(n1012) );
  AO7 U2727 ( .A(n4899), .B(n4621), .C(n4246), .Z(n1010) );
  ND3 U2728 ( .A(n4465), .B(n4796), .C(n4242), .Z(n1016) );
  NR3 U2729 ( .A(n4300), .B(n4928), .C(n4639), .Z(n994) );
  ND3 U2730 ( .A(n4255), .B(n4883), .C(n4566), .Z(n996) );
  MUX21L U2731 ( .A(n4809), .B(n2022), .S(n4621), .Z(n993) );
  NR3 U2732 ( .A(n3850), .B(n3960), .C(n3931), .Z(n3328) );
  IVP U2733 ( .A(n991), .Z(n3850) );
  AO7 U2734 ( .A(n4923), .B(n4624), .C(n4202), .Z(n991) );
  MUX41 U2735 ( .D0(n1519), .D1(n1501), .D2(n1510), .D3(n1493), .A(n3873), .B(
        n3884), .Z(N129) );
  MUX41 U2736 ( .D0(n986), .D1(n971), .D2(n980), .D3(n963), .A(n3872), .B(
        n3882), .Z(N181) );
  ND4 U2737 ( .A(n3710), .B(n3709), .C(n3708), .D(n3707), .Z(n963) );
  MUX21L U2738 ( .A(n3705), .B(n3706), .S(n3922), .Z(n3707) );
  MUX21L U2739 ( .A(n3701), .B(n3702), .S(n3923), .Z(n3709) );
  MUX21L U2740 ( .A(n3699), .B(n3700), .S(n4004), .Z(n3710) );
  AO7 U2741 ( .A(n4936), .B(n4576), .C(n4121), .Z(n1487) );
  MUX21L U2742 ( .A(n4256), .B(n1919), .S(n4627), .Z(n1490) );
  MUX21L U2743 ( .A(n4576), .B(n4936), .S(n4263), .Z(n1488) );
  MUX21L U2744 ( .A(n4765), .B(n4477), .S(n4216), .Z(n1507) );
  MUX21L U2745 ( .A(n4467), .B(n2590), .S(n4212), .Z(n1506) );
  MUX21L U2746 ( .A(n2524), .B(n2523), .S(n4595), .Z(n1505) );
  NR3 U2747 ( .A(n45), .B(n3957), .C(n3922), .Z(n3699) );
  NR2 U2748 ( .A(n1990), .B(n1989), .Z(n1992) );
  ND2 U2749 ( .A(n3081), .B(n3080), .Z(n984) );
  MUX21L U2750 ( .A(n4918), .B(n4612), .S(n4272), .Z(n983) );
  MUX21L U2751 ( .A(n2927), .B(n4740), .S(n4614), .Z(n982) );
  AN3 U2752 ( .A(n964), .B(n3994), .C(n3915), .Z(n3433) );
  MUX21L U2753 ( .A(n2023), .B(n4621), .S(n4297), .Z(n964) );
  ND2 U2754 ( .A(n4926), .B(n4621), .Z(n2023) );
  ND2 U2755 ( .A(n1746), .B(n1745), .Z(n958) );
  ND2 U2756 ( .A(n4573), .B(n4289), .Z(n1745) );
  MUX21L U2757 ( .A(n1744), .B(n4289), .S(n4934), .Z(n1746) );
  ND2 U2758 ( .A(n1791), .B(n1790), .Z(n959) );
  ND2 U2759 ( .A(n4936), .B(n4263), .Z(n1790) );
  EO U2760 ( .A(n4563), .B(n4263), .Z(n1791) );
  MUX41 U2761 ( .D0(n1485), .D1(n1469), .D2(n1477), .D3(n1460), .A(n3872), .B(
        n3883), .Z(N128) );
  NR2 U2762 ( .A(n4221), .B(n4865), .Z(n1470) );
  AO7 U2763 ( .A(n4943), .B(n4225), .C(n4405), .Z(n1471) );
  MUX41 U2764 ( .D0(n957), .D1(n940), .D2(n948), .D3(n936), .A(n3872), .B(
        n3882), .Z(N180) );
  ND4 U2765 ( .A(n3753), .B(n3752), .C(n3751), .D(n3750), .Z(n940) );
  AO2 U2766 ( .A(n3743), .B(n3957), .C(n3742), .D(n3957), .Z(n3751) );
  MUX21L U2767 ( .A(n3744), .B(n3745), .S(n3921), .Z(n3753) );
  MUX21L U2768 ( .A(n3747), .B(n3746), .S(n3921), .Z(n3752) );
  NR2 U2769 ( .A(n4626), .B(n4291), .Z(n1453) );
  AN3 U2770 ( .A(n4563), .B(n4209), .C(n4885), .Z(n1458) );
  ND2 U2771 ( .A(n1735), .B(n1734), .Z(n1454) );
  NR2 U2772 ( .A(n4898), .B(n4052), .Z(n945) );
  NR2 U2773 ( .A(n4902), .B(n4486), .Z(n947) );
  NR2 U2774 ( .A(n4568), .B(n4222), .Z(n941) );
  MUX21L U2775 ( .A(n3749), .B(n3748), .S(n3921), .Z(n3750) );
  AN3 U2776 ( .A(n3996), .B(n938), .C(n3952), .Z(n3749) );
  ND2 U2777 ( .A(n4636), .B(n4297), .Z(n937) );
  MUX41 U2778 ( .D0(n1452), .D1(n1434), .D2(n1443), .D3(n1426), .A(n3873), .B(
        n3883), .Z(N127) );
  NR2 U2779 ( .A(n4003), .B(n47), .Z(n3745) );
  EN U2780 ( .A(n4888), .B(n4639), .Z(n2183) );
  ND4 U2781 ( .A(n3698), .B(n3697), .C(n3696), .D(n3695), .Z(n1426) );
  MUX21L U2782 ( .A(n3687), .B(n3688), .S(n3956), .Z(n3698) );
  MUX21L U2783 ( .A(n3690), .B(n3689), .S(n3923), .Z(n3697) );
  MUX21L U2784 ( .A(n3693), .B(n3694), .S(n3925), .Z(n3695) );
  ND2 U2785 ( .A(n1910), .B(n1909), .Z(n933) );
  MUX21L U2786 ( .A(n1980), .B(n4623), .S(n4295), .Z(n935) );
  MUX21L U2787 ( .A(n4836), .B(n1718), .S(n4290), .Z(n929) );
  NR3 U2788 ( .A(n4003), .B(n2376), .C(n3957), .Z(n3744) );
  ND2 U2789 ( .A(n4570), .B(n4220), .Z(n2376) );
  ND2 U2790 ( .A(n1861), .B(n1860), .Z(n1423) );
  ND2 U2791 ( .A(n4259), .B(n4527), .Z(n1860) );
  EO U2792 ( .A(n4893), .B(n4259), .Z(n1861) );
  ND2 U2793 ( .A(n1750), .B(n1749), .Z(n1422) );
  ND2 U2794 ( .A(n4265), .B(n4517), .Z(n1749) );
  MUX21L U2795 ( .A(n4934), .B(n1748), .S(n4573), .Z(n1750) );
  NR2 U2796 ( .A(n4003), .B(n4958), .Z(n3743) );
  MUX41 U2797 ( .D0(n928), .D1(n913), .D2(n920), .D3(n908), .A(n3872), .B(
        n3882), .Z(N179) );
  NR3 U2798 ( .A(n3956), .B(n4003), .C(n46), .Z(n3689) );
  NR2 U2799 ( .A(n1823), .B(n1822), .Z(n1825) );
  ND4 U2800 ( .A(n3813), .B(n3812), .C(n3811), .D(n3810), .Z(n920) );
  MUX21L U2801 ( .A(n3802), .B(n3803), .S(n3999), .Z(n3813) );
  MUX21L U2802 ( .A(n3804), .B(n3805), .S(n3922), .Z(n3812) );
  MUX21L U2803 ( .A(n3808), .B(n3809), .S(n3921), .Z(n3810) );
  MUX21L U2804 ( .A(n2885), .B(n2884), .S(n4616), .Z(n1446) );
  MUX21L U2805 ( .A(n4786), .B(n4439), .S(n4235), .Z(n1450) );
  MUX21L U2806 ( .A(n4751), .B(n4618), .S(n4248), .Z(n1445) );
  NR2 U2807 ( .A(n3956), .B(n3852), .Z(n3690) );
  IVP U2808 ( .A(n1425), .Z(n3852) );
  AO7 U2809 ( .A(n4925), .B(n4540), .C(n2014), .Z(n1425) );
  ND2 U2810 ( .A(n4622), .B(n4296), .Z(n2014) );
  EN U2811 ( .A(n4893), .B(n4227), .Z(n915) );
  MUX21L U2812 ( .A(n3785), .B(n3784), .S(n3922), .Z(n3786) );
  AN3 U2813 ( .A(n3953), .B(n912), .C(n3997), .Z(n3785) );
  AN3 U2814 ( .A(n3997), .B(n3953), .C(n909), .Z(n3784) );
  ND2 U2815 ( .A(n2235), .B(n2234), .Z(n912) );
  MUX41 U2816 ( .D0(n1420), .D1(n1403), .D2(n1411), .D3(n1395), .A(n3871), .B(
        n3883), .Z(N126) );
  EN U2817 ( .A(n4890), .B(n4636), .Z(n436) );
  NR2 U2818 ( .A(n3957), .B(n48), .Z(n3783) );
  ND2 U2819 ( .A(n4287), .B(n4559), .Z(n2317) );
  MUX21L U2820 ( .A(n4257), .B(n1911), .S(n4939), .Z(n905) );
  MUX21L U2821 ( .A(n4835), .B(n1719), .S(n4572), .Z(n901) );
  ND2 U2822 ( .A(n1983), .B(n1982), .Z(n907) );
  MUX21L U2823 ( .A(n4591), .B(n2438), .S(n4942), .Z(n914) );
  ND2 U2824 ( .A(n4591), .B(n4159), .Z(n2438) );
  NR3 U2825 ( .A(n49), .B(n3958), .C(n3922), .Z(n3802) );
  ND2 U2826 ( .A(n4903), .B(n4486), .Z(n2755) );
  EN U2827 ( .A(n4562), .B(n4294), .Z(n437) );
  NR2 U2828 ( .A(n4000), .B(n3957), .Z(n3778) );
  NR2 U2829 ( .A(n4000), .B(n3957), .Z(n3779) );
  MUX41 U2830 ( .D0(n900), .D1(n886), .D2(n892), .D3(n879), .A(n3872), .B(
        n3882), .Z(N178) );
  ND4 U2831 ( .A(n3837), .B(n3836), .C(n3835), .D(n3834), .Z(n892) );
  MUX21L U2832 ( .A(n3826), .B(n3827), .S(n3998), .Z(n3837) );
  MUX21L U2833 ( .A(n3828), .B(n3829), .S(n3923), .Z(n3836) );
  MUX21L U2834 ( .A(n3833), .B(n3832), .S(n3958), .Z(n3834) );
  ND2 U2835 ( .A(n4897), .B(n4483), .Z(n1409) );
  MUX21L U2836 ( .A(n4941), .B(n4222), .S(n4569), .Z(n1404) );
  AN3 U2837 ( .A(n1390), .B(n3952), .C(n3915), .Z(n3395) );
  ND3 U2838 ( .A(n1710), .B(n1709), .C(n1708), .Z(n1390) );
  ND2 U2839 ( .A(n4109), .B(n4520), .Z(n1709) );
  ND2 U2840 ( .A(n4933), .B(n4521), .Z(n1710) );
  NR3 U2841 ( .A(n3922), .B(n3958), .C(n3858), .Z(n3826) );
  IVP U2842 ( .A(n891), .Z(n3858) );
  AO7 U2843 ( .A(n4602), .B(n4040), .C(n2773), .Z(n891) );
  ND2 U2844 ( .A(n4903), .B(n4245), .Z(n2773) );
  NR3 U2845 ( .A(n50), .B(n3997), .C(n3958), .Z(n3829) );
  ND2 U2846 ( .A(n4464), .B(n4851), .Z(n2546) );
  ND2 U2847 ( .A(n2319), .B(n2318), .Z(n885) );
  AO7 U2848 ( .A(n4298), .B(n4544), .C(n2042), .Z(n880) );
  ND2 U2849 ( .A(n2140), .B(n2139), .Z(n881) );
  MUX21L U2850 ( .A(n4530), .B(n1912), .S(n4257), .Z(n876) );
  ND2 U2851 ( .A(n1809), .B(n1808), .Z(n874) );
  MUX21L U2852 ( .A(n4623), .B(n1984), .S(n4924), .Z(n878) );
  AN3 U2853 ( .A(n3916), .B(n888), .C(n3996), .Z(n3833) );
  ND2 U2854 ( .A(n2494), .B(n2493), .Z(n888) );
  ND2 U2855 ( .A(n4226), .B(n4401), .Z(n2493) );
  MUX21L U2856 ( .A(n4944), .B(n2492), .S(n4593), .Z(n2494) );
  MUX41 U2857 ( .D0(n1389), .D1(n1373), .D2(n1381), .D3(n1365), .A(n3872), .B(
        n3883), .Z(N125) );
  ND2 U2858 ( .A(n4617), .B(n4747), .Z(n1382) );
  MUX21L U2859 ( .A(n3070), .B(n4601), .S(n4251), .Z(n1386) );
  MUX21L U2860 ( .A(n4273), .B(n2950), .S(n4613), .Z(n1384) );
  AN3 U2861 ( .A(n4733), .B(n3952), .C(n3915), .Z(n3396) );
  ND2 U2862 ( .A(n4606), .B(n4050), .Z(n889) );
  MUX21L U2863 ( .A(n4820), .B(n1903), .S(n4258), .Z(n1363) );
  ND2 U2864 ( .A(n1789), .B(n1788), .Z(n1360) );
  EO U2865 ( .A(n4890), .B(n4571), .Z(n1359) );
  MUX41 U2866 ( .D0(n871), .D1(n857), .D2(n864), .D3(n849), .A(n3873), .B(
        n3882), .Z(N177) );
  NR3 U2867 ( .A(n53), .B(n3960), .C(n3931), .Z(n3338) );
  ND2 U2868 ( .A(n4923), .B(n4293), .Z(n1965) );
  MUX41 U2869 ( .D0(n1358), .D1(n1344), .D2(n1352), .D3(n1337), .A(LogIn2[47]), 
        .B(n3883), .Z(N124) );
  NR2 U2870 ( .A(n4581), .B(n4092), .Z(n868) );
  MUX21L U2871 ( .A(n4084), .B(n4584), .S(n4909), .Z(n869) );
  ND2 U2872 ( .A(n2834), .B(n4101), .Z(n865) );
  ND3 U2873 ( .A(n2156), .B(n2155), .C(n2154), .Z(n853) );
  EO U2874 ( .A(n4561), .B(n4300), .Z(n851) );
  MUX21L U2875 ( .A(n4554), .B(n2268), .S(n4285), .Z(n855) );
  NR3 U2876 ( .A(n51), .B(n3955), .C(n3926), .Z(n3576) );
  ND2 U2877 ( .A(n4443), .B(n4781), .Z(n3149) );
  ND2 U2878 ( .A(n4162), .B(n4412), .Z(n1345) );
  MUX21L U2879 ( .A(n4482), .B(n4761), .S(n4219), .Z(n1351) );
  ND2 U2880 ( .A(n4610), .B(n2623), .Z(n1349) );
  AN3 U2881 ( .A(n1353), .B(n3914), .C(n3951), .Z(n3577) );
  NR2 U2882 ( .A(n4618), .B(n4248), .Z(n1353) );
  MUX41 U2883 ( .D0(n844), .D1(n829), .D2(n836), .D3(n823), .A(n3873), .B(
        n3882), .Z(N176) );
  OR3 U2884 ( .A(n4290), .B(n4933), .C(n4572), .Z(n438) );
  NR2 U2885 ( .A(n4014), .B(n3851), .Z(n3348) );
  IVP U2886 ( .A(n822), .Z(n3851) );
  AO4 U2887 ( .A(n4623), .B(n4295), .C(n4924), .D(n4295), .Z(n822) );
  MUX41 U2888 ( .D0(n1329), .D1(n1311), .D2(n1320), .D3(n1303), .A(n3871), .B(
        n3883), .Z(N123) );
  MUX21L U2889 ( .A(n4408), .B(n2440), .S(n4223), .Z(n830) );
  EO U2890 ( .A(n4891), .B(n4610), .Z(n832) );
  ND3 U2891 ( .A(n2497), .B(n2496), .C(n2495), .Z(n831) );
  NR2 U2892 ( .A(n4920), .B(n4598), .Z(n840) );
  NR3 U2893 ( .A(n4276), .B(n4915), .C(n4615), .Z(n838) );
  AO7 U2894 ( .A(n4238), .B(n4435), .C(n4911), .Z(n843) );
  ND3 U2895 ( .A(n3355), .B(n3354), .C(n3353), .Z(n823) );
  MUX21L U2896 ( .A(n3351), .B(n3352), .S(n4014), .Z(n3354) );
  MUX21L U2897 ( .A(n3348), .B(n3347), .S(n3930), .Z(n3353) );
  MUX21L U2898 ( .A(n3349), .B(n3350), .S(n3960), .Z(n3355) );
  ND2 U2899 ( .A(n1967), .B(n1966), .Z(n821) );
  ND2 U2900 ( .A(n4923), .B(n4294), .Z(n1967) );
  ND2 U2901 ( .A(n4625), .B(n4294), .Z(n1966) );
  NR3 U2902 ( .A(n55), .B(n3960), .C(n3931), .Z(n3300) );
  ND2 U2903 ( .A(n4626), .B(n4204), .Z(n1938) );
  ND2 U2904 ( .A(n2579), .B(n4060), .Z(n1315) );
  ND2 U2905 ( .A(n2654), .B(n2653), .Z(n1317) );
  ND2 U2906 ( .A(n2483), .B(n2482), .Z(n1314) );
  AN3 U2907 ( .A(n845), .B(n3915), .C(n3951), .Z(n3339) );
  ND3 U2908 ( .A(n4517), .B(n4833), .C(n4117), .Z(n845) );
  NR3 U2909 ( .A(n56), .B(n4013), .C(n3960), .Z(n3304) );
  ND2 U2910 ( .A(n4537), .B(n4812), .Z(n1976) );
  MUX41 U2911 ( .D0(n820), .D1(n806), .D2(n812), .D3(n801), .A(n3873), .B(
        n3882), .Z(N175) );
  ND2 U2912 ( .A(n3359), .B(n3358), .Z(n801) );
  NR2 U2913 ( .A(n3960), .B(n4072), .Z(n3347) );
  OR3 U2914 ( .A(n4288), .B(n4955), .C(n4633), .Z(n439) );
  ND2 U2915 ( .A(n4088), .B(n4779), .Z(n817) );
  ND2 U2916 ( .A(n4922), .B(n4096), .Z(n816) );
  ND2 U2917 ( .A(n4909), .B(n4584), .Z(n818) );
  MUX41 U2918 ( .D0(n1297), .D1(n1279), .D2(n1288), .D3(n1271), .A(n3871), .B(
        n3883), .Z(N122) );
  ND4 U2919 ( .A(n3318), .B(n3317), .C(n3316), .D(n3315), .Z(n1271) );
  NR3 U2920 ( .A(n3856), .B(n3999), .C(n3954), .Z(n3517) );
  IVP U2921 ( .A(n811), .Z(n3856) );
  AO7 U2922 ( .A(n4903), .B(n4042), .C(n4603), .Z(n811) );
  ND2 U2923 ( .A(n2402), .B(n2401), .Z(n1280) );
  MUX21L U2924 ( .A(n2529), .B(n4946), .S(n4228), .Z(n1283) );
  ND2 U2925 ( .A(n2485), .B(n2484), .Z(n1282) );
  AO7 U2926 ( .A(n4237), .B(n4790), .C(n4587), .Z(n1296) );
  MUX21L U2927 ( .A(n4090), .B(n4445), .S(n4907), .Z(n1294) );
  MUX21L U2928 ( .A(n4751), .B(n4249), .S(n4618), .Z(n1290) );
  NR2 U2929 ( .A(n4641), .B(n4297), .Z(n802) );
  MUX41 U2930 ( .D0(n799), .D1(n786), .D2(n790), .D3(n784), .A(n3873), .B(
        n3882), .Z(N174) );
  ND2 U2931 ( .A(n3361), .B(n3360), .Z(n784) );
  AN3 U2932 ( .A(n807), .B(n3914), .C(n3952), .Z(n3514) );
  ND2 U2933 ( .A(n4071), .B(n4404), .Z(n807) );
  MUX41 U2934 ( .D0(n1266), .D1(n1249), .D2(n1258), .D3(n1243), .A(n3872), .B(
        n3883), .Z(N121) );
  ND2 U2935 ( .A(n3324), .B(n3323), .Z(n1243) );
  ND4 U2936 ( .A(n3741), .B(n3740), .C(n3739), .D(n3738), .Z(n1249) );
  MUX21L U2937 ( .A(n3730), .B(n3731), .S(n4000), .Z(n3741) );
  MUX21L U2938 ( .A(n3734), .B(n3735), .S(n4004), .Z(n3739) );
  MUX21L U2939 ( .A(n3732), .B(n3733), .S(n3922), .Z(n3740) );
  AO7 U2940 ( .A(n4907), .B(n4445), .C(n4089), .Z(n796) );
  ND2 U2941 ( .A(n2818), .B(n2817), .Z(n791) );
  MUX21L U2942 ( .A(n3235), .B(n3234), .S(n4588), .Z(n798) );
  AN3 U2943 ( .A(n788), .B(n3994), .C(n3951), .Z(n3526) );
  AO7 U2944 ( .A(n4949), .B(n4610), .C(n4212), .Z(n788) );
  ND2 U2945 ( .A(n3476), .B(n3475), .Z(n786) );
  EO U2946 ( .A(n3953), .B(n3928), .Z(n3475) );
  MUX21L U2947 ( .A(n3474), .B(n3473), .S(n3928), .Z(n3476) );
  NR2 U2948 ( .A(n4016), .B(n413), .Z(n3474) );
  ND2 U2949 ( .A(n2404), .B(n2403), .Z(n1250) );
  MUX21L U2950 ( .A(n4410), .B(n2432), .S(n4223), .Z(n1251) );
  ND2 U2951 ( .A(n2517), .B(n2516), .Z(n1252) );
  NR2 U2952 ( .A(n4638), .B(n4282), .Z(n1247) );
  IVP U2953 ( .A(n782), .Z(n3861) );
  ND2 U2954 ( .A(n2882), .B(n4141), .Z(n775) );
  MUX21L U2955 ( .A(n4788), .B(n4080), .S(n4586), .Z(n780) );
  MUX21L U2956 ( .A(n3412), .B(n3411), .S(n3871), .Z(n3414) );
  NR2 U2957 ( .A(n3885), .B(n59), .Z(n3411) );
  NR2 U2958 ( .A(n3885), .B(n3861), .Z(n3412) );
  ND2 U2959 ( .A(n2087), .B(n2086), .Z(n1244) );
  ND2 U2960 ( .A(n4929), .B(n4278), .Z(n2087) );
  ND2 U2961 ( .A(n4577), .B(n4278), .Z(n2086) );
  NR3 U2962 ( .A(n4236), .B(n3957), .C(n3924), .Z(n3730) );
  NR3 U2963 ( .A(n4300), .B(n3998), .C(n3927), .Z(n3522) );
  MUX21L U2964 ( .A(n3321), .B(n3322), .S(n3931), .Z(n3323) );
  NR3 U2965 ( .A(n3960), .B(n4014), .C(n3849), .Z(n3322) );
  ND3 U2966 ( .A(n4533), .B(n4817), .C(n4205), .Z(n1242) );
  MUX21L U2967 ( .A(n3533), .B(n3532), .S(n3954), .Z(n3537) );
  NR2 U2968 ( .A(n3998), .B(n2324), .Z(n3533) );
  NR2 U2969 ( .A(n3927), .B(n60), .Z(n3532) );
  MUX41 U2970 ( .D0(n1240), .D1(n1223), .D2(n1232), .D3(n1221), .A(n3872), .B(
        n3883), .Z(N120) );
  AO7 U2971 ( .A(n417), .B(n3326), .C(n3325), .Z(n1221) );
  NR2 U2972 ( .A(n4911), .B(n4587), .Z(n1239) );
  ND2 U2973 ( .A(n4618), .B(n4249), .Z(n1234) );
  MUX21L U2974 ( .A(n4767), .B(n3003), .S(n4269), .Z(n1236) );
  ND3 U2975 ( .A(n3447), .B(n3446), .C(n3445), .Z(n1223) );
  MUX21L U2976 ( .A(n3440), .B(n3959), .S(n4016), .Z(n3446) );
  MUX21L U2977 ( .A(n3442), .B(n3441), .S(n3958), .Z(n3447) );
  MUX21L U2978 ( .A(n3443), .B(n3444), .S(n3958), .Z(n3445) );
  ND2 U2979 ( .A(n2089), .B(n2088), .Z(n1222) );
  ND2 U2980 ( .A(n4929), .B(n4278), .Z(n2089) );
  ND2 U2981 ( .A(n4577), .B(n4278), .Z(n2088) );
  OR3 U2982 ( .A(n4287), .B(n4955), .C(n4634), .Z(n440) );
  NR2 U2983 ( .A(n4016), .B(n413), .Z(n3442) );
  NR2 U2984 ( .A(n3954), .B(n3927), .Z(n3534) );
  AN3 U2985 ( .A(n766), .B(n3913), .C(n3951), .Z(n3621) );
  AO4 U2986 ( .A(n4618), .B(n4249), .C(n4895), .D(n4249), .Z(n766) );
  ND2 U2987 ( .A(n3725), .B(n3724), .Z(N119) );
  AO2 U2988 ( .A(n3885), .B(n1211), .C(n3885), .D(n3871), .Z(n3725) );
  MUX21L U2989 ( .A(n3723), .B(n1205), .S(n3871), .Z(n3724) );
  NR3 U2990 ( .A(n3177), .B(n3955), .C(n3925), .Z(n3620) );
  ND3 U2991 ( .A(n4234), .B(n4784), .C(n4585), .Z(n3177) );
  MUX21L U2992 ( .A(n3632), .B(n3631), .S(n3955), .Z(n3637) );
  NR2 U2993 ( .A(n4002), .B(n62), .Z(n3632) );
  NR3 U2994 ( .A(n4002), .B(n414), .C(n3925), .Z(n3631) );
  NR2 U2995 ( .A(n3885), .B(n3863), .Z(n3723) );
  IVP U2996 ( .A(n1220), .Z(n3863) );
  MUX21L U2997 ( .A(n4614), .B(n4145), .S(n4916), .Z(n1214) );
  NR2 U2998 ( .A(n3958), .B(n3929), .Z(n3440) );
  NR3 U2999 ( .A(n3856), .B(n3998), .C(n3953), .Z(n3495) );
  NR2 U3000 ( .A(n3929), .B(n4106), .Z(n3441) );
  NR2 U3001 ( .A(n3956), .B(n3848), .Z(n3630) );
  IVP U3002 ( .A(n761), .Z(n3848) );
  AO4 U3003 ( .A(n4615), .B(n4275), .C(n4915), .D(n4275), .Z(n761) );
  NR3 U3004 ( .A(n61), .B(n3953), .C(n3928), .Z(n3491) );
  ND2 U3005 ( .A(n4480), .B(n4763), .Z(n2707) );
  ND2 U3006 ( .A(n2091), .B(n2090), .Z(n1204) );
  ND2 U3007 ( .A(n4929), .B(n4278), .Z(n2091) );
  ND2 U3008 ( .A(n4577), .B(n4278), .Z(n2090) );
  NR2 U3009 ( .A(n3884), .B(n3862), .Z(n3404) );
  IVP U3010 ( .A(n1203), .Z(n3862) );
  AO7 U3011 ( .A(n4895), .B(n4099), .C(n4618), .Z(n1196) );
  AN3 U3012 ( .A(n3951), .B(n762), .C(n3995), .Z(n3633) );
  NR2 U3013 ( .A(n4599), .B(n4268), .Z(n762) );
  OR3 U3014 ( .A(n4214), .B(n4897), .C(n4608), .Z(n441) );
  NR2 U3015 ( .A(n4016), .B(n4242), .Z(n3449) );
  OR3 U3016 ( .A(n4226), .B(n4944), .C(n4593), .Z(n442) );
  AN3 U3017 ( .A(n3952), .B(n1192), .C(n3994), .Z(n3504) );
  ND2 U3018 ( .A(n2642), .B(n4055), .Z(n1192) );
  ND2 U3019 ( .A(n4896), .B(n4609), .Z(n2642) );
  ND3 U3020 ( .A(n3508), .B(n3507), .C(n3506), .Z(n1194) );
  MUX21L U3021 ( .A(n3500), .B(n3501), .S(n3928), .Z(n3507) );
  MUX21L U3022 ( .A(n3504), .B(n3505), .S(n3928), .Z(n3506) );
  MUX21L U3023 ( .A(n3503), .B(n3502), .S(n3953), .Z(n3508) );
  NR2 U3024 ( .A(n3997), .B(n4230), .Z(n3503) );
  NR2 U3025 ( .A(n3884), .B(n3864), .Z(n3403) );
  IVP U3026 ( .A(n1191), .Z(n3864) );
  AO3 U3027 ( .A(n4015), .B(n3849), .C(n3930), .D(n3959), .Z(n1191) );
  NR2 U3028 ( .A(n4002), .B(n3956), .Z(n3634) );
  NR2 U3029 ( .A(n4003), .B(n3849), .Z(n3675) );
  MUX21L U3030 ( .A(n4585), .B(n3181), .S(n4909), .Z(n758) );
  ND2 U3031 ( .A(n4585), .B(n4083), .Z(n3181) );
  NR2 U3032 ( .A(n3998), .B(n3953), .Z(n3505) );
  NR2 U3033 ( .A(n3924), .B(n65), .Z(n3639) );
  ND2 U3034 ( .A(n4239), .B(n4434), .Z(n3243) );
  AO7 U3035 ( .A(n4253), .B(n4447), .C(n4776), .Z(n1187) );
  AO7 U3036 ( .A(n4920), .B(n4457), .C(n4269), .Z(n1186) );
  NR3 U3037 ( .A(n4246), .B(n4900), .C(n4616), .Z(n1183) );
  ND2 U3038 ( .A(n3566), .B(n3565), .Z(n1182) );
  NR2 U3039 ( .A(n3927), .B(n3564), .Z(n3566) );
  MUX21L U3040 ( .A(n1181), .B(n3563), .S(n3954), .Z(n3565) );
  NR2 U3041 ( .A(n4004), .B(n3955), .Z(n3564) );
  ND2 U3042 ( .A(n2643), .B(n4055), .Z(n1180) );
  ND2 U3043 ( .A(n4896), .B(n4609), .Z(n2643) );
  EO U3044 ( .A(n4890), .B(n4240), .Z(n443) );
  MUX21L U3045 ( .A(n3839), .B(n3838), .S(n3924), .Z(n3847) );
  NR2 U3046 ( .A(n3997), .B(n3849), .Z(n3838) );
  NR3 U3047 ( .A(n3997), .B(n68), .C(n3958), .Z(n3839) );
  AN3 U3048 ( .A(n4038), .B(n3914), .C(n3951), .Z(n3587) );
  MUX21L U3049 ( .A(n3842), .B(n3843), .S(n3997), .Z(n3845) );
  ND2 U3050 ( .A(n2941), .B(n2940), .Z(n1168) );
  ND2 U3051 ( .A(n3958), .B(n3922), .Z(n3844) );
  MUX21L U3052 ( .A(n3598), .B(n3597), .S(n3955), .Z(n3603) );
  NR3 U3053 ( .A(n4000), .B(n71), .C(n3926), .Z(n3597) );
  NR2 U3054 ( .A(n4000), .B(n418), .Z(n3598) );
  MUX21L U3055 ( .A(n3599), .B(n3600), .S(n3926), .Z(n3601) );
  NR2 U3056 ( .A(n4001), .B(n3955), .Z(n3600) );
  AN3 U3057 ( .A(n3951), .B(n1165), .C(n3995), .Z(n3599) );
  NR2 U3058 ( .A(n4598), .B(n4269), .Z(n1165) );
  MUX21L U3059 ( .A(n3606), .B(n3607), .S(n3955), .Z(n3608) );
  NR2 U3060 ( .A(n3925), .B(n73), .Z(n3607) );
  NR3 U3061 ( .A(n3926), .B(n4001), .C(n74), .Z(n3606) );
  MUX21L U3062 ( .A(n3613), .B(n3612), .S(n3955), .Z(n3614) );
  ND2 U3063 ( .A(n3610), .B(n1160), .Z(n3612) );
  ND2 U3064 ( .A(n3611), .B(n1162), .Z(n3613) );
  NR2 U3065 ( .A(n4001), .B(n3925), .Z(n3610) );
  NR2 U3066 ( .A(n4001), .B(n3925), .Z(n3611) );
  NR2 U3067 ( .A(n3885), .B(n119), .Z(n3727) );
  ND3 U3068 ( .A(n4003), .B(n505), .C(n3956), .Z(n3670) );
  MUX41 U3069 ( .D0(n750), .D1(n733), .D2(n741), .D3(n725), .A(n3873), .B(
        n3882), .Z(N229) );
  MUX21L U3070 ( .A(n3453), .B(n3454), .S(n3958), .Z(n3462) );
  NR2 U3071 ( .A(n4016), .B(n413), .Z(n3454) );
  NR3 U3072 ( .A(n4016), .B(n433), .C(n3929), .Z(n3453) );
  ND2 U3073 ( .A(n3729), .B(n3728), .Z(N220) );
  AO2 U3074 ( .A(n3885), .B(n504), .C(n3885), .D(n3871), .Z(n3729) );
  MUX21L U3075 ( .A(n3727), .B(n502), .S(n3871), .Z(n3728) );
  ND3 U3076 ( .A(n3543), .B(n3542), .C(n3541), .Z(n504) );
  NR3 U3077 ( .A(n124), .B(n4010), .C(n3954), .Z(n3485) );
  ND2 U3078 ( .A(n4422), .B(n4862), .Z(n2160) );
  NR3 U3079 ( .A(n2324), .B(n3959), .C(n3930), .Z(n3373) );
  NR2 U3080 ( .A(n4003), .B(n3860), .Z(n3684) );
  IVP U3081 ( .A(n494), .Z(n3860) );
  AO4 U3082 ( .A(n4589), .B(n4239), .C(n4912), .D(n4239), .Z(n494) );
  NR2 U3083 ( .A(n3957), .B(n125), .Z(n3795) );
  ND2 U3084 ( .A(n4955), .B(n4633), .Z(n2323) );
  NR2 U3085 ( .A(n3424), .B(n3423), .Z(n3426) );
  NR2 U3086 ( .A(n4015), .B(n3959), .Z(n3424) );
  NR2 U3087 ( .A(n3959), .B(n433), .Z(n3423) );
  ND2 U3088 ( .A(n2618), .B(n2617), .Z(n647) );
  EO U3089 ( .A(n4884), .B(n4226), .Z(n645) );
  AO7 U3090 ( .A(n4940), .B(n4627), .C(n4135), .Z(n600) );
  ND2 U3091 ( .A(n1729), .B(n1728), .Z(n596) );
  ND3 U3092 ( .A(n2009), .B(n2008), .C(n2007), .Z(n602) );
  AN3 U3093 ( .A(n3953), .B(n669), .C(n3996), .Z(n3484) );
  ND3 U3094 ( .A(n2238), .B(n2237), .C(n2236), .Z(n669) );
  ND2 U3095 ( .A(n4637), .B(n4186), .Z(n2236) );
  ND2 U3096 ( .A(n4637), .B(n4952), .Z(n2238) );
  AN3 U3097 ( .A(n3951), .B(n420), .C(n3994), .Z(n3557) );
  MUX41 U3098 ( .D0(n720), .D1(n702), .D2(n711), .D3(n697), .A(n3873), .B(
        n3882), .Z(N228) );
  ND4 U3099 ( .A(n3722), .B(n3721), .C(n3720), .D(n3719), .Z(n697) );
  MUX41 U3100 ( .D0(n690), .D1(n672), .D2(n681), .D3(n666), .A(n3873), .B(
        n3881), .Z(N227) );
  MUX41 U3101 ( .D0(n659), .D1(n643), .D2(n650), .D3(n635), .A(n3873), .B(
        n3881), .Z(N226) );
  MUX41 U3102 ( .D0(n627), .D1(n612), .D2(n620), .D3(n603), .A(n3873), .B(
        n3881), .Z(N225) );
  MUX41 U3103 ( .D0(n595), .D1(n578), .D2(n587), .D3(n569), .A(n3873), .B(
        n3881), .Z(N224) );
  MUX41 U3104 ( .D0(n539), .D1(n524), .D2(n530), .D3(n522), .A(n3873), .B(
        n3881), .Z(N222) );
  ND2 U3105 ( .A(n3426), .B(n3425), .Z(n524) );
  ND2 U3106 ( .A(n3392), .B(n3391), .Z(n522) );
  MUX21L U3107 ( .A(n3678), .B(n498), .S(n3924), .Z(n3683) );
  NR3 U3108 ( .A(n4247), .B(n4897), .C(n4620), .Z(n498) );
  MUX21L U3109 ( .A(n3797), .B(n3796), .S(n3921), .Z(n3798) );
  AN3 U3110 ( .A(n3953), .B(n701), .C(n3997), .Z(n3797) );
  AN3 U3111 ( .A(n3996), .B(n3952), .C(n698), .Z(n3796) );
  ND2 U3112 ( .A(n2216), .B(n2215), .Z(n701) );
  MUX21L U3113 ( .A(n3711), .B(n3712), .S(n4004), .Z(n3722) );
  NR3 U3114 ( .A(n126), .B(n3957), .C(n3924), .Z(n3711) );
  ND2 U3115 ( .A(n3686), .B(n3685), .Z(n495) );
  AO6 U3116 ( .A(n4003), .B(n3956), .C(n3924), .Z(n3686) );
  MUX21L U3117 ( .A(n3684), .B(n493), .S(n3956), .Z(n3685) );
  ND2 U3118 ( .A(n3139), .B(n3138), .Z(n493) );
  AN3 U3119 ( .A(n545), .B(n3953), .C(n3994), .Z(n3457) );
  ND2 U3120 ( .A(n2249), .B(n4184), .Z(n545) );
  ND2 U3121 ( .A(n4953), .B(n4636), .Z(n2249) );
  AO4 U3122 ( .A(n4641), .B(n4298), .C(n4926), .D(n4298), .Z(n543) );
  NR3 U3123 ( .A(n4796), .B(n3959), .C(n3930), .Z(n3363) );
  NR2 U3124 ( .A(n3999), .B(n3957), .Z(n3790) );
  NR2 U3125 ( .A(n3999), .B(n3957), .Z(n3791) );
  NR2 U3126 ( .A(n3999), .B(n4641), .Z(n3793) );
  AN3 U3127 ( .A(n565), .B(n3915), .C(n3952), .Z(n3374) );
  ND3 U3128 ( .A(n4517), .B(n4833), .C(n4117), .Z(n565) );
  ND2 U3129 ( .A(n3954), .B(n496), .Z(n3479) );
  ND2 U3130 ( .A(n2253), .B(n4183), .Z(n496) );
  ND2 U3131 ( .A(n4953), .B(n4636), .Z(n2253) );
  ND2 U3132 ( .A(n3954), .B(n509), .Z(n3477) );
  ND2 U3133 ( .A(n2251), .B(n4184), .Z(n509) );
  ND2 U3134 ( .A(n4953), .B(n4636), .Z(n2251) );
  NR2 U3135 ( .A(n3999), .B(n3954), .Z(n3558) );
  AN3 U3136 ( .A(n721), .B(n3915), .C(n3951), .Z(n3364) );
  ND2 U3137 ( .A(n4116), .B(n4518), .Z(n721) );
  AN3 U3138 ( .A(n525), .B(n3914), .C(n3994), .Z(n3556) );
  ND3 U3139 ( .A(n4411), .B(n4860), .C(n4161), .Z(n525) );
  AN3 U3140 ( .A(n514), .B(n3995), .C(n3914), .Z(n3659) );
  ND3 U3141 ( .A(n4495), .B(n4752), .C(n4100), .Z(n514) );
  AN3 U3142 ( .A(n1643), .B(n3939), .C(n3996), .Z(n3819) );
  MUX21L U3143 ( .A(n2698), .B(n2697), .S(n4903), .Z(n1643) );
  ND2 U3144 ( .A(n4049), .B(n4478), .Z(n2698) );
  ND2 U3145 ( .A(n4606), .B(n4048), .Z(n2697) );
  AN3 U3146 ( .A(n1641), .B(n3939), .C(n3996), .Z(n3818) );
  NR2 U3147 ( .A(n4225), .B(n4856), .Z(n1641) );
  MUX21L U3148 ( .A(n3757), .B(n3756), .S(n3924), .Z(n3765) );
  NR2 U3149 ( .A(n4002), .B(n40), .Z(n3756) );
  AN3 U3150 ( .A(n1128), .B(n3972), .C(n3952), .Z(n3757) );
  AN3 U3151 ( .A(n1129), .B(n3940), .C(n3996), .Z(n3759) );
  MUX21L U3152 ( .A(n2334), .B(n4870), .S(n4633), .Z(n1129) );
  ND2 U3153 ( .A(n4288), .B(n4870), .Z(n2334) );
  IVP U3154 ( .A(n23), .Z(n3953) );
  IVP U3155 ( .A(n23), .Z(n3958) );
  IVP U3156 ( .A(n3939), .Z(n3969) );
  AN3 U3157 ( .A(n1072), .B(n3893), .C(n3994), .Z(n3544) );
  ND2 U3158 ( .A(n4898), .B(n2738), .Z(n1072) );
  ND2 U3159 ( .A(n4604), .B(n4242), .Z(n2738) );
  IVP U3160 ( .A(n3939), .Z(n3964) );
  IVP U3161 ( .A(n3943), .Z(n3955) );
  IVP U3162 ( .A(n3944), .Z(n3957) );
  IVP U3163 ( .A(n23), .Z(n3952) );
  IVP U3164 ( .A(n3939), .Z(n3965) );
  IVP U3165 ( .A(n3892), .Z(n3921) );
  IVP U3166 ( .A(n3887), .Z(n3916) );
  IVP U3167 ( .A(n3887), .Z(n3919) );
  IVP U3168 ( .A(n3973), .Z(n3998) );
  IVP U3169 ( .A(n3893), .Z(n3923) );
  IVP U3170 ( .A(n3975), .Z(n3997) );
  IVP U3171 ( .A(n3974), .Z(n3996) );
  IVP U3172 ( .A(n3886), .Z(n3920) );
  IVP U3173 ( .A(n3974), .Z(n4002) );
  IVP U3174 ( .A(n3975), .Z(n4013) );
  NR2 U3175 ( .A(n3998), .B(n3892), .Z(n3814) );
  IVP U3176 ( .A(n3949), .Z(n3954) );
  IVP U3177 ( .A(n3975), .Z(n4008) );
  IVP U3178 ( .A(n3975), .Z(n4009) );
  IVP U3179 ( .A(n3888), .Z(n3924) );
  IVP U3180 ( .A(n3975), .Z(n4012) );
  ND4 U3181 ( .A(n3655), .B(n3654), .C(n3653), .D(n3652), .Z(n1051) );
  ND4 U3182 ( .A(n1049), .B(n3956), .C(n3892), .D(n3979), .Z(n3652) );
  MUX21L U3183 ( .A(n3651), .B(n3650), .S(n3956), .Z(n3653) );
  MUX21L U3184 ( .A(n3648), .B(n3649), .S(n3956), .Z(n3654) );
  AN3 U3185 ( .A(n1050), .B(n3891), .C(n3995), .Z(n3648) );
  ND2 U3186 ( .A(n3170), .B(n3169), .Z(n1050) );
  ND3 U3187 ( .A(n4584), .B(n4086), .C(n4908), .Z(n3169) );
  MUX21L U3188 ( .A(n3167), .B(n3168), .S(n4584), .Z(n3170) );
  MUX21L U3189 ( .A(n3646), .B(n3647), .S(n4002), .Z(n3655) );
  AN3 U3190 ( .A(n1047), .B(n3944), .C(n3913), .Z(n3646) );
  AN3 U3191 ( .A(n1046), .B(n3944), .C(n3914), .Z(n3647) );
  ND2 U3192 ( .A(n4271), .B(n4735), .Z(n1047) );
  IVP U3193 ( .A(n3972), .Z(n3994) );
  IVP U3194 ( .A(n3888), .Z(n3927) );
  IVP U3195 ( .A(n3973), .Z(n3999) );
  IVP U3196 ( .A(n26), .Z(n3871) );
  AN3 U3197 ( .A(n1530), .B(n3979), .C(n3915), .Z(n3771) );
  MUX21L U3198 ( .A(n2056), .B(n4927), .S(n4299), .Z(n1530) );
  ND2 U3199 ( .A(n4927), .B(n4640), .Z(n2056) );
  AN3 U3200 ( .A(n1048), .B(n3889), .C(n3995), .Z(n3650) );
  MUX21L U3201 ( .A(n4206), .B(n4452), .S(n4922), .Z(n1048) );
  IVP U3202 ( .A(n3939), .Z(n3968) );
  IVP U3203 ( .A(n3945), .Z(n3956) );
  IVP U3204 ( .A(n3867), .Z(n3872) );
  IVP U3205 ( .A(n24), .Z(n3884) );
  IVP U3206 ( .A(n3886), .Z(n3914) );
  ND4 U3207 ( .A(n3336), .B(n3335), .C(n3334), .D(n3333), .Z(n992) );
  ND4 U3208 ( .A(n990), .B(n3960), .C(n3912), .D(n3992), .Z(n3333) );
  MUX21L U3209 ( .A(n3327), .B(n3328), .S(n4014), .Z(n3336) );
  MUX21L U3210 ( .A(n3329), .B(n3330), .S(n4014), .Z(n3335) );
  MUX21L U3211 ( .A(n3332), .B(n3331), .S(n3931), .Z(n3334) );
  NR3 U3212 ( .A(n44), .B(n4014), .C(n3960), .Z(n3332) );
  AN3 U3213 ( .A(n988), .B(n3942), .C(n3995), .Z(n3331) );
  IVP U3214 ( .A(n3879), .Z(n3883) );
  IVP U3215 ( .A(n3888), .Z(n3925) );
  IVP U3216 ( .A(n3979), .Z(n3995) );
  AN3 U3217 ( .A(n989), .B(n3887), .C(n3951), .Z(n3330) );
  MUX21L U3218 ( .A(n4825), .B(n1837), .S(n4630), .Z(n989) );
  ND2 U3219 ( .A(n4126), .B(n4825), .Z(n1837) );
  IVP U3220 ( .A(n3887), .Z(n3917) );
  ND4 U3221 ( .A(n3439), .B(n3438), .C(n3437), .D(n3436), .Z(n971) );
  ND4 U3222 ( .A(n968), .B(n3959), .C(n3907), .D(n3988), .Z(n3436) );
  MUX21L U3223 ( .A(n3432), .B(n3433), .S(n3959), .Z(n3438) );
  MUX21L U3224 ( .A(n3430), .B(n3431), .S(n4015), .Z(n3439) );
  AN3 U3225 ( .A(n1533), .B(n3980), .C(n3952), .Z(n3768) );
  ND2 U3226 ( .A(n4557), .B(n4871), .Z(n1533) );
  AN3 U3227 ( .A(n966), .B(n3945), .C(n3915), .Z(n3430) );
  ND2 U3228 ( .A(n2153), .B(n2152), .Z(n966) );
  ND2 U3229 ( .A(n4950), .B(n4423), .Z(n2152) );
  MUX21L U3230 ( .A(n2151), .B(n4138), .S(n4949), .Z(n2153) );
  MUX21L U3231 ( .A(n3435), .B(n3434), .S(n3959), .Z(n3437) );
  NR3 U3232 ( .A(n3929), .B(n4016), .C(n3854), .Z(n3435) );
  AN3 U3233 ( .A(n967), .B(n3889), .C(n3994), .Z(n3434) );
  IVP U3234 ( .A(n970), .Z(n3854) );
  MUX21L U3235 ( .A(n3703), .B(n3704), .S(n4004), .Z(n3708) );
  AN3 U3236 ( .A(n4384), .B(n3948), .C(n3914), .Z(n3703) );
  ND2 U3237 ( .A(n1841), .B(n1840), .Z(n960) );
  IVP U3238 ( .A(n3947), .Z(n3960) );
  IVP U3239 ( .A(n3973), .Z(n4000) );
  IVP U3240 ( .A(n3973), .Z(n4001) );
  IVP U3241 ( .A(n3886), .Z(n3915) );
  AN3 U3242 ( .A(n4733), .B(n3949), .C(n3916), .Z(n3327) );
  AN3 U3243 ( .A(n965), .B(n3941), .C(n3915), .Z(n3431) );
  AO7 U3244 ( .A(n4930), .B(n4190), .C(n4578), .Z(n965) );
  AN3 U3245 ( .A(n969), .B(n3889), .C(n3994), .Z(n3432) );
  MUX21L U3246 ( .A(n4868), .B(n4420), .S(n4289), .Z(n969) );
  AN3 U3247 ( .A(n961), .B(n3977), .C(n3952), .Z(n3701) );
  ND2 U3248 ( .A(n1908), .B(n1907), .Z(n961) );
  ND2 U3249 ( .A(n4939), .B(n4529), .Z(n1907) );
  MUX21L U3250 ( .A(n1906), .B(n4134), .S(n4939), .Z(n1908) );
  AN3 U3251 ( .A(n962), .B(n3948), .C(n3995), .Z(n3705) );
  EN U3252 ( .A(n4885), .B(n4293), .Z(n962) );
  IVP U3253 ( .A(n3889), .Z(n3931) );
  IVP U3254 ( .A(n3976), .Z(n4014) );
  IVP U3255 ( .A(n3974), .Z(n4007) );
  IVP U3256 ( .A(n3946), .Z(n3959) );
  IVP U3257 ( .A(n3975), .Z(n4011) );
  IVP U3258 ( .A(n3974), .Z(n4004) );
  IVP U3259 ( .A(n3880), .Z(n3882) );
  IVP U3260 ( .A(n3943), .Z(n3951) );
  AN3 U3261 ( .A(n939), .B(n3940), .C(n3996), .Z(n3747) );
  ND2 U3262 ( .A(n2315), .B(n2314), .Z(n939) );
  ND2 U3263 ( .A(n4634), .B(n4871), .Z(n2314) );
  MUX21L U3264 ( .A(n2313), .B(n4177), .S(n4634), .Z(n2315) );
  IVP U3265 ( .A(n3910), .Z(n3922) );
  IVP U3266 ( .A(n3889), .Z(n3929) );
  IVP U3267 ( .A(n3976), .Z(n4015) );
  IVP U3268 ( .A(n3976), .Z(n4016) );
  MUX21L U3269 ( .A(n3692), .B(n3691), .S(n3923), .Z(n3696) );
  AN3 U3270 ( .A(n1424), .B(n3977), .C(n3952), .Z(n3692) );
  EN U3271 ( .A(n4884), .B(n4627), .Z(n1424) );
  IVP U3272 ( .A(n3939), .Z(n3967) );
  IVP U3273 ( .A(n3974), .Z(n4003) );
  NR2 U3274 ( .A(n4004), .B(n3893), .Z(n3742) );
  ND4 U3275 ( .A(n3789), .B(n3788), .C(n3787), .D(n3786), .Z(n913) );
  MUX21L U3276 ( .A(n3781), .B(n3780), .S(n3923), .Z(n3789) );
  MUX21L U3277 ( .A(n3783), .B(n3782), .S(n3921), .Z(n3788) );
  AO2 U3278 ( .A(n3779), .B(n3892), .C(n3778), .D(n911), .Z(n3787) );
  AN3 U3279 ( .A(n4210), .B(n3940), .C(n3996), .Z(n3746) );
  MUX21L U3280 ( .A(n3806), .B(n3807), .S(n3999), .Z(n3811) );
  AN3 U3281 ( .A(n916), .B(n3940), .C(n3916), .Z(n3806) );
  AN3 U3282 ( .A(n4562), .B(n4208), .C(n4890), .Z(n917) );
  IVP U3283 ( .A(n3939), .Z(n3963) );
  IVP U3284 ( .A(n3887), .Z(n3918) );
  ND4 U3285 ( .A(n3402), .B(n3401), .C(n3400), .D(n3399), .Z(n1395) );
  ND4 U3286 ( .A(n1394), .B(n3959), .C(n3908), .D(n3989), .Z(n3399) );
  MUX21L U3287 ( .A(n3395), .B(n3396), .S(n4015), .Z(n3401) );
  MUX21L U3288 ( .A(n3398), .B(n3397), .S(n3959), .Z(n3400) );
  AN3 U3289 ( .A(n919), .B(n3940), .C(n3997), .Z(n3808) );
  MUX21L U3290 ( .A(n4217), .B(n4897), .S(n4605), .Z(n919) );
  AN3 U3291 ( .A(n918), .B(n3976), .C(n3953), .Z(n3804) );
  MUX21L U3292 ( .A(n4898), .B(n4608), .S(n4214), .Z(n918) );
  AN3 U3293 ( .A(n910), .B(n3940), .C(n3996), .Z(n3782) );
  EO U3294 ( .A(n4887), .B(n4280), .Z(n910) );
  MUX21L U3295 ( .A(n3393), .B(n3394), .S(n4015), .Z(n3402) );
  AN3 U3296 ( .A(n1392), .B(n3946), .C(n3915), .Z(n3393) );
  AN3 U3297 ( .A(n1391), .B(n3942), .C(n3915), .Z(n3394) );
  MUX21L U3298 ( .A(n4430), .B(n1799), .S(n4936), .Z(n1392) );
  AN3 U3299 ( .A(n1393), .B(n3888), .C(n3994), .Z(n3397) );
  ND2 U3300 ( .A(n1885), .B(n1884), .Z(n1393) );
  ND2 U3301 ( .A(n4258), .B(n4628), .Z(n1884) );
  MUX21L U3302 ( .A(n1883), .B(n4823), .S(n4629), .Z(n1885) );
  MUX21L U3303 ( .A(n3830), .B(n3831), .S(n3922), .Z(n3835) );
  AN3 U3304 ( .A(n887), .B(n3976), .C(n3953), .Z(n3831) );
  ND2 U3305 ( .A(n2710), .B(n2709), .Z(n890) );
  NR2 U3306 ( .A(n3923), .B(n3977), .Z(n3687) );
  AN3 U3307 ( .A(n4734), .B(n3978), .C(n3953), .Z(n3780) );
  IVP U3308 ( .A(n3975), .Z(n4010) );
  IVP U3309 ( .A(n3889), .Z(n3930) );
  NR2 U3310 ( .A(n3925), .B(n3947), .Z(n3827) );
  ND4 U3311 ( .A(n3584), .B(n3583), .C(n3582), .D(n3581), .Z(n1358) );
  ND4 U3312 ( .A(n1357), .B(n3955), .C(n3901), .D(n3983), .Z(n3581) );
  MUX21L U3313 ( .A(n3577), .B(n3578), .S(n4000), .Z(n3583) );
  MUX21L U3314 ( .A(n3575), .B(n3576), .S(n4000), .Z(n3584) );
  ND4 U3315 ( .A(n3346), .B(n3345), .C(n3344), .D(n3343), .Z(n849) );
  ND4 U3316 ( .A(n848), .B(n3960), .C(n3911), .D(n3991), .Z(n3343) );
  MUX21L U3317 ( .A(n3339), .B(n3340), .S(n4014), .Z(n3345) );
  MUX21L U3318 ( .A(n3337), .B(n3338), .S(n4014), .Z(n3346) );
  AN3 U3319 ( .A(n1355), .B(n3941), .C(n3914), .Z(n3575) );
  MUX21L U3320 ( .A(n2952), .B(n2951), .S(n4917), .Z(n1355) );
  ND2 U3321 ( .A(n4149), .B(n4507), .Z(n2952) );
  ND2 U3322 ( .A(n4273), .B(n4507), .Z(n2951) );
  AN3 U3323 ( .A(n847), .B(n3887), .C(n3951), .Z(n3340) );
  AO7 U3324 ( .A(n4937), .B(n4630), .C(n4260), .Z(n847) );
  MUX21L U3325 ( .A(n3580), .B(n3579), .S(n3926), .Z(n3582) );
  NR3 U3326 ( .A(n52), .B(n4000), .C(n3955), .Z(n3580) );
  AN3 U3327 ( .A(n1354), .B(n3941), .C(n3995), .Z(n3579) );
  MUX21L U3328 ( .A(n3342), .B(n3341), .S(n3931), .Z(n3344) );
  AN3 U3329 ( .A(n846), .B(n3941), .C(n3994), .Z(n3341) );
  NR3 U3330 ( .A(n54), .B(n4014), .C(n3960), .Z(n3342) );
  NR2 U3331 ( .A(n4574), .B(n4265), .Z(n846) );
  IVP U3332 ( .A(n3939), .Z(n3966) );
  AN3 U3333 ( .A(n1356), .B(n3911), .C(n3951), .Z(n3578) );
  AO7 U3334 ( .A(n4267), .B(n4770), .C(n3045), .Z(n1356) );
  ND2 U3335 ( .A(n4921), .B(n4599), .Z(n3045) );
  AN3 U3336 ( .A(n4210), .B(n3948), .C(n3916), .Z(n3337) );
  ND4 U3337 ( .A(n3308), .B(n3307), .C(n3306), .D(n3305), .Z(n1303) );
  MUX21L U3338 ( .A(n3304), .B(n3303), .S(n3931), .Z(n3306) );
  ND4 U3339 ( .A(n1302), .B(n3960), .C(n3904), .D(n3980), .Z(n3305) );
  MUX21L U3340 ( .A(n3299), .B(n3300), .S(n4013), .Z(n3308) );
  MUX21L U3341 ( .A(n3301), .B(n3302), .S(n4013), .Z(n3307) );
  AN3 U3342 ( .A(n1298), .B(n3916), .C(n3951), .Z(n3301) );
  AN3 U3343 ( .A(n1301), .B(n3886), .C(n3951), .Z(n3302) );
  ND3 U3344 ( .A(n4518), .B(n4833), .C(n4116), .Z(n1298) );
  IVP U3345 ( .A(n3974), .Z(n4006) );
  AN3 U3346 ( .A(n1300), .B(n3941), .C(n3916), .Z(n3299) );
  ND2 U3347 ( .A(n1829), .B(n1828), .Z(n1300) );
  ND2 U3348 ( .A(n4937), .B(n4261), .Z(n1829) );
  ND2 U3349 ( .A(n4631), .B(n4261), .Z(n1828) );
  AN3 U3350 ( .A(n1299), .B(n3950), .C(n3995), .Z(n3303) );
  AO4 U3351 ( .A(n4574), .B(n4265), .C(n4935), .D(n4265), .Z(n1299) );
  IVP U3352 ( .A(n3939), .Z(n3962) );
  IVP U3353 ( .A(n3870), .Z(n3873) );
  IVP U3354 ( .A(n3888), .Z(n3926) );
  NR2 U3355 ( .A(n3960), .B(n3911), .Z(n3352) );
  ND4 U3356 ( .A(n3521), .B(n3520), .C(n3519), .D(n3518), .Z(n812) );
  MUX21L U3357 ( .A(n3517), .B(n3516), .S(n3928), .Z(n3519) );
  ND4 U3358 ( .A(n810), .B(n3954), .C(n3903), .D(n3985), .Z(n3518) );
  MUX21L U3359 ( .A(n3514), .B(n3515), .S(n3998), .Z(n3520) );
  ND4 U3360 ( .A(n3472), .B(n3471), .C(n3470), .D(n3469), .Z(n806) );
  ND3 U3361 ( .A(n805), .B(n3988), .C(n3906), .Z(n3469) );
  MUX21L U3362 ( .A(n3467), .B(n3468), .S(n3929), .Z(n3470) );
  MUX21L U3363 ( .A(n3465), .B(n3466), .S(n3958), .Z(n3471) );
  AN3 U3364 ( .A(n809), .B(n3891), .C(n3951), .Z(n3515) );
  ND2 U3365 ( .A(n2640), .B(n2639), .Z(n809) );
  ND2 U3366 ( .A(n4609), .B(n4214), .Z(n2639) );
  MUX21L U3367 ( .A(n2638), .B(n4214), .S(n4894), .Z(n2640) );
  AN3 U3368 ( .A(n804), .B(n3993), .C(n3952), .Z(n3467) );
  ND2 U3369 ( .A(n4638), .B(n4282), .Z(n804) );
  MUX21L U3370 ( .A(n3512), .B(n3513), .S(n3997), .Z(n3521) );
  NR3 U3371 ( .A(n57), .B(n3953), .C(n3928), .Z(n3513) );
  AN3 U3372 ( .A(n808), .B(n3943), .C(n3914), .Z(n3512) );
  MUX21L U3373 ( .A(n3463), .B(n3464), .S(n4016), .Z(n3472) );
  NR2 U3374 ( .A(n3958), .B(n3929), .Z(n3463) );
  AN3 U3375 ( .A(n803), .B(n3942), .C(n3915), .Z(n3464) );
  ND2 U3376 ( .A(n2143), .B(n4136), .Z(n803) );
  MUX21L U3377 ( .A(n3356), .B(n3357), .S(n3930), .Z(n3359) );
  AN3 U3378 ( .A(n3942), .B(n3981), .C(n4022), .Z(n3357) );
  ND2 U3379 ( .A(n1969), .B(n1968), .Z(n800) );
  NR2 U3380 ( .A(n3930), .B(n3949), .Z(n3351) );
  ND4 U3381 ( .A(n3531), .B(n3530), .C(n3529), .D(n3528), .Z(n790) );
  ND3 U3382 ( .A(n412), .B(n3948), .C(n3927), .Z(n3528) );
  MUX21L U3383 ( .A(n3522), .B(n3523), .S(n3953), .Z(n3531) );
  MUX21L U3384 ( .A(n3526), .B(n3527), .S(n3927), .Z(n3529) );
  ND3 U3385 ( .A(n1268), .B(n3950), .C(n3931), .Z(n3315) );
  ND2 U3386 ( .A(n1831), .B(n1830), .Z(n1268) );
  ND2 U3387 ( .A(n4937), .B(n4261), .Z(n1831) );
  ND2 U3388 ( .A(n4631), .B(n4261), .Z(n1830) );
  MUX21L U3389 ( .A(n3309), .B(n3310), .S(n3960), .Z(n3318) );
  NR3 U3390 ( .A(n58), .B(n4013), .C(n3931), .Z(n3309) );
  AN3 U3391 ( .A(n1267), .B(n3990), .C(n3916), .Z(n3310) );
  MUX21L U3392 ( .A(n3313), .B(n3314), .S(n3931), .Z(n3316) );
  NR2 U3393 ( .A(n3960), .B(n3992), .Z(n3314) );
  AN3 U3394 ( .A(n1269), .B(n3995), .C(n3951), .Z(n3313) );
  NR2 U3395 ( .A(n4631), .B(n4260), .Z(n1269) );
  MUX21L U3396 ( .A(n3311), .B(n3312), .S(n4013), .Z(n3317) );
  AN3 U3397 ( .A(n1270), .B(n3886), .C(n3951), .Z(n3311) );
  NR2 U3398 ( .A(n3960), .B(n408), .Z(n3312) );
  ND3 U3399 ( .A(n4532), .B(n4817), .C(n4206), .Z(n1270) );
  MUX21L U3400 ( .A(n3524), .B(n3525), .S(n3998), .Z(n3530) );
  AN3 U3401 ( .A(n789), .B(n3891), .C(n3951), .Z(n3524) );
  NR2 U3402 ( .A(n3953), .B(n409), .Z(n3525) );
  ND2 U3403 ( .A(n2690), .B(n2689), .Z(n789) );
  IVP U3404 ( .A(n3889), .Z(n3928) );
  AN3 U3405 ( .A(n4022), .B(n3942), .C(n3994), .Z(n3516) );
  AN3 U3406 ( .A(n787), .B(n3976), .C(n3914), .Z(n3523) );
  NR2 U3407 ( .A(n4591), .B(n4223), .Z(n787) );
  MUX21L U3408 ( .A(n3736), .B(n3737), .S(n3922), .Z(n3738) );
  AN3 U3409 ( .A(n1248), .B(n3940), .C(n3996), .Z(n3736) );
  AO4 U3410 ( .A(n4578), .B(n4279), .C(n4930), .D(n4279), .Z(n1245) );
  ND2 U3411 ( .A(n2144), .B(n4137), .Z(n785) );
  ND2 U3412 ( .A(n4931), .B(n4580), .Z(n2144) );
  ND2 U3413 ( .A(n3414), .B(n3413), .Z(N173) );
  ND3 U3414 ( .A(n773), .B(n3867), .C(n3884), .Z(n3413) );
  NR2 U3415 ( .A(n4016), .B(n3945), .Z(n3468) );
  ND3 U3416 ( .A(n3910), .B(n3949), .C(n783), .Z(n3361) );
  AO7 U3417 ( .A(n4923), .B(n4626), .C(n4292), .Z(n783) );
  ND2 U3418 ( .A(n3959), .B(n3911), .Z(n3358) );
  AO3 U3419 ( .A(n417), .B(n3538), .C(n3537), .D(n3536), .Z(n773) );
  ND2 U3420 ( .A(n3903), .B(n3945), .Z(n3538) );
  MUX21L U3421 ( .A(n3534), .B(n3535), .S(n3999), .Z(n3536) );
  NR2 U3422 ( .A(n3953), .B(n3985), .Z(n3527) );
  ND2 U3423 ( .A(n3948), .B(n3989), .Z(n3421) );
  ND2 U3424 ( .A(n772), .B(n3949), .Z(n3420) );
  AO4 U3425 ( .A(n4578), .B(n4280), .C(n4930), .D(n4280), .Z(n772) );
  AN3 U3426 ( .A(n4210), .B(n3977), .C(n3952), .Z(n3732) );
  MUX21L U3427 ( .A(n3319), .B(n3320), .S(n4014), .Z(n3324) );
  NR2 U3428 ( .A(n3931), .B(n3950), .Z(n3320) );
  NR3 U3429 ( .A(n413), .B(n3960), .C(n3931), .Z(n3319) );
  ND2 U3430 ( .A(n3726), .B(n3866), .Z(N172) );
  MUX21L U3431 ( .A(n771), .B(n765), .S(n3885), .Z(n3726) );
  ND4 U3432 ( .A(n3628), .B(n3627), .C(n3626), .D(n3625), .Z(n771) );
  ND4 U3433 ( .A(n770), .B(n3955), .C(n3897), .D(n3981), .Z(n3625) );
  MUX21L U3434 ( .A(n3619), .B(n3620), .S(n4001), .Z(n3628) );
  MUX21L U3435 ( .A(n3621), .B(n3622), .S(n4001), .Z(n3627) );
  AN3 U3436 ( .A(n1246), .B(n3940), .C(n3915), .Z(n3734) );
  ND2 U3437 ( .A(n4188), .B(n4547), .Z(n1246) );
  MUX21L U3438 ( .A(n3624), .B(n3623), .S(n3925), .Z(n3626) );
  NR3 U3439 ( .A(n3186), .B(n4002), .C(n3955), .Z(n3624) );
  AN3 U3440 ( .A(n767), .B(n3950), .C(n3995), .Z(n3623) );
  ND2 U3441 ( .A(n3416), .B(n3415), .Z(N171) );
  ND2 U3442 ( .A(n3885), .B(n3867), .Z(n3416) );
  NR2 U3443 ( .A(n3927), .B(n3950), .Z(n3535) );
  ND4 U3444 ( .A(n3499), .B(n3498), .C(n3497), .D(n3496), .Z(n1211) );
  MUX21L U3445 ( .A(n3495), .B(n3494), .S(n3928), .Z(n3497) );
  ND4 U3446 ( .A(n1210), .B(n3954), .C(n3905), .D(n3986), .Z(n3496) );
  MUX21L U3447 ( .A(n3490), .B(n3491), .S(n3997), .Z(n3499) );
  AN3 U3448 ( .A(n769), .B(n3891), .C(n3951), .Z(n3622) );
  NR2 U3449 ( .A(n4268), .B(n4455), .Z(n769) );
  AN3 U3450 ( .A(n768), .B(n3950), .C(n3920), .Z(n3619) );
  AO7 U3451 ( .A(n4918), .B(n4612), .C(n4272), .Z(n768) );
  ND3 U3452 ( .A(n3950), .B(n3991), .C(n3910), .Z(n3360) );
  ND2 U3453 ( .A(n764), .B(n3867), .Z(n3415) );
  ND3 U3454 ( .A(n3637), .B(n3636), .C(n3635), .Z(n764) );
  MUX21L U3455 ( .A(n3633), .B(n3634), .S(n3925), .Z(n3635) );
  MUX21L U3456 ( .A(n3629), .B(n3630), .S(n3925), .Z(n3636) );
  MUX21L U3457 ( .A(n3492), .B(n3493), .S(n3997), .Z(n3498) );
  AN3 U3458 ( .A(n1206), .B(n3914), .C(n3952), .Z(n3492) );
  AN3 U3459 ( .A(n1209), .B(n3890), .C(n3952), .Z(n3493) );
  NR2 U3460 ( .A(n4591), .B(n4223), .Z(n1206) );
  AO7 U3461 ( .A(n3849), .B(n3540), .C(n3539), .Z(n765) );
  ND2 U3462 ( .A(n3902), .B(n3985), .Z(n3540) );
  ND2 U3463 ( .A(n3903), .B(n3945), .Z(n3539) );
  AN3 U3464 ( .A(n1208), .B(n3941), .C(n3914), .Z(n3490) );
  NR3 U3465 ( .A(n4228), .B(n4947), .C(n4596), .Z(n1208) );
  AN3 U3466 ( .A(n763), .B(n3950), .C(n3995), .Z(n3629) );
  ND3 U3467 ( .A(n3180), .B(n3179), .C(n3178), .Z(n763) );
  ND2 U3468 ( .A(n4083), .B(n4441), .Z(n3179) );
  ND2 U3469 ( .A(n4909), .B(n4441), .Z(n3180) );
  ND2 U3470 ( .A(n3452), .B(n3451), .Z(n1205) );
  MUX21L U3471 ( .A(n3906), .B(n3450), .S(n3958), .Z(n3451) );
  MUX21L U3472 ( .A(n3449), .B(n3448), .S(n3929), .Z(n3452) );
  ND2 U3473 ( .A(n3406), .B(n3405), .Z(N118) );
  ND3 U3474 ( .A(n1194), .B(n3870), .C(n3884), .Z(n3405) );
  MUX21L U3475 ( .A(n3404), .B(n3403), .S(n3871), .Z(n3406) );
  IVP U3476 ( .A(n3880), .Z(n3885) );
  AO3 U3477 ( .A(n4003), .B(n3677), .C(n3892), .D(n3676), .Z(n760) );
  ND2 U3478 ( .A(n3944), .B(n759), .Z(n3677) );
  MUX21L U3479 ( .A(n3674), .B(n3675), .S(n3956), .Z(n3676) );
  ND2 U3480 ( .A(n3241), .B(n3240), .Z(n759) );
  AN3 U3481 ( .A(n1207), .B(n3941), .C(n3993), .Z(n3494) );
  ND3 U3482 ( .A(n4399), .B(n4853), .C(n4065), .Z(n1207) );
  ND2 U3483 ( .A(n3912), .B(n3950), .Z(n3325) );
  ND2 U3484 ( .A(n3912), .B(n3992), .Z(n3326) );
  MUX21L U3485 ( .A(n3408), .B(n3407), .S(n3884), .Z(N117) );
  ND2 U3486 ( .A(n1182), .B(n3870), .Z(n3407) );
  ND2 U3487 ( .A(n1190), .B(n3870), .Z(n3408) );
  ND2 U3488 ( .A(n3641), .B(n3640), .Z(n757) );
  ND2 U3489 ( .A(n3956), .B(n3896), .Z(n3640) );
  MUX21L U3490 ( .A(n3639), .B(n3638), .S(n4002), .Z(n3641) );
  NR2 U3491 ( .A(n3925), .B(n3859), .Z(n3638) );
  AN3 U3492 ( .A(n1193), .B(n3944), .C(n3994), .Z(n3500) );
  ND2 U3493 ( .A(n4044), .B(n4485), .Z(n1193) );
  MUX21L U3494 ( .A(n3410), .B(n3409), .S(n3884), .Z(N116) );
  ND2 U3495 ( .A(n1174), .B(n3870), .Z(n3409) );
  ND2 U3496 ( .A(n1179), .B(n3869), .Z(n3410) );
  ND4 U3497 ( .A(n3594), .B(n3593), .C(n3592), .D(n3591), .Z(n1179) );
  ND4 U3498 ( .A(n1178), .B(n3955), .C(n3901), .D(n3983), .Z(n3591) );
  MUX21L U3499 ( .A(n3587), .B(n3588), .S(n4000), .Z(n3593) );
  MUX21L U3500 ( .A(n3590), .B(n3589), .S(n3926), .Z(n3592) );
  MUX21L U3501 ( .A(n3585), .B(n3586), .S(n4000), .Z(n3594) );
  NR3 U3502 ( .A(n66), .B(n3955), .C(n3926), .Z(n3586) );
  AN3 U3503 ( .A(n1176), .B(n3941), .C(n3914), .Z(n3585) );
  AN3 U3504 ( .A(n1175), .B(n3941), .C(n3995), .Z(n3589) );
  ND2 U3505 ( .A(n2939), .B(n2938), .Z(n1175) );
  ND2 U3506 ( .A(n4916), .B(n4274), .Z(n2939) );
  ND2 U3507 ( .A(n4613), .B(n4274), .Z(n2938) );
  AN3 U3508 ( .A(n1177), .B(n3896), .C(n3951), .Z(n3588) );
  MUX21L U3509 ( .A(n4269), .B(n3005), .S(n4920), .Z(n1177) );
  ND2 U3510 ( .A(n4269), .B(n4457), .Z(n3005) );
  ND4 U3511 ( .A(n3847), .B(n3846), .C(n3845), .D(n3844), .Z(n1172) );
  ND3 U3512 ( .A(n3511), .B(n3510), .C(n3509), .Z(n1174) );
  ND2 U3513 ( .A(n3904), .B(n3986), .Z(n3511) );
  ND2 U3514 ( .A(n3904), .B(n3947), .Z(n3509) );
  ND2 U3515 ( .A(n1173), .B(n3898), .Z(n3510) );
  ND2 U3516 ( .A(n3643), .B(n3642), .Z(n755) );
  ND3 U3517 ( .A(n3895), .B(n3945), .C(n4002), .Z(n3642) );
  ND3 U3518 ( .A(n3896), .B(n3950), .C(n754), .Z(n3643) );
  AO4 U3519 ( .A(n4588), .B(n4239), .C(n4912), .D(n4588), .Z(n754) );
  MUX21L U3520 ( .A(n3840), .B(n3841), .S(n3958), .Z(n3846) );
  AN3 U3521 ( .A(n1171), .B(n3890), .C(n3996), .Z(n3840) );
  MUX21L U3522 ( .A(n4456), .B(n3006), .S(n4269), .Z(n1169) );
  ND3 U3523 ( .A(n3603), .B(n3602), .C(n3601), .Z(n1167) );
  ND3 U3524 ( .A(n4590), .B(n4073), .C(n4909), .Z(n753) );
  MUX21L U3525 ( .A(n3595), .B(n3596), .S(n3926), .Z(n3602) );
  NR2 U3526 ( .A(n3955), .B(n3849), .Z(n3596) );
  AN3 U3527 ( .A(n1166), .B(n3950), .C(n3995), .Z(n3595) );
  ND2 U3528 ( .A(n3246), .B(n3245), .Z(n752) );
  ND2 U3529 ( .A(n4076), .B(n4794), .Z(n3246) );
  AO2 U3530 ( .A(n3605), .B(n4001), .C(n3604), .D(n4001), .Z(n3609) );
  NR2 U3531 ( .A(n3926), .B(n3946), .Z(n3604) );
  NR2 U3532 ( .A(n3926), .B(n76), .Z(n3605) );
  ND2 U3533 ( .A(n3609), .B(n3608), .Z(n1164) );
  AN3 U3534 ( .A(n3865), .B(n3874), .C(n1163), .Z(n444) );
  NR2 U3535 ( .A(n4588), .B(n4239), .Z(n751) );
  MUX21L U3536 ( .A(n4584), .B(n4234), .S(n4908), .Z(n1161) );
  MUX21L U3537 ( .A(n3616), .B(n3615), .S(n4001), .Z(n1159) );
  ND3 U3538 ( .A(n3900), .B(n3950), .C(n1158), .Z(n3615) );
  ND2 U3539 ( .A(n3211), .B(n4079), .Z(n1158) );
  EO U3540 ( .A(n4892), .B(n4587), .Z(n3211) );
  MUX21L U3541 ( .A(n3618), .B(n3617), .S(n4001), .Z(n1157) );
  ND3 U3542 ( .A(n3899), .B(n3943), .C(n1156), .Z(n3618) );
  MUX21L U3543 ( .A(n4238), .B(n3226), .S(n4587), .Z(n1156) );
  ND2 U3544 ( .A(n4237), .B(n4790), .Z(n3226) );
  ND3 U3545 ( .A(n3899), .B(n3950), .C(n1155), .Z(n3617) );
  AO4 U3546 ( .A(n4584), .B(n4234), .C(n4908), .D(n4234), .Z(n1155) );
  ND3 U3547 ( .A(n3900), .B(n3944), .C(n4078), .Z(n3616) );
  ND2 U3548 ( .A(n3285), .B(n3284), .Z(n1154) );
  EN U3549 ( .A(n4890), .B(n4241), .Z(n3285) );
  EO U3550 ( .A(n4564), .B(n4241), .Z(n3284) );
  MUX21L U3551 ( .A(n4911), .B(n4587), .S(n4238), .Z(n1153) );
  ND2 U3552 ( .A(n3228), .B(n3227), .Z(n1152) );
  ND2 U3553 ( .A(n4078), .B(n4436), .Z(n3228) );
  ND2 U3554 ( .A(n4911), .B(n4077), .Z(n3227) );
  AO4 U3555 ( .A(n4587), .B(n4238), .C(n4911), .D(n4238), .Z(n1151) );
  NR2 U3556 ( .A(n4588), .B(n4238), .Z(n1150) );
  NR2 U3557 ( .A(n3871), .B(n122), .Z(n3572) );
  ND2 U3558 ( .A(n3923), .B(n3947), .Z(n3681) );
  ND4 U3559 ( .A(n3371), .B(n3370), .C(n3369), .D(n3368), .Z(n725) );
  MUX21L U3560 ( .A(n3362), .B(n3363), .S(n4014), .Z(n3371) );
  ND4 U3561 ( .A(n724), .B(n3959), .C(n3910), .D(n3991), .Z(n3368) );
  MUX21L U3562 ( .A(n3364), .B(n3365), .S(n4015), .Z(n3370) );
  ND4 U3563 ( .A(n3462), .B(n3461), .C(n3460), .D(n3459), .Z(n547) );
  ND3 U3564 ( .A(n544), .B(n3988), .C(n3929), .Z(n3459) );
  MUX21L U3565 ( .A(n3455), .B(n3456), .S(n3958), .Z(n3461) );
  MUX21L U3566 ( .A(n3457), .B(n3458), .S(n3929), .Z(n3460) );
  ND4 U3567 ( .A(n3665), .B(n3664), .C(n3663), .D(n3662), .Z(n520) );
  ND4 U3568 ( .A(n518), .B(n3956), .C(n3894), .D(n3978), .Z(n3662) );
  MUX21L U3569 ( .A(n3656), .B(n3657), .S(n4002), .Z(n3665) );
  MUX21L U3570 ( .A(n3658), .B(n3659), .S(n3956), .Z(n3664) );
  AN3 U3571 ( .A(n519), .B(n3891), .C(n3995), .Z(n3658) );
  ND2 U3572 ( .A(n3209), .B(n3208), .Z(n519) );
  ND2 U3573 ( .A(n4910), .B(n4237), .Z(n3208) );
  EO U3574 ( .A(n4564), .B(n4237), .Z(n3209) );
  ND3 U3575 ( .A(n500), .B(n3978), .C(n3945), .Z(n3680) );
  ND2 U3576 ( .A(n3298), .B(n4073), .Z(n500) );
  EO U3577 ( .A(n4890), .B(n4601), .Z(n3298) );
  MUX41 U3578 ( .D0(n564), .D1(n547), .D2(n555), .D3(n542), .A(n3873), .B(
        n3881), .Z(N223) );
  AO3 U3579 ( .A(n3909), .B(n3387), .C(n3386), .D(n3385), .Z(n542) );
  MUX41 U3580 ( .D0(n520), .D1(n510), .D2(n513), .D3(n128), .A(n3872), .B(
        n3881), .Z(N221) );
  AO7 U3581 ( .A(n3987), .B(n3477), .C(n3906), .Z(n510) );
  ND4 U3582 ( .A(n3571), .B(n3570), .C(n3569), .D(n3568), .Z(n513) );
  MUX21L U3583 ( .A(n3668), .B(n3669), .S(n4003), .Z(n3672) );
  NR2 U3584 ( .A(n3924), .B(n3950), .Z(n3669) );
  NR3 U3585 ( .A(n3924), .B(n3956), .C(n123), .Z(n3668) );
  MUX21L U3586 ( .A(n3666), .B(n3667), .S(n4003), .Z(n3673) );
  NR2 U3587 ( .A(n3924), .B(n3849), .Z(n3667) );
  AN3 U3588 ( .A(n506), .B(n3950), .C(n3914), .Z(n3666) );
  MUX21L U3589 ( .A(n3679), .B(n3978), .S(n3923), .Z(n3682) );
  ND2 U3590 ( .A(n3137), .B(n3136), .Z(n499) );
  ND2 U3591 ( .A(n4907), .B(n4232), .Z(n3137) );
  MUX21L U3592 ( .A(n3367), .B(n3366), .S(n3930), .Z(n3369) );
  AN3 U3593 ( .A(n722), .B(n3942), .C(n3994), .Z(n3366) );
  NR3 U3594 ( .A(n120), .B(n4015), .C(n3959), .Z(n3367) );
  ND2 U3595 ( .A(n1768), .B(n1767), .Z(n722) );
  MUX21L U3596 ( .A(n3661), .B(n3660), .S(n3956), .Z(n3663) );
  AN3 U3597 ( .A(n517), .B(n3890), .C(n3995), .Z(n3660) );
  NR3 U3598 ( .A(n3924), .B(n4003), .C(n121), .Z(n3661) );
  AO4 U3599 ( .A(n4599), .B(n4267), .C(n4921), .D(n4267), .Z(n517) );
  ND2 U3600 ( .A(n3574), .B(n3573), .Z(N219) );
  ND2 U3601 ( .A(n497), .B(n3871), .Z(n3573) );
  MUX21L U3602 ( .A(n3572), .B(n3871), .S(n3885), .Z(n3574) );
  AO7 U3603 ( .A(n3987), .B(n3479), .C(n3905), .Z(n497) );
  NR2 U3604 ( .A(n3390), .B(n3389), .Z(n3392) );
  NR2 U3605 ( .A(n3930), .B(n3990), .Z(n3390) );
  NR2 U3606 ( .A(n3930), .B(n508), .Z(n3389) );
  ND4 U3607 ( .A(n3801), .B(n3800), .C(n3799), .D(n3798), .Z(n702) );
  MUX21L U3608 ( .A(n3793), .B(n3792), .S(n3920), .Z(n3801) );
  AO2 U3609 ( .A(n3791), .B(n3893), .C(n3790), .D(n700), .Z(n3799) );
  MUX21L U3610 ( .A(n3795), .B(n3794), .S(n3922), .Z(n3800) );
  ND4 U3611 ( .A(n3489), .B(n3488), .C(n3487), .D(n3486), .Z(n672) );
  ND4 U3612 ( .A(n668), .B(n3954), .C(n3928), .D(n3986), .Z(n3486) );
  MUX21L U3613 ( .A(n3480), .B(n3481), .S(n4016), .Z(n3489) );
  MUX21L U3614 ( .A(n3484), .B(n3485), .S(n3928), .Z(n3487) );
  ND4 U3615 ( .A(n3381), .B(n3380), .C(n3379), .D(n3378), .Z(n569) );
  ND4 U3616 ( .A(n4242), .B(n3959), .C(n3909), .D(n3990), .Z(n3378) );
  MUX21L U3617 ( .A(n3372), .B(n3373), .S(n4015), .Z(n3381) );
  MUX21L U3618 ( .A(n3374), .B(n3375), .S(n4015), .Z(n3380) );
  ND4 U3619 ( .A(n3562), .B(n3561), .C(n3560), .D(n3559), .Z(n530) );
  MUX21L U3620 ( .A(n3555), .B(n3556), .S(n3954), .Z(n3561) );
  ND3 U3621 ( .A(n529), .B(n3984), .C(n3942), .Z(n3559) );
  MUX21L U3622 ( .A(n3557), .B(n3558), .S(n3927), .Z(n3560) );
  AN3 U3623 ( .A(n723), .B(n3909), .C(n3952), .Z(n3365) );
  ND2 U3624 ( .A(n1879), .B(n1878), .Z(n723) );
  ND2 U3625 ( .A(n1875), .B(n4938), .Z(n1878) );
  MUX21L U3626 ( .A(n1876), .B(n1877), .S(n4938), .Z(n1879) );
  AN3 U3627 ( .A(n699), .B(n3984), .C(n3953), .Z(n3792) );
  MUX21L U3628 ( .A(n2063), .B(n4928), .S(n4300), .Z(n699) );
  ND2 U3629 ( .A(n4928), .B(n4546), .Z(n2063) );
  AN3 U3630 ( .A(n670), .B(n3890), .C(n3953), .Z(n3480) );
  EO U3631 ( .A(n4566), .B(n4285), .Z(n670) );
  AN3 U3632 ( .A(n568), .B(n3909), .C(n3952), .Z(n3375) );
  AO4 U3633 ( .A(n4630), .B(n4260), .C(n4938), .D(n4260), .Z(n568) );
  AN3 U3634 ( .A(n516), .B(n3950), .C(n3914), .Z(n3656) );
  ND2 U3635 ( .A(n2994), .B(n4152), .Z(n516) );
  ND2 U3636 ( .A(n4919), .B(n4597), .Z(n2994) );
  ND3 U3637 ( .A(n507), .B(n3895), .C(n3956), .Z(n3671) );
  ND2 U3638 ( .A(n3135), .B(n3134), .Z(n507) );
  ND2 U3639 ( .A(n4907), .B(n4232), .Z(n3135) );
  ND2 U3640 ( .A(n4583), .B(n4232), .Z(n3134) );
  ND3 U3641 ( .A(n3429), .B(n3428), .C(n3427), .Z(n492) );
  ND2 U3642 ( .A(n3907), .B(n3989), .Z(n3429) );
  ND2 U3643 ( .A(n3908), .B(n3948), .Z(n3427) );
  ND2 U3644 ( .A(n491), .B(n3907), .Z(n3428) );
  MUX21L U3645 ( .A(n3715), .B(n3716), .S(n4004), .Z(n3720) );
  AN3 U3646 ( .A(n693), .B(n3940), .C(n3915), .Z(n3715) );
  ND3 U3647 ( .A(n1882), .B(n1881), .C(n1880), .Z(n694) );
  MUX21L U3648 ( .A(n3717), .B(n3718), .S(n3922), .Z(n3719) );
  AN3 U3649 ( .A(n696), .B(n3940), .C(n3996), .Z(n3717) );
  AO4 U3650 ( .A(n4575), .B(n4264), .C(n4935), .D(n4264), .Z(n692) );
  MUX21L U3651 ( .A(n3482), .B(n3483), .S(n3954), .Z(n3488) );
  AN3 U3652 ( .A(n671), .B(n3890), .C(n3993), .Z(n3482) );
  AN3 U3653 ( .A(n3993), .B(n3914), .C(n667), .Z(n3483) );
  ND2 U3654 ( .A(n4633), .B(n4288), .Z(n671) );
  MUX21L U3655 ( .A(n3377), .B(n3376), .S(n3930), .Z(n3379) );
  AN3 U3656 ( .A(n566), .B(n3941), .C(n3994), .Z(n3376) );
  NR3 U3657 ( .A(n127), .B(n4015), .C(n3959), .Z(n3377) );
  NR3 U3658 ( .A(n4264), .B(n4935), .C(n4575), .Z(n566) );
  MUX21L U3659 ( .A(n3382), .B(n3383), .S(n3959), .Z(n3386) );
  AN3 U3660 ( .A(n540), .B(n3973), .C(n3915), .Z(n3383) );
  NR2 U3661 ( .A(n3930), .B(n419), .Z(n3382) );
  NR3 U3662 ( .A(n4289), .B(n4933), .C(n4572), .Z(n540) );
  MUX21L U3663 ( .A(n3553), .B(n3554), .S(n3927), .Z(n3562) );
  AN3 U3664 ( .A(n527), .B(n3984), .C(n3951), .Z(n3553) );
  NR2 U3665 ( .A(n3954), .B(n3855), .Z(n3554) );
  AO4 U3666 ( .A(n4608), .B(n4215), .C(n4900), .D(n4215), .Z(n527) );
  MUX21L U3667 ( .A(n3567), .B(n3984), .S(n3927), .Z(n3568) );
  AN3 U3668 ( .A(n3953), .B(n420), .C(n3995), .Z(n3567) );
  ND2 U3669 ( .A(n3419), .B(n3418), .Z(N218) );
  MUX21L U3670 ( .A(n3417), .B(n3865), .S(n3885), .Z(n3419) );
  ND2 U3671 ( .A(n495), .B(n3865), .Z(n3418) );
  ND2 U3672 ( .A(n512), .B(n3943), .Z(n3570) );
  NR3 U3673 ( .A(n4218), .B(n4894), .C(n4605), .Z(n512) );
  AO2 U3674 ( .A(n511), .B(n3926), .C(n3926), .D(n3947), .Z(n3569) );
  NR3 U3675 ( .A(n4222), .B(n4941), .C(n4567), .Z(n511) );
  AN3 U3676 ( .A(n4884), .B(n3940), .C(n3997), .Z(n3794) );
  AN3 U3677 ( .A(n515), .B(n3950), .C(n3914), .Z(n3657) );
  AO7 U3678 ( .A(n4915), .B(n4615), .C(n4275), .Z(n515) );
  MUX21L U3679 ( .A(n3388), .B(n3909), .S(n3959), .Z(n3391) );
  AN3 U3680 ( .A(n521), .B(n3973), .C(n3915), .Z(n3388) );
  NR2 U3681 ( .A(n4576), .B(n4262), .Z(n521) );
  ND2 U3682 ( .A(n503), .B(n3901), .Z(n3542) );
  ND2 U3683 ( .A(n4610), .B(n4211), .Z(n503) );
  AO7 U3684 ( .A(n3987), .B(n3478), .C(n3905), .Z(n502) );
  ND2 U3685 ( .A(n3954), .B(n501), .Z(n3478) );
  ND2 U3686 ( .A(n2252), .B(n4183), .Z(n501) );
  ND2 U3687 ( .A(n4953), .B(n4636), .Z(n2252) );
  MUX21L U3688 ( .A(n3713), .B(n3714), .S(n3924), .Z(n3721) );
  AN3 U3689 ( .A(n695), .B(n3977), .C(n3952), .Z(n3713) );
  ND2 U3690 ( .A(n4116), .B(n4518), .Z(n691) );
  MUX21L U3691 ( .A(n3422), .B(n3946), .S(n3929), .Z(n3425) );
  AN3 U3692 ( .A(n3994), .B(n523), .C(n3952), .Z(n3422) );
  ND2 U3693 ( .A(n2250), .B(n4184), .Z(n523) );
  ND2 U3694 ( .A(n4953), .B(n4636), .Z(n2250) );
  ND3 U3695 ( .A(n4623), .B(n4295), .C(n4924), .Z(n508) );
  AN3 U3696 ( .A(n4563), .B(n3942), .C(n3915), .Z(n3362) );
  AN3 U3697 ( .A(n4397), .B(n3941), .C(n3914), .Z(n3481) );
  MUX21L U3698 ( .A(n3384), .B(n3948), .S(n4015), .Z(n3385) );
  AN3 U3699 ( .A(n4026), .B(n3888), .C(n3952), .Z(n3384) );
  AO7 U3700 ( .A(n3849), .B(n3645), .C(n3644), .Z(n490) );
  ND2 U3701 ( .A(n3894), .B(n3979), .Z(n3645) );
  IVP U3702 ( .A(n3939), .Z(n3961) );
  IVP U3703 ( .A(n3974), .Z(n4005) );
  AN3 U3704 ( .A(n567), .B(n3947), .C(n3915), .Z(n3372) );
  ND2 U3705 ( .A(n4125), .B(n4524), .Z(n567) );
  AN3 U3706 ( .A(n546), .B(n3890), .C(n3994), .Z(n3455) );
  ND3 U3707 ( .A(n4420), .B(n4867), .C(n4172), .Z(n546) );
  AN3 U3708 ( .A(n528), .B(n3891), .C(n3994), .Z(n3555) );
  ND3 U3709 ( .A(n4485), .B(n4759), .C(n4044), .Z(n528) );
  NR2 U3710 ( .A(n4016), .B(n3949), .Z(n3458) );
  ND2 U3711 ( .A(n541), .B(n3948), .Z(n3387) );
  ND2 U3712 ( .A(n4125), .B(n4525), .Z(n541) );
  ND2 U3713 ( .A(n3902), .B(n3943), .Z(n3541) );
  ND2 U3714 ( .A(n3902), .B(n3984), .Z(n3543) );
  ND2 U3715 ( .A(n3893), .B(n3946), .Z(n3644) );
  ND2 U3716 ( .A(n3942), .B(n3983), .Z(n3571) );
  IVP U3717 ( .A(LogIn2[44]), .Z(n3939) );
  IVP U3718 ( .A(n4959), .Z(n4964) );
  IVP U3719 ( .A(n4985), .Z(n4969) );
  IVP U3720 ( .A(n4960), .Z(n4961) );
  IVP U3721 ( .A(n4960), .Z(n4963) );
  IVP U3722 ( .A(n4959), .Z(n4966) );
  IVP U3723 ( .A(n4960), .Z(n4962) );
  IVP U3724 ( .A(n4959), .Z(n4965) );
  IVP U3725 ( .A(LogIn2[40]), .Z(n4968) );
  IVP U3726 ( .A(n4970), .Z(n4967) );
  IVP U3727 ( .A(n3971), .Z(n3940) );
  IVP U3728 ( .A(n3971), .Z(n3949) );
  IVP U3729 ( .A(n3970), .Z(n3942) );
  IVP U3730 ( .A(n3970), .Z(n3945) );
  IVP U3731 ( .A(n3959), .Z(n3941) );
  IVP U3732 ( .A(n3970), .Z(n3946) );
  IVP U3733 ( .A(n3970), .Z(n3947) );
  IVP U3734 ( .A(n3971), .Z(n3948) );
  IVP U3735 ( .A(n3971), .Z(n3950) );
  IVP U3736 ( .A(LogIn2[44]), .Z(n3943) );
  IVP U3737 ( .A(LogIn2[47]), .Z(n3867) );
  IVP U3738 ( .A(LogIn2[44]), .Z(n3944) );
  IVP U3739 ( .A(LogIn2[47]), .Z(n3870) );
  IVP U3740 ( .A(LogIn2[47]), .Z(n3866) );
  IVP U3741 ( .A(LogIn2[47]), .Z(n3869) );
  IVP U3742 ( .A(LogIn2[47]), .Z(n3865) );
  IVP U3743 ( .A(LogIn2[47]), .Z(n3868) );
  IVP U3744 ( .A(n5049), .Z(n5048) );
  IVP U3745 ( .A(n5049), .Z(n5046) );
  IVP U3746 ( .A(n5049), .Z(n5047) );
  IVP U3747 ( .A(n5053), .Z(n5031) );
  IVP U3748 ( .A(n5052), .Z(n5032) );
  IVP U3749 ( .A(n5052), .Z(n5033) );
  IVP U3750 ( .A(n5051), .Z(n5034) );
  IVP U3751 ( .A(n5053), .Z(n5030) );
  IVP U3752 ( .A(n5053), .Z(n5029) );
  IVP U3753 ( .A(n5051), .Z(n5035) );
  IVP U3754 ( .A(n5051), .Z(n5036) );
  IVP U3755 ( .A(n5051), .Z(n5037) );
  IVP U3756 ( .A(n5051), .Z(n5038) );
  IVP U3757 ( .A(n5050), .Z(n5039) );
  IVP U3758 ( .A(n5050), .Z(n5040) );
  IVP U3759 ( .A(n5050), .Z(n5041) );
  IVP U3760 ( .A(n5050), .Z(n5042) );
  IVP U3761 ( .A(n5050), .Z(n5043) );
  IVP U3762 ( .A(n5054), .Z(n5025) );
  IVP U3763 ( .A(n5054), .Z(n5026) );
  IVP U3764 ( .A(n5054), .Z(n5027) );
  IVP U3765 ( .A(n5054), .Z(n5028) );
  IVP U3766 ( .A(n5049), .Z(n5044) );
  IVP U3767 ( .A(n5049), .Z(n5045) );
  IVP U3768 ( .A(n4968), .Z(n4959) );
  IVP U3769 ( .A(n4969), .Z(n4960) );
  IVP U3770 ( .A(n3943), .Z(n3971) );
  IVP U3771 ( .A(n3944), .Z(n3970) );
  AO5 U3772 ( .A(n446), .B(n447), .C(n5062), .Z(n445) );
  FA1A U3773 ( .A(Term31[26]), .B(Term11[114]), .CI(
        \add_1_root_sub_1_root_add_225_2/carry[2] ), .CO(
        \add_1_root_sub_1_root_add_225_2/carry[3] ), .S(N280) );
  FA1A U3774 ( .A(Term31[24]), .B(Term11[112]), .CI(FractionBit[23]), .CO(
        \add_1_root_sub_1_root_add_225_2/carry[1] ), .S(N278) );
  FA1A U3775 ( .A(Term31[25]), .B(Term11[113]), .CI(
        \add_1_root_sub_1_root_add_225_2/carry[1] ), .CO(
        \add_1_root_sub_1_root_add_225_2/carry[2] ), .S(N279) );
  IV U3776 ( .A(n448), .Z(n449) );
  IV U3777 ( .A(n464), .Z(n465) );
  IV U3778 ( .A(n468), .Z(n469) );
  IV U3779 ( .A(n470), .Z(n471) );
  IV U3780 ( .A(n474), .Z(n475) );
  IV U3781 ( .A(n476), .Z(n477) );
  IV U3782 ( .A(n478), .Z(n479) );
  IV U3783 ( .A(n480), .Z(n481) );
  IV U3784 ( .A(n482), .Z(n483) );
  MUX81P U3785 ( .D0(n538), .D1(n534), .D2(n536), .D3(n532), .D4(n537), .D5(
        n533), .D6(n535), .D7(n531), .A(n3913), .B(n3969), .C(n3999), .Z(n539)
         );
  MUX81P U3786 ( .D0(n554), .D1(n4062), .D2(n552), .D3(n549), .D4(n553), .D5(
        n550), .D6(n551), .D7(n548), .A(n3917), .B(n3965), .C(n4016), .Z(n555)
         );
  MUX81P U3787 ( .D0(n563), .D1(n559), .D2(n561), .D3(n557), .D4(n562), .D5(
        n558), .D6(n560), .D7(n556), .A(n3917), .B(n3960), .C(n4004), .Z(n564)
         );
  MUX81P U3788 ( .D0(n577), .D1(n573), .D2(n575), .D3(n571), .D4(n576), .D5(
        n572), .D6(n574), .D7(n570), .A(n3917), .B(n3961), .C(n4004), .Z(n578)
         );
  MUX81P U3789 ( .D0(n586), .D1(n582), .D2(n584), .D3(n580), .D4(n585), .D5(
        n581), .D6(n583), .D7(n579), .A(n3917), .B(n3961), .C(n4004), .Z(n587)
         );
  MUX81P U3790 ( .D0(n594), .D1(n4932), .D2(n592), .D3(n589), .D4(n593), .D5(
        n590), .D6(n591), .D7(n588), .A(n3917), .B(n3961), .C(n4004), .Z(n595)
         );
  MUX81P U3791 ( .D0(n602), .D1(n598), .D2(n600), .D3(n596), .D4(n601), .D5(
        n597), .D6(n599), .D7(n4109), .A(n3917), .B(n3961), .C(n4004), .Z(n603) );
  MUX81P U3792 ( .D0(n611), .D1(n607), .D2(n609), .D3(n605), .D4(n610), .D5(
        n606), .D6(n608), .D7(n604), .A(n3917), .B(n3961), .C(n4005), .Z(n612)
         );
  MUX81P U3793 ( .D0(n4932), .D1(n616), .D2(n618), .D3(n614), .D4(n619), .D5(
        n615), .D6(n617), .D7(n613), .A(n3917), .B(n3961), .C(n4005), .Z(n620)
         );
  MUX81P U3794 ( .D0(n626), .D1(n420), .D2(n624), .D3(n621), .D4(n625), .D5(
        n622), .D6(n623), .D7(n4932), .A(n3917), .B(n3961), .C(n4005), .Z(n627) );
  MUX81P U3795 ( .D0(n634), .D1(n630), .D2(n632), .D3(n628), .D4(n633), .D5(
        n629), .D6(n631), .D7(n4521), .A(n3917), .B(n3961), .C(n4005), .Z(n635) );
  MUX81P U3796 ( .D0(n4931), .D1(n639), .D2(n641), .D3(n637), .D4(n642), .D5(
        n638), .D6(n640), .D7(n636), .A(n3917), .B(n3961), .C(n4005), .Z(n643)
         );
  MUX81P U3797 ( .D0(n420), .D1(n646), .D2(n648), .D3(n644), .D4(n649), .D5(
        n645), .D6(n647), .D7(n4931), .A(n3917), .B(n3961), .C(n4005), .Z(n650) );
  MUX81P U3798 ( .D0(n658), .D1(n654), .D2(n656), .D3(n652), .D4(n657), .D5(
        n653), .D6(n655), .D7(n651), .A(n3917), .B(n3961), .C(n4005), .Z(n659)
         );
  MUX81P U3799 ( .D0(n665), .D1(n661), .D2(n663), .D3(n660), .D4(n664), .D5(
        n4922), .D6(n662), .D7(n4839), .A(n3917), .B(n3961), .C(n4005), .Z(
        n666) );
  MUX81P U3800 ( .D0(n680), .D1(n676), .D2(n678), .D3(n674), .D4(n679), .D5(
        n675), .D6(n677), .D7(n673), .A(n3918), .B(n3962), .C(n4005), .Z(n681)
         );
  MUX81P U3801 ( .D0(n689), .D1(n685), .D2(n687), .D3(n683), .D4(n688), .D5(
        n684), .D6(n686), .D7(n682), .A(n3918), .B(n3962), .C(n4005), .Z(n690)
         );
  MUX81P U3802 ( .D0(n710), .D1(n706), .D2(n708), .D3(n704), .D4(n709), .D5(
        n705), .D6(n707), .D7(n703), .A(n3918), .B(n3962), .C(n4005), .Z(n711)
         );
  MUX81P U3803 ( .D0(n719), .D1(n715), .D2(n717), .D3(n713), .D4(n718), .D5(
        n714), .D6(n716), .D7(n712), .A(n3918), .B(n3962), .C(n4005), .Z(n720)
         );
  MUX81P U3804 ( .D0(n732), .D1(n729), .D2(n4931), .D3(n727), .D4(n731), .D5(
        n728), .D6(n730), .D7(n726), .A(n3918), .B(n3962), .C(n4006), .Z(n733)
         );
  MUX81P U3805 ( .D0(n740), .D1(n737), .D2(n739), .D3(n735), .D4(n434), .D5(
        n736), .D6(n738), .D7(n734), .A(n3918), .B(n3962), .C(n4006), .Z(n741)
         );
  MUX81P U3806 ( .D0(n749), .D1(n745), .D2(n747), .D3(n743), .D4(n748), .D5(
        n744), .D6(n746), .D7(n742), .A(n3918), .B(n3962), .C(n4006), .Z(n750)
         );
  MUX81P U3807 ( .D0(n781), .D1(n777), .D2(n779), .D3(n775), .D4(n780), .D5(
        n776), .D6(n778), .D7(n774), .A(n3918), .B(n3962), .C(n4006), .Z(n782)
         );
  MUX81P U3808 ( .D0(n798), .D1(n794), .D2(n796), .D3(n792), .D4(n797), .D5(
        n793), .D6(n795), .D7(n791), .A(n3918), .B(n3962), .C(n4006), .Z(n799)
         );
  MUX81P U3809 ( .D0(n819), .D1(n815), .D2(n817), .D3(n814), .D4(n818), .D5(
        n4932), .D6(n816), .D7(n813), .A(n3918), .B(n3962), .C(n4006), .Z(n820) );
  MUX81P U3810 ( .D0(n4170), .D1(n4138), .D2(n827), .D3(n825), .D4(n828), .D5(
        n826), .D6(n407), .D7(n824), .A(n3918), .B(n3962), .C(n4006), .Z(n829)
         );
  MUX81P U3811 ( .D0(n835), .D1(n4597), .D2(n833), .D3(n830), .D4(n834), .D5(
        n831), .D6(n832), .D7(n4165), .A(n3918), .B(n3962), .C(n4006), .Z(n836) );
  MUX81P U3812 ( .D0(n843), .D1(n839), .D2(n841), .D3(n4597), .D4(n842), .D5(
        n838), .D6(n840), .D7(n837), .A(n3918), .B(n3963), .C(n4006), .Z(n844)
         );
  MUX81P U3813 ( .D0(n4418), .D1(n853), .D2(n855), .D3(n851), .D4(n856), .D5(
        n852), .D6(n854), .D7(n850), .A(n3918), .B(n3963), .C(n4006), .Z(n857)
         );
  MUX81P U3814 ( .D0(n863), .D1(n860), .D2(n861), .D3(n858), .D4(n862), .D5(
        n859), .D6(n4932), .D7(n4412), .A(n3918), .B(n3963), .C(n4006), .Z(
        n864) );
  MUX81P U3815 ( .D0(n870), .D1(n866), .D2(n868), .D3(n4932), .D4(n869), .D5(
        n429), .D6(n867), .D7(n865), .A(n3918), .B(n3963), .C(n4006), .Z(n871)
         );
  MUX81P U3816 ( .D0(n878), .D1(n874), .D2(n876), .D3(n872), .D4(n877), .D5(
        n873), .D6(n875), .D7(n4108), .A(n3918), .B(n3963), .C(n4007), .Z(n879) );
  MUX81P U3817 ( .D0(n4840), .D1(n882), .D2(n884), .D3(n4639), .D4(n885), .D5(
        n881), .D6(n883), .D7(n880), .A(n3918), .B(n3963), .C(n4007), .Z(n886)
         );
  MUX81P U3818 ( .D0(n899), .D1(n895), .D2(n897), .D3(n894), .D4(n898), .D5(
        n427), .D6(n896), .D7(n893), .A(n3918), .B(n3963), .C(n4007), .Z(n900)
         );
  MUX81P U3819 ( .D0(n907), .D1(n903), .D2(n905), .D3(n901), .D4(n906), .D5(
        n902), .D6(n904), .D7(n4522), .A(n3918), .B(n3963), .C(n4007), .Z(n908) );
  MUX81P U3820 ( .D0(n927), .D1(n924), .D2(n426), .D3(n922), .D4(n926), .D5(
        n923), .D6(n925), .D7(n921), .A(n3918), .B(n3963), .C(n4007), .Z(n928)
         );
  MUX81P U3821 ( .D0(n935), .D1(n931), .D2(n933), .D3(n929), .D4(n934), .D5(
        n930), .D6(n932), .D7(n4838), .A(n3918), .B(n3963), .C(n4007), .Z(n936) );
  MUX81P U3822 ( .D0(n947), .D1(n944), .D2(n945), .D3(n942), .D4(n946), .D5(
        n943), .D6(n425), .D7(n941), .A(n3918), .B(n3963), .C(n4007), .Z(n948)
         );
  MUX81P U3823 ( .D0(n956), .D1(n952), .D2(n954), .D3(n950), .D4(n955), .D5(
        n951), .D6(n953), .D7(n949), .A(n3918), .B(n3963), .C(n4007), .Z(n957)
         );
  MUX81P U3824 ( .D0(n979), .D1(n975), .D2(n977), .D3(n973), .D4(n978), .D5(
        n974), .D6(n976), .D7(n972), .A(n3919), .B(n3964), .C(n4007), .Z(n980)
         );
  MUX81P U3825 ( .D0(n4435), .D1(n983), .D2(n984), .D3(n4617), .D4(n985), .D5(
        n982), .D6(n4254), .D7(n981), .A(n3919), .B(n3964), .C(n4007), .Z(n986) );
  MUX81P U3826 ( .D0(n1000), .D1(n996), .D2(n998), .D3(n994), .D4(n999), .D5(
        n995), .D6(n997), .D7(n993), .A(n3919), .B(n3964), .C(n4007), .Z(n1001) );
  MUX81P U3827 ( .D0(n1008), .D1(n1005), .D2(n1006), .D3(n1003), .D4(n1007), 
        .D5(n1004), .D6(n4931), .D7(n1002), .A(n3919), .B(n3964), .C(n4007), 
        .Z(n1009) );
  MUX81P U3828 ( .D0(n1016), .D1(n1013), .D2(n1015), .D3(n1011), .D4(n423), 
        .D5(n1012), .D6(n1014), .D7(n1010), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1017) );
  MUX81P U3829 ( .D0(n1025), .D1(n1021), .D2(n1023), .D3(n1019), .D4(n1024), 
        .D5(n1020), .D6(n1022), .D7(n1018), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1026) );
  MUX81P U3830 ( .D0(n1034), .D1(n1030), .D2(n1032), .D3(n1028), .D4(n1033), 
        .D5(n1029), .D6(n1031), .D7(n1027), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1035) );
  MUX81P U3831 ( .D0(n1043), .D1(n1039), .D2(n1041), .D3(n1037), .D4(n1042), 
        .D5(n1038), .D6(n1040), .D7(n1036), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1044) );
  MUX81P U3832 ( .D0(n1059), .D1(n1055), .D2(n1057), .D3(n1053), .D4(n1058), 
        .D5(n1054), .D6(n1056), .D7(n1052), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1060) );
  MUX81P U3833 ( .D0(n1068), .D1(n1064), .D2(n1066), .D3(n1062), .D4(n1067), 
        .D5(n1063), .D6(n1065), .D7(n1061), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1069) );
  MUX81P U3834 ( .D0(n1080), .D1(n1076), .D2(n1078), .D3(n1075), .D4(n1079), 
        .D5(n422), .D6(n1077), .D7(n1074), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1081) );
  MUX81P U3835 ( .D0(n1088), .D1(n1084), .D2(n1086), .D3(n1082), .D4(n1087), 
        .D5(n1083), .D6(n1085), .D7(n4522), .A(n3919), .B(n3964), .C(n4008), 
        .Z(n1089) );
  MUX81P U3836 ( .D0(n1097), .D1(n1093), .D2(n1095), .D3(n1091), .D4(n1096), 
        .D5(n1092), .D6(n1094), .D7(n1090), .A(n3919), .B(n3965), .C(n4008), 
        .Z(n1098) );
  MUX81P U3837 ( .D0(n1105), .D1(n1102), .D2(n412), .D3(n1100), .D4(n1104), 
        .D5(n1101), .D6(n1103), .D7(n1099), .A(n3919), .B(n3965), .C(n4008), 
        .Z(n1106) );
  MUX81P U3838 ( .D0(n1114), .D1(n1110), .D2(n1112), .D3(n1108), .D4(n1113), 
        .D5(n1109), .D6(n1111), .D7(n1107), .A(n3919), .B(n3965), .C(n4008), 
        .Z(n1115) );
  MUX81P U3839 ( .D0(n1123), .D1(n1119), .D2(n1121), .D3(n1117), .D4(n1122), 
        .D5(n1118), .D6(n1120), .D7(n1116), .A(n3919), .B(n3965), .C(n4008), 
        .Z(n1124) );
  MUX81P U3840 ( .D0(n1139), .D1(n1135), .D2(n1137), .D3(n1133), .D4(n1138), 
        .D5(n1134), .D6(n1136), .D7(n1132), .A(n3920), .B(n3965), .C(n4009), 
        .Z(n1140) );
  MUX81P U3841 ( .D0(n1148), .D1(n1144), .D2(n1146), .D3(n1142), .D4(n1147), 
        .D5(n1143), .D6(n1145), .D7(n1141), .A(n3919), .B(n3965), .C(n4009), 
        .Z(n1149) );
  MUX81P U3842 ( .D0(n1189), .D1(n1185), .D2(n1187), .D3(n4251), .D4(n1188), 
        .D5(n1184), .D6(n1186), .D7(n1183), .A(n3920), .B(n3965), .C(n4009), 
        .Z(n1190) );
  MUX81P U3843 ( .D0(n1202), .D1(n1198), .D2(n1200), .D3(n1196), .D4(n1201), 
        .D5(n1197), .D6(n1199), .D7(n1195), .A(n3919), .B(n3965), .C(n4009), 
        .Z(n1203) );
  MUX81P U3844 ( .D0(n1219), .D1(n1215), .D2(n1217), .D3(n1213), .D4(n1218), 
        .D5(n1214), .D6(n1216), .D7(n1212), .A(n3919), .B(n3965), .C(n4009), 
        .Z(n1220) );
  MUX81P U3845 ( .D0(n1231), .D1(n1227), .D2(n1229), .D3(n1225), .D4(n1230), 
        .D5(n1226), .D6(n1228), .D7(n1224), .A(n3920), .B(n3965), .C(n4009), 
        .Z(n1232) );
  MUX81P U3846 ( .D0(n1239), .D1(n432), .D2(n1237), .D3(n1234), .D4(n1238), 
        .D5(n1235), .D6(n1236), .D7(n1233), .A(n3920), .B(n3965), .C(n4009), 
        .Z(n1240) );
  MUX81P U3847 ( .D0(n1257), .D1(n1253), .D2(n1255), .D3(n1251), .D4(n1256), 
        .D5(n1252), .D6(n1254), .D7(n1250), .A(n3919), .B(n3966), .C(n4009), 
        .Z(n1258) );
  MUX81P U3848 ( .D0(n1265), .D1(n431), .D2(n1263), .D3(n1260), .D4(n1264), 
        .D5(n1261), .D6(n1262), .D7(n1259), .A(n3920), .B(n3966), .C(n4009), 
        .Z(n1266) );
  MUX81P U3849 ( .D0(n4419), .D1(n1275), .D2(n1277), .D3(n1273), .D4(n1278), 
        .D5(n1274), .D6(n1276), .D7(n1272), .A(n3920), .B(n3966), .C(n4009), 
        .Z(n1279) );
  MUX81P U3850 ( .D0(n1287), .D1(n1283), .D2(n1285), .D3(n1281), .D4(n1286), 
        .D5(n1282), .D6(n1284), .D7(n1280), .A(n3919), .B(n3966), .C(n4009), 
        .Z(n1288) );
  MUX81P U3851 ( .D0(n1296), .D1(n1292), .D2(n1294), .D3(n1290), .D4(n1295), 
        .D5(n1291), .D6(n1293), .D7(n1289), .A(n3920), .B(n3966), .C(n4009), 
        .Z(n1297) );
  MUX81P U3852 ( .D0(n1310), .D1(n4567), .D2(n1308), .D3(n1305), .D4(n1309), 
        .D5(n1306), .D6(n1307), .D7(n1304), .A(n3920), .B(n3966), .C(n4010), 
        .Z(n1311) );
  MUX81P U3853 ( .D0(n1319), .D1(n1315), .D2(n1317), .D3(n1313), .D4(n1318), 
        .D5(n1314), .D6(n1316), .D7(n1312), .A(n3919), .B(n3966), .C(n4010), 
        .Z(n1320) );
  MUX81P U3854 ( .D0(n1328), .D1(n1324), .D2(n1326), .D3(n1322), .D4(n1327), 
        .D5(n1323), .D6(n1325), .D7(n1321), .A(n3920), .B(n3966), .C(n4010), 
        .Z(n1329) );
  MUX81P U3855 ( .D0(n1336), .D1(n1332), .D2(n1334), .D3(n1330), .D4(n1335), 
        .D5(n1331), .D6(n1333), .D7(n4107), .A(n3920), .B(n3966), .C(n4010), 
        .Z(n1337) );
  MUX81P U3856 ( .D0(n1343), .D1(n4839), .D2(n1342), .D3(n1339), .D4(n4632), 
        .D5(n1340), .D6(n1341), .D7(n1338), .A(n3920), .B(n3966), .C(n4010), 
        .Z(n1344) );
  MUX81P U3857 ( .D0(n430), .D1(n1348), .D2(n1350), .D3(n1346), .D4(n1351), 
        .D5(n1347), .D6(n1349), .D7(n1345), .A(n3920), .B(n3966), .C(n4010), 
        .Z(n1352) );
  MUX81P U3858 ( .D0(n1364), .D1(n1361), .D2(n1363), .D3(n1359), .D4(n4931), 
        .D5(n1360), .D6(n1362), .D7(n4523), .A(n3920), .B(n3966), .C(n4010), 
        .Z(n1365) );
  MUX81P U3859 ( .D0(n1372), .D1(n4277), .D2(n1370), .D3(n1367), .D4(n1371), 
        .D5(n1368), .D6(n1369), .D7(n1366), .A(n3920), .B(n3967), .C(n4010), 
        .Z(n1373) );
  MUX81P U3860 ( .D0(n1380), .D1(n1376), .D2(n1378), .D3(n1374), .D4(n1379), 
        .D5(n1375), .D6(n1377), .D7(n428), .A(n3920), .B(n3967), .C(n4010), 
        .Z(n1381) );
  MUX81P U3861 ( .D0(n1388), .D1(n1384), .D2(n1386), .D3(n1382), .D4(n1387), 
        .D5(n1383), .D6(n1385), .D7(n4883), .A(n3920), .B(n3967), .C(n4010), 
        .Z(n1389) );
  MUX81P U3862 ( .D0(n1402), .D1(n4137), .D2(n1400), .D3(n1397), .D4(n1401), 
        .D5(n1398), .D6(n1399), .D7(n1396), .A(n3920), .B(n3967), .C(n4010), 
        .Z(n1403) );
  MUX81P U3863 ( .D0(n1410), .D1(n3071), .D2(n1408), .D3(n1405), .D4(n1409), 
        .D5(n1406), .D6(n1407), .D7(n1404), .A(n3920), .B(n3967), .C(n4011), 
        .Z(n1411) );
  MUX81P U3864 ( .D0(n1419), .D1(n1415), .D2(n1417), .D3(n1413), .D4(n1418), 
        .D5(n1414), .D6(n1416), .D7(n1412), .A(n3920), .B(n3967), .C(n4011), 
        .Z(n1420) );
  MUX81P U3865 ( .D0(n1433), .D1(n1429), .D2(n1431), .D3(n1427), .D4(n1432), 
        .D5(n1428), .D6(n1430), .D7(n4931), .A(n3919), .B(n3967), .C(n4011), 
        .Z(n1434) );
  MUX81P U3866 ( .D0(n1442), .D1(n1438), .D2(n1440), .D3(n1436), .D4(n1441), 
        .D5(n1437), .D6(n1439), .D7(n1435), .A(n3920), .B(n3967), .C(n4011), 
        .Z(n1443) );
  MUX81P U3867 ( .D0(n1451), .D1(n1447), .D2(n1449), .D3(n1445), .D4(n1450), 
        .D5(n1446), .D6(n1448), .D7(n1444), .A(n3920), .B(n3967), .C(n4011), 
        .Z(n1452) );
  MUX81P U3868 ( .D0(n1459), .D1(n1456), .D2(n4839), .D3(n1454), .D4(n1458), 
        .D5(n1455), .D6(n1457), .D7(n1453), .A(n3919), .B(n3967), .C(n4011), 
        .Z(n1460) );
  MUX81P U3869 ( .D0(n1468), .D1(n1464), .D2(n1466), .D3(n1462), .D4(n1467), 
        .D5(n1463), .D6(n1465), .D7(n1461), .A(n3917), .B(n3967), .C(n4011), 
        .Z(n1469) );
  MUX81P U3870 ( .D0(n1476), .D1(n1472), .D2(n1474), .D3(n1471), .D4(n1475), 
        .D5(n2541), .D6(n1473), .D7(n1470), .A(n3917), .B(n3967), .C(n4011), 
        .Z(n1477) );
  MUX81P U3871 ( .D0(n1484), .D1(n4571), .D2(n1482), .D3(n1479), .D4(n1483), 
        .D5(n1480), .D6(n1481), .D7(n1478), .A(n3917), .B(n3968), .C(n4011), 
        .Z(n1485) );
  MUX81P U3872 ( .D0(n1492), .D1(n1488), .D2(n1490), .D3(n1486), .D4(n1491), 
        .D5(n1487), .D6(n1489), .D7(n424), .A(n3917), .B(n3968), .C(n4011), 
        .Z(n1493) );
  MUX81P U3873 ( .D0(n1500), .D1(n1497), .D2(n1499), .D3(n1495), .D4(n4558), 
        .D5(n1496), .D6(n1498), .D7(n1494), .A(n3917), .B(n3968), .C(n4011), 
        .Z(n1501) );
  MUX81P U3874 ( .D0(n1509), .D1(n1505), .D2(n1507), .D3(n1503), .D4(n1508), 
        .D5(n1504), .D6(n1506), .D7(n1502), .A(n3917), .B(n3968), .C(n4011), 
        .Z(n1510) );
  MUX81P U3875 ( .D0(n1518), .D1(n1514), .D2(n1516), .D3(n1512), .D4(n1517), 
        .D5(n1513), .D6(n1515), .D7(n1511), .A(n3917), .B(n3968), .C(n4012), 
        .Z(n1519) );
  MUX81P U3876 ( .D0(n1527), .D1(n1523), .D2(n1525), .D3(n1521), .D4(n1526), 
        .D5(n1522), .D6(n1524), .D7(n1520), .A(n3917), .B(n3968), .C(n4012), 
        .Z(n1528) );
  MUX81P U3877 ( .D0(n1543), .D1(n1539), .D2(n1541), .D3(n1537), .D4(n1542), 
        .D5(n1538), .D6(n1540), .D7(n1536), .A(n3917), .B(n3968), .C(n4012), 
        .Z(n1544) );
  MUX81P U3878 ( .D0(n1552), .D1(n1548), .D2(n1550), .D3(n1546), .D4(n1551), 
        .D5(n1547), .D6(n1549), .D7(n1545), .A(n3916), .B(n3968), .C(n4012), 
        .Z(n1553) );
  MUX81P U3879 ( .D0(n1561), .D1(n1557), .D2(n1559), .D3(n1555), .D4(n1560), 
        .D5(n1556), .D6(n1558), .D7(n1554), .A(n3916), .B(n3968), .C(n4012), 
        .Z(n1562) );
  MUX81P U3880 ( .D0(n1570), .D1(n1566), .D2(n1568), .D3(n1564), .D4(n1569), 
        .D5(n1565), .D6(n1567), .D7(n1563), .A(n3916), .B(n3968), .C(n4012), 
        .Z(n1571) );
  MUX81P U3881 ( .D0(n1579), .D1(n1575), .D2(n1577), .D3(n1573), .D4(n1578), 
        .D5(n1574), .D6(n1576), .D7(n1572), .A(n3916), .B(n3968), .C(n4012), 
        .Z(n1580) );
  MUX81P U3882 ( .D0(n1588), .D1(n1584), .D2(n1586), .D3(n1582), .D4(n1587), 
        .D5(n1583), .D6(n1585), .D7(n1581), .A(n3916), .B(n3968), .C(n4012), 
        .Z(n1589) );
  MUX81P U3883 ( .D0(n1597), .D1(n1593), .D2(n1595), .D3(n1591), .D4(n1596), 
        .D5(n1592), .D6(n1594), .D7(n1590), .A(n3916), .B(n3969), .C(n4012), 
        .Z(n1598) );
  MUX81P U3884 ( .D0(n1606), .D1(n1602), .D2(n1604), .D3(n1600), .D4(n1605), 
        .D5(n1601), .D6(n1603), .D7(n1599), .A(n3916), .B(n3969), .C(n4012), 
        .Z(n1607) );
  MUX81P U3885 ( .D0(n4818), .D1(n424), .D2(n406), .D3(n1608), .D4(n1611), 
        .D5(n1609), .D6(n1610), .D7(n2556), .A(n3916), .B(n3969), .C(n4012), 
        .Z(n1612) );
  MUX81P U3886 ( .D0(n1620), .D1(n1616), .D2(n1618), .D3(n1614), .D4(n1619), 
        .D5(n1615), .D6(n1617), .D7(n1613), .A(n3916), .B(n3969), .C(n4012), 
        .Z(n1621) );
  MUX81P U3887 ( .D0(n1629), .D1(n1625), .D2(n1627), .D3(n1623), .D4(n1628), 
        .D5(n1624), .D6(n1626), .D7(n1622), .A(n3916), .B(n3969), .C(n4013), 
        .Z(n1630) );
  MUX81P U3888 ( .D0(n1638), .D1(n1634), .D2(n1636), .D3(n1632), .D4(n1637), 
        .D5(n1633), .D6(n1635), .D7(n1631), .A(n3916), .B(n3969), .C(n4013), 
        .Z(n1639) );
  MUX81P U3889 ( .D0(n1653), .D1(n1649), .D2(n1651), .D3(n1647), .D4(n1652), 
        .D5(n1648), .D6(n1650), .D7(n1646), .A(n3916), .B(n3969), .C(n4013), 
        .Z(n1654) );
  MUX81P U3890 ( .D0(n1662), .D1(n1658), .D2(n1660), .D3(n1656), .D4(n1661), 
        .D5(n1657), .D6(n1659), .D7(n1655), .A(n3916), .B(n3969), .C(n4013), 
        .Z(n1663) );
  MUX81P U3891 ( .D0(n1671), .D1(n1667), .D2(n1669), .D3(n1665), .D4(n1670), 
        .D5(n1666), .D6(n1668), .D7(n1664), .A(n3916), .B(n3969), .C(n4013), 
        .Z(n1672) );
  MUX81P U3892 ( .D0(n1679), .D1(n1676), .D2(n1678), .D3(n1674), .D4(n421), 
        .D5(n1675), .D6(n1677), .D7(n1673), .A(n3916), .B(n3969), .C(n4013), 
        .Z(n1680) );
  MUX81P U3893 ( .D0(n1688), .D1(n1684), .D2(n1686), .D3(n1682), .D4(n1687), 
        .D5(n1683), .D6(n1685), .D7(n1681), .A(n3916), .B(n3969), .C(n4013), 
        .Z(n1689) );
  AN2P U3894 ( .A(n4209), .B(n4890), .Z(n1702) );
  AN2P U3895 ( .A(n4566), .B(n4209), .Z(n1738) );
  AN2P U3896 ( .A(n4891), .B(n4209), .Z(n1757) );
  AN2P U3897 ( .A(n4891), .B(n4209), .Z(n1761) );
  AN2P U3898 ( .A(n4891), .B(n4565), .Z(n1765) );
  AN2P U3899 ( .A(n4891), .B(n4564), .Z(n1772) );
  AN2P U3900 ( .A(n4564), .B(n4208), .Z(n1778) );
  AN2P U3901 ( .A(n4892), .B(n4563), .Z(n1804) );
  AN2P U3902 ( .A(n4892), .B(n4563), .Z(n1813) );
  AN2P U3903 ( .A(n4892), .B(n4563), .Z(n1816) );
  AN2P U3904 ( .A(n4892), .B(n4210), .Z(n1838) );
  AN2P U3905 ( .A(n4892), .B(n4207), .Z(n1842) );
  AN2P U3906 ( .A(n4566), .B(n4208), .Z(n1877) );
  AN2P U3907 ( .A(n4564), .B(n4209), .Z(n1906) );
  AN2P U3908 ( .A(n4884), .B(n4209), .Z(n1933) );
  AN2P U3909 ( .A(n4884), .B(n4563), .Z(n1947) );
  AN2P U3910 ( .A(n4562), .B(n4208), .Z(n1981) );
  AN2P U3911 ( .A(n4207), .B(n4561), .Z(n1994) );
  AN2P U3912 ( .A(n4886), .B(n4208), .Z(n2029) );
  AN2P U3913 ( .A(n4886), .B(n4560), .Z(n2036) );
  AN2P U3914 ( .A(n4886), .B(n4560), .Z(n2039) );
  AN2P U3915 ( .A(n4887), .B(n4561), .Z(n2065) );
  AN2P U3916 ( .A(n4562), .B(n4209), .Z(n2072) );
  AN2P U3917 ( .A(n4208), .B(n4887), .Z(n2093) );
  AN2P U3918 ( .A(n4562), .B(n4887), .Z(n2109) );
  AN2P U3919 ( .A(n4887), .B(n4208), .Z(n2116) );
  AN2P U3920 ( .A(n4208), .B(n4888), .Z(n2121) );
  AN2P U3921 ( .A(n4888), .B(n4561), .Z(n2131) );
  AN2P U3922 ( .A(n4210), .B(n4888), .Z(n2145) );
  AN2P U3923 ( .A(n4560), .B(n4209), .Z(n2151) );
  AN2P U3924 ( .A(n4560), .B(n4208), .Z(n2175) );
  AN2P U3925 ( .A(n4889), .B(n4563), .Z(n2200) );
  AN2P U3926 ( .A(n4889), .B(n4563), .Z(n2205) );
  AN2P U3927 ( .A(n4889), .B(n4208), .Z(n2209) );
  AN2P U3928 ( .A(n4889), .B(n4564), .Z(n2213) );
  AN2P U3929 ( .A(n4889), .B(n4565), .Z(n2228) );
  AN2P U3930 ( .A(n4565), .B(n4208), .Z(n2233) );
  AN2P U3931 ( .A(n4564), .B(n4209), .Z(n2276) );
  AN2P U3932 ( .A(n4565), .B(n4209), .Z(n2289) );
  AN2P U3933 ( .A(n4887), .B(n4565), .Z(n2294) );
  AN2P U3934 ( .A(n4889), .B(n4210), .Z(n2308) );
  AN2P U3935 ( .A(n4889), .B(n4210), .Z(n2313) );
  AN2P U3936 ( .A(n4566), .B(n4210), .Z(n2324) );
  AN2P U3937 ( .A(n4565), .B(n4210), .Z(n2337) );
  AN2P U3938 ( .A(n4888), .B(n4210), .Z(n2364) );
  AN2P U3939 ( .A(n4209), .B(n4887), .Z(n2380) );
  AN2P U3940 ( .A(n4887), .B(n4565), .Z(n2386) );
  AN2P U3941 ( .A(n4565), .B(n4887), .Z(n2394) );
  AN2P U3942 ( .A(n4886), .B(n4208), .Z(n2424) );
  AN2P U3943 ( .A(n4886), .B(n4208), .Z(n2428) );
  AN2P U3944 ( .A(n4566), .B(n4208), .Z(n2435) );
  AN2P U3945 ( .A(n4566), .B(n4208), .Z(n2441) );
  AN2P U3946 ( .A(n4563), .B(n4208), .Z(n2507) );
  AN2P U3947 ( .A(n4892), .B(n4562), .Z(n2519) );
  AN2P U3948 ( .A(n4892), .B(n4561), .Z(n2541) );
  AN2P U3949 ( .A(n4561), .B(n4209), .Z(n2553) );
  AN2P U3950 ( .A(n4892), .B(n4561), .Z(n2556) );
  AN2P U3951 ( .A(n4892), .B(n4561), .Z(n2562) );
  AN2P U3952 ( .A(n4209), .B(n4891), .Z(n2582) );
  AN2P U3953 ( .A(n4210), .B(n4891), .Z(n2591) );
  AN2P U3954 ( .A(n4210), .B(n4891), .Z(n2597) );
  AN2P U3955 ( .A(n4563), .B(n4208), .Z(n2614) );
  AN2P U3956 ( .A(n4561), .B(n4207), .Z(n2655) );
  AN2P U3957 ( .A(n4891), .B(n4208), .Z(n2661) );
  AN2P U3958 ( .A(n4891), .B(n4560), .Z(n2670) );
  AN2P U3959 ( .A(n4560), .B(n4210), .Z(n2728) );
  AN2P U3960 ( .A(n4884), .B(n4561), .Z(n2734) );
  AN2P U3961 ( .A(n4885), .B(n4210), .Z(n2748) );
  AN2P U3962 ( .A(n4886), .B(n4209), .Z(n2757) );
  AN2P U3963 ( .A(n4886), .B(n4562), .Z(n2774) );
  AN2P U3964 ( .A(n4887), .B(n4562), .Z(n2790) );
  AN2P U3965 ( .A(n4562), .B(n4888), .Z(n2804) );
  AN2P U3966 ( .A(n4208), .B(n4564), .Z(n2855) );
  AN2P U3967 ( .A(n4889), .B(n4564), .Z(n2860) );
  AN2P U3968 ( .A(n4889), .B(n4564), .Z(n2865) );
  AN2P U3969 ( .A(n4564), .B(n4208), .Z(n2872) );
  AN2P U3970 ( .A(n4565), .B(n4889), .Z(n2888) );
  AN2P U3971 ( .A(n4565), .B(n4889), .Z(n2895) );
  AN2P U3972 ( .A(n4889), .B(n4208), .Z(n2905) );
  AN2P U3973 ( .A(n4207), .B(n4566), .Z(n2920) );
  AN2P U3974 ( .A(n4888), .B(n4208), .Z(n2956) );
  AN2P U3975 ( .A(n4887), .B(n4208), .Z(n2969) );
  AN2P U3976 ( .A(n4886), .B(n4209), .Z(n3015) );
  AN2P U3977 ( .A(n4886), .B(n4209), .Z(n3025) );
  AN2P U3978 ( .A(n4209), .B(n4560), .Z(n3040) );
  AN2P U3979 ( .A(n4885), .B(n4209), .Z(n3067) );
  AN2P U3980 ( .A(n4885), .B(n4561), .Z(n3071) );
  AN2P U3981 ( .A(n4885), .B(n4209), .Z(n3084) );
  AN2P U3982 ( .A(n4562), .B(n4885), .Z(n3093) );
  AN2P U3983 ( .A(n4884), .B(n4562), .Z(n3097) );
  AN2P U3984 ( .A(n4209), .B(n4562), .Z(n3103) );
  AN2P U3985 ( .A(n4562), .B(n4209), .Z(n3108) );
  AN2P U3986 ( .A(n4884), .B(n4562), .Z(n3114) );
  AN2P U3987 ( .A(n4893), .B(n4207), .Z(n3167) );
  AN2P U3988 ( .A(n4892), .B(n4207), .Z(n3186) );
  AN2P U3989 ( .A(n4891), .B(n4565), .Z(n3217) );
  AN2P U3990 ( .A(n4566), .B(n4891), .Z(n3253) );
  AN2P U3991 ( .A(n4566), .B(n4209), .Z(n3263) );
  AN2P U3992 ( .A(n4565), .B(n4209), .Z(n3275) );
  AN2P U3993 ( .A(n3951), .B(n1242), .Z(n3321) );
  AN2P U3994 ( .A(n821), .B(n3994), .Z(n3349) );
  AN2P U3995 ( .A(n3994), .B(n800), .Z(n3356) );
  AN2P U3996 ( .A(n3871), .B(n492), .Z(n3417) );
  AN2P U3997 ( .A(n3915), .B(n1222), .Z(n3444) );
  AN2P U3998 ( .A(n1204), .B(n3953), .Z(n3448) );
  AN2P U3999 ( .A(n3994), .B(n3915), .Z(n3450) );
  AN2P U4000 ( .A(n543), .B(n3915), .Z(n3456) );
  AN2P U4001 ( .A(n802), .B(n3915), .Z(n3466) );
  AN2P U4002 ( .A(n3993), .B(n785), .Z(n3473) );
  AN2P U4003 ( .A(n3994), .B(n1180), .Z(n3563) );
  OR2 U4004 ( .A(n79), .B(n3614), .Z(n1163) );
  AN2P U4005 ( .A(n3995), .B(n758), .Z(n3674) );
  AN2P U4006 ( .A(n3995), .B(n3951), .Z(n3678) );
  AN2P U4007 ( .A(n3951), .B(n499), .Z(n3679) );
  AN2P U4008 ( .A(n3995), .B(n3914), .Z(n3688) );
  AN2P U4009 ( .A(n1421), .B(n3952), .Z(n3691) );
  AN2P U4010 ( .A(n1423), .B(n3995), .Z(n3693) );
  AN2P U4011 ( .A(n3995), .B(n1422), .Z(n3694) );
  AN2P U4012 ( .A(n3952), .B(n3914), .Z(n3700) );
  AN2P U4013 ( .A(n958), .B(n3952), .Z(n3702) );
  AN2P U4014 ( .A(n3952), .B(n960), .Z(n3704) );
  AN2P U4015 ( .A(n3995), .B(n959), .Z(n3706) );
  AN2P U4016 ( .A(n3952), .B(n3914), .Z(n3712) );
  AN2P U4017 ( .A(n691), .B(n3952), .Z(n3714) );
  AN2P U4018 ( .A(n3952), .B(n694), .Z(n3716) );
  AN2P U4019 ( .A(n3996), .B(n692), .Z(n3718) );
  AN2P U4020 ( .A(n3952), .B(n3915), .Z(n3731) );
  AN2P U4021 ( .A(n1244), .B(n3952), .Z(n3733) );
  AN2P U4022 ( .A(n3952), .B(n1247), .Z(n3735) );
  AN2P U4023 ( .A(n3996), .B(n1245), .Z(n3737) );
  AN2P U4024 ( .A(n937), .B(n3952), .Z(n3748) );
  AN2P U4025 ( .A(n1531), .B(n3996), .Z(n3770) );
  AN2P U4026 ( .A(n3997), .B(n1532), .Z(n3773) );
  AN2P U4027 ( .A(n3953), .B(n3915), .Z(n3803) );
  AN2P U4028 ( .A(n914), .B(n3953), .Z(n3805) );
  AN2P U4029 ( .A(n3953), .B(n917), .Z(n3807) );
  AN2P U4030 ( .A(n3996), .B(n915), .Z(n3809) );
  AN2P U4031 ( .A(n1640), .B(n3952), .Z(n3820) );
  AN2P U4032 ( .A(n889), .B(n3953), .Z(n3828) );
  AN2P U4033 ( .A(n890), .B(n3996), .Z(n3830) );
  AN2P U4034 ( .A(n4734), .B(n3996), .Z(n3832) );
  AN2P U4035 ( .A(n1169), .B(n3996), .Z(n3841) );
  AN2P U4036 ( .A(n1170), .B(n3952), .Z(n3842) );
  AN2P U4037 ( .A(n3917), .B(n1168), .Z(n3843) );
  IVA U4038 ( .A(n3881), .Z(n3874) );
  IVA U4039 ( .A(n3881), .Z(n3875) );
  IVA U4040 ( .A(n3881), .Z(n3876) );
  IVA U4041 ( .A(n3885), .Z(n3877) );
  IVA U4042 ( .A(n3885), .Z(n3878) );
  IVA U4043 ( .A(LogIn2[46]), .Z(n3879) );
  IVA U4044 ( .A(LogIn2[46]), .Z(n3880) );
  IVA U4045 ( .A(n3878), .Z(n3881) );
  IVA U4046 ( .A(n3933), .Z(n3886) );
  IVA U4047 ( .A(n3933), .Z(n3887) );
  IVA U4048 ( .A(n3938), .Z(n3888) );
  IVA U4049 ( .A(n3913), .Z(n3889) );
  IVA U4050 ( .A(n3926), .Z(n3890) );
  IVA U4051 ( .A(n3938), .Z(n3891) );
  IVA U4052 ( .A(LogIn2[45]), .Z(n3892) );
  IVA U4053 ( .A(LogIn2[45]), .Z(n3893) );
  IVA U4054 ( .A(n3935), .Z(n3894) );
  IVA U4055 ( .A(n3934), .Z(n3895) );
  IVA U4056 ( .A(n3934), .Z(n3896) );
  IVA U4057 ( .A(n3934), .Z(n3897) );
  IVA U4058 ( .A(n3934), .Z(n3898) );
  IVA U4059 ( .A(n3934), .Z(n3899) );
  IVA U4060 ( .A(n3934), .Z(n3900) );
  IVA U4061 ( .A(n3935), .Z(n3901) );
  IVA U4062 ( .A(n3935), .Z(n3902) );
  IVA U4063 ( .A(n3935), .Z(n3903) );
  IVA U4064 ( .A(n3936), .Z(n3904) );
  IVA U4065 ( .A(n3936), .Z(n3905) );
  IVA U4066 ( .A(n3936), .Z(n3906) );
  IVA U4067 ( .A(n3937), .Z(n3907) );
  IVA U4068 ( .A(n3937), .Z(n3908) );
  IVA U4069 ( .A(n3937), .Z(n3909) );
  IVA U4070 ( .A(n3938), .Z(n3910) );
  IVA U4071 ( .A(n3938), .Z(n3911) );
  IVA U4072 ( .A(n3938), .Z(n3912) );
  IV U4073 ( .A(n3886), .Z(n3913) );
  IVA U4074 ( .A(n3932), .Z(n3933) );
  IVA U4075 ( .A(n3890), .Z(n3934) );
  IVA U4076 ( .A(n3890), .Z(n3935) );
  IVA U4077 ( .A(n3890), .Z(n3936) );
  IVA U4078 ( .A(n3894), .Z(n3937) );
  IVA U4079 ( .A(n3893), .Z(n3938) );
  IVA U4080 ( .A(n4003), .Z(n3972) );
  IVA U4081 ( .A(LogIn2[43]), .Z(n3973) );
  IVA U4082 ( .A(LogIn2[43]), .Z(n3974) );
  IVA U4083 ( .A(LogIn2[43]), .Z(n3975) );
  IVA U4084 ( .A(n4021), .Z(n3976) );
  IVA U4085 ( .A(n3993), .Z(n3977) );
  IVA U4086 ( .A(n4017), .Z(n3978) );
  IVA U4087 ( .A(n4017), .Z(n3979) );
  IVA U4088 ( .A(n4017), .Z(n3980) );
  IVA U4089 ( .A(n4018), .Z(n3981) );
  IVA U4090 ( .A(n4018), .Z(n3982) );
  IVA U4091 ( .A(n4018), .Z(n3983) );
  IVA U4092 ( .A(n4019), .Z(n3984) );
  IVA U4093 ( .A(n4019), .Z(n3985) );
  IVA U4094 ( .A(n4019), .Z(n3986) );
  IVA U4095 ( .A(n4020), .Z(n3987) );
  IVA U4096 ( .A(n4020), .Z(n3988) );
  IVA U4097 ( .A(n4020), .Z(n3989) );
  IVA U4098 ( .A(n4021), .Z(n3990) );
  IVA U4099 ( .A(n4021), .Z(n3991) );
  IVA U4100 ( .A(n4021), .Z(n3992) );
  IV U4101 ( .A(n3972), .Z(n3993) );
  IVA U4102 ( .A(n3972), .Z(n4017) );
  IVA U4103 ( .A(n3991), .Z(n4018) );
  IVA U4104 ( .A(n3990), .Z(n4019) );
  IVA U4105 ( .A(n3977), .Z(n4020) );
  IVA U4106 ( .A(n3972), .Z(n4021) );
  IVA U4107 ( .A(n4322), .Z(n4022) );
  IVA U4108 ( .A(n4322), .Z(n4023) );
  IVA U4109 ( .A(n4323), .Z(n4024) );
  IVA U4110 ( .A(n4323), .Z(n4025) );
  IVA U4111 ( .A(n4323), .Z(n4026) );
  IVA U4112 ( .A(n4324), .Z(n4027) );
  IVA U4113 ( .A(n4324), .Z(n4028) );
  IVA U4114 ( .A(n4324), .Z(n4029) );
  IVA U4115 ( .A(n4325), .Z(n4030) );
  IVA U4116 ( .A(n4325), .Z(n4031) );
  IVA U4117 ( .A(n4325), .Z(n4032) );
  IVA U4118 ( .A(n4326), .Z(n4033) );
  IVA U4119 ( .A(n4326), .Z(n4034) );
  IVA U4120 ( .A(n4326), .Z(n4035) );
  IVA U4121 ( .A(n4327), .Z(n4036) );
  IVA U4122 ( .A(n4327), .Z(n4037) );
  IVA U4123 ( .A(n4327), .Z(n4038) );
  IVA U4124 ( .A(n4328), .Z(n4039) );
  IVA U4125 ( .A(n4328), .Z(n4040) );
  IVA U4126 ( .A(n4328), .Z(n4041) );
  IVA U4127 ( .A(n4329), .Z(n4042) );
  IVA U4128 ( .A(n4329), .Z(n4043) );
  IVA U4129 ( .A(n4329), .Z(n4044) );
  IVA U4130 ( .A(n4330), .Z(n4045) );
  IVA U4131 ( .A(n4330), .Z(n4046) );
  IVA U4132 ( .A(n4330), .Z(n4047) );
  IVA U4133 ( .A(n4331), .Z(n4048) );
  IVA U4134 ( .A(n4331), .Z(n4049) );
  IVA U4135 ( .A(n4331), .Z(n4050) );
  IVA U4136 ( .A(n4332), .Z(n4051) );
  IVA U4137 ( .A(n4332), .Z(n4052) );
  IVA U4138 ( .A(n4332), .Z(n4053) );
  IVA U4139 ( .A(n4333), .Z(n4054) );
  IVA U4140 ( .A(n4333), .Z(n4055) );
  IVA U4141 ( .A(n4333), .Z(n4056) );
  IVA U4142 ( .A(n4334), .Z(n4057) );
  IVA U4143 ( .A(n4334), .Z(n4058) );
  IVA U4144 ( .A(n4334), .Z(n4059) );
  IVA U4145 ( .A(n4335), .Z(n4060) );
  IVA U4146 ( .A(n4335), .Z(n4061) );
  IVA U4147 ( .A(n4335), .Z(n4062) );
  IVA U4148 ( .A(n4336), .Z(n4063) );
  IVA U4149 ( .A(n4336), .Z(n4064) );
  IVA U4150 ( .A(n4336), .Z(n4065) );
  IVA U4151 ( .A(n4337), .Z(n4066) );
  IVA U4152 ( .A(n4337), .Z(n4067) );
  IVA U4153 ( .A(n4337), .Z(n4068) );
  IVA U4154 ( .A(n4338), .Z(n4069) );
  IVA U4155 ( .A(n4338), .Z(n4070) );
  IVA U4156 ( .A(n4338), .Z(n4071) );
  IVA U4157 ( .A(n4339), .Z(n4072) );
  IVA U4158 ( .A(n4339), .Z(n4073) );
  IVA U4159 ( .A(n4339), .Z(n4074) );
  IVA U4160 ( .A(n4340), .Z(n4075) );
  IVA U4161 ( .A(n4340), .Z(n4076) );
  IVA U4162 ( .A(n4340), .Z(n4077) );
  IVA U4163 ( .A(n4341), .Z(n4078) );
  IVA U4164 ( .A(n4341), .Z(n4079) );
  IVA U4165 ( .A(n4341), .Z(n4080) );
  IVA U4166 ( .A(n4342), .Z(n4081) );
  IVA U4167 ( .A(n4342), .Z(n4082) );
  IVA U4168 ( .A(n4342), .Z(n4083) );
  IVA U4169 ( .A(n4343), .Z(n4084) );
  IVA U4170 ( .A(n4343), .Z(n4085) );
  IVA U4171 ( .A(n4343), .Z(n4086) );
  IVA U4172 ( .A(n4344), .Z(n4087) );
  IVA U4173 ( .A(n4344), .Z(n4088) );
  IVA U4174 ( .A(n4344), .Z(n4089) );
  IVA U4175 ( .A(n4345), .Z(n4090) );
  IVA U4176 ( .A(n4345), .Z(n4091) );
  IVA U4177 ( .A(n4345), .Z(n4092) );
  IVA U4178 ( .A(n4346), .Z(n4093) );
  IVA U4179 ( .A(n4346), .Z(n4094) );
  IVA U4180 ( .A(n4346), .Z(n4095) );
  IVA U4181 ( .A(n4347), .Z(n4096) );
  IVA U4182 ( .A(n4347), .Z(n4097) );
  IVA U4183 ( .A(n4347), .Z(n4098) );
  IVA U4184 ( .A(n4348), .Z(n4099) );
  IVA U4185 ( .A(n4348), .Z(n4100) );
  IVA U4186 ( .A(n4348), .Z(n4101) );
  IVA U4187 ( .A(n4349), .Z(n4102) );
  IVA U4188 ( .A(n4349), .Z(n4103) );
  IVA U4189 ( .A(n4349), .Z(n4104) );
  IVA U4190 ( .A(n4350), .Z(n4105) );
  IVA U4191 ( .A(n4350), .Z(n4106) );
  IVA U4192 ( .A(n4350), .Z(n4107) );
  IVA U4193 ( .A(n4351), .Z(n4108) );
  IVA U4194 ( .A(n4351), .Z(n4109) );
  IVA U4195 ( .A(n4351), .Z(n4110) );
  IVA U4196 ( .A(n4352), .Z(n4111) );
  IVA U4197 ( .A(n4352), .Z(n4112) );
  IVA U4198 ( .A(n4352), .Z(n4113) );
  IVA U4199 ( .A(n4353), .Z(n4114) );
  IVA U4200 ( .A(n4353), .Z(n4115) );
  IVA U4201 ( .A(n4353), .Z(n4116) );
  IVA U4202 ( .A(n4354), .Z(n4117) );
  IVA U4203 ( .A(n4354), .Z(n4118) );
  IVA U4204 ( .A(n4354), .Z(n4119) );
  IVA U4205 ( .A(n4355), .Z(n4120) );
  IVA U4206 ( .A(n4355), .Z(n4121) );
  IVA U4207 ( .A(n4355), .Z(n4122) );
  IVA U4208 ( .A(n4356), .Z(n4123) );
  IVA U4209 ( .A(n4356), .Z(n4124) );
  IVA U4210 ( .A(n4356), .Z(n4125) );
  IVA U4211 ( .A(n4357), .Z(n4126) );
  IVA U4212 ( .A(n4357), .Z(n4127) );
  IVA U4213 ( .A(n4357), .Z(n4128) );
  IVA U4214 ( .A(n4358), .Z(n4129) );
  IVA U4215 ( .A(n4358), .Z(n4130) );
  IVA U4216 ( .A(n4358), .Z(n4131) );
  IVA U4217 ( .A(n4359), .Z(n4132) );
  IVA U4218 ( .A(n4359), .Z(n4133) );
  IVA U4219 ( .A(n4359), .Z(n4134) );
  IVA U4220 ( .A(n4360), .Z(n4135) );
  IVA U4221 ( .A(n4360), .Z(n4136) );
  IVA U4222 ( .A(n4360), .Z(n4137) );
  IVA U4223 ( .A(n4361), .Z(n4138) );
  IVA U4224 ( .A(n4361), .Z(n4139) );
  IVA U4225 ( .A(n4361), .Z(n4140) );
  IVA U4226 ( .A(n4362), .Z(n4141) );
  IVA U4227 ( .A(n4362), .Z(n4142) );
  IVA U4228 ( .A(n4362), .Z(n4143) );
  IVA U4229 ( .A(n4363), .Z(n4144) );
  IVA U4230 ( .A(n4363), .Z(n4145) );
  IVA U4231 ( .A(n4363), .Z(n4146) );
  IVA U4232 ( .A(n4364), .Z(n4147) );
  IVA U4233 ( .A(n4364), .Z(n4148) );
  IVA U4234 ( .A(n4364), .Z(n4149) );
  IVA U4235 ( .A(n4365), .Z(n4150) );
  IVA U4236 ( .A(n4365), .Z(n4151) );
  IVA U4237 ( .A(n4365), .Z(n4152) );
  IVA U4238 ( .A(n4366), .Z(n4153) );
  IVA U4239 ( .A(n4366), .Z(n4154) );
  IVA U4240 ( .A(n4366), .Z(n4155) );
  IVA U4241 ( .A(n4367), .Z(n4156) );
  IVA U4242 ( .A(n4367), .Z(n4157) );
  IVA U4243 ( .A(n4367), .Z(n4158) );
  IVA U4244 ( .A(n4368), .Z(n4159) );
  IVA U4245 ( .A(n4368), .Z(n4160) );
  IVA U4246 ( .A(n4368), .Z(n4161) );
  IVA U4247 ( .A(n4369), .Z(n4162) );
  IVA U4248 ( .A(n4369), .Z(n4163) );
  IVA U4249 ( .A(n4369), .Z(n4164) );
  IVA U4250 ( .A(n4370), .Z(n4165) );
  IVA U4251 ( .A(n4370), .Z(n4166) );
  IVA U4252 ( .A(n4370), .Z(n4167) );
  IVA U4253 ( .A(n4371), .Z(n4168) );
  IVA U4254 ( .A(n4371), .Z(n4169) );
  IVA U4255 ( .A(n4371), .Z(n4170) );
  IVA U4256 ( .A(n4372), .Z(n4171) );
  IVA U4257 ( .A(n4372), .Z(n4172) );
  IVA U4258 ( .A(n4372), .Z(n4173) );
  IVA U4259 ( .A(n4373), .Z(n4174) );
  IVA U4260 ( .A(n4373), .Z(n4175) );
  IVA U4261 ( .A(n4373), .Z(n4176) );
  IVA U4262 ( .A(n4374), .Z(n4177) );
  IVA U4263 ( .A(n4374), .Z(n4178) );
  IVA U4264 ( .A(n4374), .Z(n4179) );
  IVA U4265 ( .A(n4375), .Z(n4180) );
  IVA U4266 ( .A(n4375), .Z(n4181) );
  IVA U4267 ( .A(n4375), .Z(n4182) );
  IVA U4268 ( .A(n4376), .Z(n4183) );
  IVA U4269 ( .A(n4376), .Z(n4184) );
  IVA U4270 ( .A(n4376), .Z(n4185) );
  IVA U4271 ( .A(n4377), .Z(n4186) );
  IVA U4272 ( .A(n4377), .Z(n4187) );
  IVA U4273 ( .A(n4377), .Z(n4188) );
  IVA U4274 ( .A(n4378), .Z(n4189) );
  IVA U4275 ( .A(n4378), .Z(n4190) );
  IVA U4276 ( .A(n4378), .Z(n4191) );
  IVA U4277 ( .A(n4379), .Z(n4192) );
  IVA U4278 ( .A(n4379), .Z(n4193) );
  IVA U4279 ( .A(n4379), .Z(n4194) );
  IVA U4280 ( .A(n4380), .Z(n4195) );
  IVA U4281 ( .A(n4380), .Z(n4196) );
  IVA U4282 ( .A(n4380), .Z(n4197) );
  IVA U4283 ( .A(n4381), .Z(n4198) );
  IVA U4284 ( .A(n4381), .Z(n4199) );
  IVA U4285 ( .A(n4381), .Z(n4200) );
  IVA U4286 ( .A(n4382), .Z(n4201) );
  IVA U4287 ( .A(n4382), .Z(n4202) );
  IVA U4288 ( .A(n4382), .Z(n4203) );
  IVA U4289 ( .A(n4383), .Z(n4204) );
  IVA U4290 ( .A(n4383), .Z(n4205) );
  IVA U4291 ( .A(n4383), .Z(n4206) );
  IV U4292 ( .A(n4030), .Z(n4207) );
  IVA U4293 ( .A(n4329), .Z(n4301) );
  IVA U4294 ( .A(n4330), .Z(n4302) );
  IVA U4295 ( .A(n4328), .Z(n4303) );
  IVA U4296 ( .A(n4359), .Z(n4304) );
  IVA U4297 ( .A(LogIn2[42]), .Z(n4305) );
  IVA U4298 ( .A(LogIn2[42]), .Z(n4306) );
  IVA U4299 ( .A(LogIn2[42]), .Z(n4307) );
  IVA U4300 ( .A(LogIn2[42]), .Z(n4308) );
  IVA U4301 ( .A(LogIn2[42]), .Z(n4309) );
  IVA U4302 ( .A(LogIn2[42]), .Z(n4310) );
  IVA U4303 ( .A(n4372), .Z(n4311) );
  IVA U4304 ( .A(n4382), .Z(n4312) );
  IVA U4305 ( .A(n4330), .Z(n4313) );
  IVA U4306 ( .A(n4336), .Z(n4314) );
  IVA U4307 ( .A(n4364), .Z(n4315) );
  IVA U4308 ( .A(LogIn2[42]), .Z(n4316) );
  IVA U4309 ( .A(n4329), .Z(n4317) );
  IVA U4310 ( .A(LogIn2[42]), .Z(n4318) );
  IVA U4311 ( .A(n4357), .Z(n4319) );
  IVA U4312 ( .A(LogIn2[42]), .Z(n4320) );
  IVA U4313 ( .A(LogIn2[42]), .Z(n4321) );
  IVA U4314 ( .A(n4321), .Z(n4322) );
  IVA U4315 ( .A(n4321), .Z(n4323) );
  IVA U4316 ( .A(n4321), .Z(n4324) );
  IVA U4317 ( .A(n4320), .Z(n4325) );
  IVA U4318 ( .A(n4320), .Z(n4326) );
  IVA U4319 ( .A(n4320), .Z(n4327) );
  IVA U4320 ( .A(n4319), .Z(n4328) );
  IVA U4321 ( .A(n4319), .Z(n4329) );
  IVA U4322 ( .A(n4319), .Z(n4330) );
  IVA U4323 ( .A(n4318), .Z(n4331) );
  IVA U4324 ( .A(n4318), .Z(n4332) );
  IVA U4325 ( .A(n4318), .Z(n4333) );
  IVA U4326 ( .A(n4317), .Z(n4334) );
  IVA U4327 ( .A(n4317), .Z(n4335) );
  IVA U4328 ( .A(n4317), .Z(n4336) );
  IVA U4329 ( .A(n4316), .Z(n4337) );
  IVA U4330 ( .A(n4316), .Z(n4338) );
  IVA U4331 ( .A(n4316), .Z(n4339) );
  IVA U4332 ( .A(n4315), .Z(n4340) );
  IVA U4333 ( .A(n4315), .Z(n4341) );
  IVA U4334 ( .A(n4315), .Z(n4342) );
  IVA U4335 ( .A(n4314), .Z(n4343) );
  IVA U4336 ( .A(n4314), .Z(n4344) );
  IVA U4337 ( .A(n4314), .Z(n4345) );
  IVA U4338 ( .A(n4313), .Z(n4346) );
  IVA U4339 ( .A(n4313), .Z(n4347) );
  IVA U4340 ( .A(n4313), .Z(n4348) );
  IVA U4341 ( .A(n4312), .Z(n4349) );
  IVA U4342 ( .A(n4312), .Z(n4350) );
  IVA U4343 ( .A(n4312), .Z(n4351) );
  IVA U4344 ( .A(n4311), .Z(n4352) );
  IVA U4345 ( .A(n4311), .Z(n4353) );
  IVA U4346 ( .A(n4311), .Z(n4354) );
  IVA U4347 ( .A(n4310), .Z(n4355) );
  IVA U4348 ( .A(n4310), .Z(n4356) );
  IVA U4349 ( .A(n4310), .Z(n4357) );
  IVA U4350 ( .A(n4309), .Z(n4358) );
  IVA U4351 ( .A(n4309), .Z(n4359) );
  IVA U4352 ( .A(n4309), .Z(n4360) );
  IVA U4353 ( .A(n4308), .Z(n4361) );
  IVA U4354 ( .A(n4308), .Z(n4362) );
  IVA U4355 ( .A(n4308), .Z(n4363) );
  IVA U4356 ( .A(n4307), .Z(n4364) );
  IVA U4357 ( .A(n4307), .Z(n4365) );
  IVA U4358 ( .A(n4307), .Z(n4366) );
  IVA U4359 ( .A(n4306), .Z(n4367) );
  IVA U4360 ( .A(n4306), .Z(n4368) );
  IVA U4361 ( .A(n4306), .Z(n4369) );
  IVA U4362 ( .A(n4305), .Z(n4370) );
  IVA U4363 ( .A(n4305), .Z(n4371) );
  IVA U4364 ( .A(n4305), .Z(n4372) );
  IVA U4365 ( .A(n4304), .Z(n4373) );
  IVA U4366 ( .A(n4304), .Z(n4374) );
  IVA U4367 ( .A(n4304), .Z(n4375) );
  IVA U4368 ( .A(n4303), .Z(n4376) );
  IVA U4369 ( .A(n4303), .Z(n4377) );
  IVA U4370 ( .A(n4303), .Z(n4378) );
  IVA U4371 ( .A(n4302), .Z(n4379) );
  IVA U4372 ( .A(n4302), .Z(n4380) );
  IVA U4373 ( .A(n4302), .Z(n4381) );
  IVA U4374 ( .A(n4301), .Z(n4382) );
  IVA U4375 ( .A(n4301), .Z(n4383) );
  IVA U4376 ( .A(n4662), .Z(n4384) );
  IVA U4377 ( .A(n4662), .Z(n4385) );
  IVA U4378 ( .A(n4663), .Z(n4386) );
  IVA U4379 ( .A(n4663), .Z(n4387) );
  IVA U4380 ( .A(n4663), .Z(n4388) );
  IVA U4381 ( .A(n4664), .Z(n4389) );
  IVA U4382 ( .A(n4664), .Z(n4390) );
  IVA U4383 ( .A(n4664), .Z(n4391) );
  IVA U4384 ( .A(n4665), .Z(n4392) );
  IVA U4385 ( .A(n4665), .Z(n4393) );
  IVA U4386 ( .A(n4665), .Z(n4394) );
  IVA U4387 ( .A(n4666), .Z(n4395) );
  IVA U4388 ( .A(n4666), .Z(n4396) );
  IVA U4389 ( .A(n4666), .Z(n4397) );
  IVA U4390 ( .A(n4667), .Z(n4398) );
  IVA U4391 ( .A(n4667), .Z(n4399) );
  IVA U4392 ( .A(n4667), .Z(n4400) );
  IVA U4393 ( .A(n4668), .Z(n4401) );
  IVA U4394 ( .A(n4668), .Z(n4402) );
  IVA U4395 ( .A(n4668), .Z(n4403) );
  IVA U4396 ( .A(n4669), .Z(n4404) );
  IVA U4397 ( .A(n4669), .Z(n4405) );
  IVA U4398 ( .A(n4669), .Z(n4406) );
  IVA U4399 ( .A(n4670), .Z(n4407) );
  IVA U4400 ( .A(n4670), .Z(n4408) );
  IVA U4401 ( .A(n4670), .Z(n4409) );
  IVA U4402 ( .A(n4671), .Z(n4410) );
  IVA U4403 ( .A(n4671), .Z(n4411) );
  IVA U4404 ( .A(n4671), .Z(n4412) );
  IVA U4405 ( .A(n4672), .Z(n4413) );
  IVA U4406 ( .A(n4672), .Z(n4414) );
  IVA U4407 ( .A(n4672), .Z(n4415) );
  IVA U4408 ( .A(n4673), .Z(n4416) );
  IVA U4409 ( .A(n4673), .Z(n4417) );
  IVA U4410 ( .A(n4673), .Z(n4418) );
  IVA U4411 ( .A(n4674), .Z(n4419) );
  IVA U4412 ( .A(n4674), .Z(n4420) );
  IVA U4413 ( .A(n4674), .Z(n4421) );
  IVA U4414 ( .A(n4675), .Z(n4422) );
  IVA U4415 ( .A(n4675), .Z(n4423) );
  IVA U4416 ( .A(n4675), .Z(n4424) );
  IVA U4417 ( .A(n4676), .Z(n4425) );
  IVA U4418 ( .A(n4676), .Z(n4426) );
  IVA U4419 ( .A(n4676), .Z(n4427) );
  IVA U4420 ( .A(n4677), .Z(n4428) );
  IVA U4421 ( .A(n4677), .Z(n4429) );
  IVA U4422 ( .A(n4677), .Z(n4430) );
  IVA U4423 ( .A(n4678), .Z(n4431) );
  IVA U4424 ( .A(n4678), .Z(n4432) );
  IVA U4425 ( .A(n4678), .Z(n4433) );
  IVA U4426 ( .A(n4679), .Z(n4434) );
  IVA U4427 ( .A(n4679), .Z(n4435) );
  IVA U4428 ( .A(n4679), .Z(n4436) );
  IVA U4429 ( .A(n4680), .Z(n4437) );
  IVA U4430 ( .A(n4680), .Z(n4438) );
  IVA U4431 ( .A(n4680), .Z(n4439) );
  IVA U4432 ( .A(n4681), .Z(n4440) );
  IVA U4433 ( .A(n4681), .Z(n4441) );
  IVA U4434 ( .A(n4681), .Z(n4442) );
  IVA U4435 ( .A(n4682), .Z(n4443) );
  IVA U4436 ( .A(n4682), .Z(n4444) );
  IVA U4437 ( .A(n4682), .Z(n4445) );
  IVA U4438 ( .A(n4683), .Z(n4446) );
  IVA U4439 ( .A(n4683), .Z(n4447) );
  IVA U4440 ( .A(n4683), .Z(n4448) );
  IVA U4441 ( .A(n4684), .Z(n4449) );
  IVA U4442 ( .A(n4684), .Z(n4450) );
  IVA U4443 ( .A(n4684), .Z(n4451) );
  IVA U4444 ( .A(n4685), .Z(n4452) );
  IVA U4445 ( .A(n4685), .Z(n4453) );
  IVA U4446 ( .A(n4685), .Z(n4454) );
  IVA U4447 ( .A(n4686), .Z(n4455) );
  IVA U4448 ( .A(n4686), .Z(n4456) );
  IVA U4449 ( .A(n4686), .Z(n4457) );
  IVA U4450 ( .A(n4687), .Z(n4458) );
  IVA U4451 ( .A(n4687), .Z(n4459) );
  IVA U4452 ( .A(n4687), .Z(n4460) );
  IVA U4453 ( .A(n4688), .Z(n4461) );
  IVA U4454 ( .A(n4688), .Z(n4462) );
  IVA U4455 ( .A(n4688), .Z(n4463) );
  IVA U4456 ( .A(n4689), .Z(n4464) );
  IVA U4457 ( .A(n4689), .Z(n4465) );
  IVA U4458 ( .A(n4689), .Z(n4466) );
  IVA U4459 ( .A(n4690), .Z(n4467) );
  IVA U4460 ( .A(n4690), .Z(n4468) );
  IVA U4461 ( .A(n4690), .Z(n4469) );
  IVA U4462 ( .A(n4691), .Z(n4470) );
  IVA U4463 ( .A(n4691), .Z(n4471) );
  IVA U4464 ( .A(n4691), .Z(n4472) );
  IVA U4465 ( .A(n4692), .Z(n4473) );
  IVA U4466 ( .A(n4692), .Z(n4474) );
  IVA U4467 ( .A(n4692), .Z(n4475) );
  IVA U4468 ( .A(n4693), .Z(n4476) );
  IVA U4469 ( .A(n4693), .Z(n4477) );
  IVA U4470 ( .A(n4693), .Z(n4478) );
  IVA U4471 ( .A(n4694), .Z(n4479) );
  IVA U4472 ( .A(n4694), .Z(n4480) );
  IVA U4473 ( .A(n4694), .Z(n4481) );
  IVA U4474 ( .A(n4695), .Z(n4482) );
  IVA U4475 ( .A(n4695), .Z(n4483) );
  IVA U4476 ( .A(n4695), .Z(n4484) );
  IVA U4477 ( .A(n4696), .Z(n4485) );
  IVA U4478 ( .A(n4696), .Z(n4486) );
  IVA U4479 ( .A(n4696), .Z(n4487) );
  IVA U4480 ( .A(n4697), .Z(n4488) );
  IVA U4481 ( .A(n4697), .Z(n4489) );
  IVA U4482 ( .A(n4697), .Z(n4490) );
  IVA U4483 ( .A(n4698), .Z(n4491) );
  IVA U4484 ( .A(n4698), .Z(n4492) );
  IVA U4485 ( .A(n4698), .Z(n4493) );
  IVA U4486 ( .A(n4699), .Z(n4494) );
  IVA U4487 ( .A(n4699), .Z(n4495) );
  IVA U4488 ( .A(n4699), .Z(n4496) );
  IVA U4489 ( .A(n4700), .Z(n4497) );
  IVA U4490 ( .A(n4700), .Z(n4498) );
  IVA U4491 ( .A(n4700), .Z(n4499) );
  IVA U4492 ( .A(n4701), .Z(n4500) );
  IVA U4493 ( .A(n4701), .Z(n4501) );
  IVA U4494 ( .A(n4701), .Z(n4502) );
  IVA U4495 ( .A(n4702), .Z(n4503) );
  IVA U4496 ( .A(n4702), .Z(n4504) );
  IVA U4497 ( .A(n4702), .Z(n4505) );
  IVA U4498 ( .A(n4703), .Z(n4506) );
  IVA U4499 ( .A(n4703), .Z(n4507) );
  IVA U4500 ( .A(n4703), .Z(n4508) );
  IVA U4501 ( .A(n4704), .Z(n4509) );
  IVA U4502 ( .A(n4704), .Z(n4510) );
  IVA U4503 ( .A(n4704), .Z(n4511) );
  IVA U4504 ( .A(n4705), .Z(n4512) );
  IVA U4505 ( .A(n4705), .Z(n4513) );
  IVA U4506 ( .A(n4705), .Z(n4514) );
  IVA U4507 ( .A(n4706), .Z(n4515) );
  IVA U4508 ( .A(n4706), .Z(n4516) );
  IVA U4509 ( .A(n4706), .Z(n4517) );
  IVA U4510 ( .A(n4707), .Z(n4518) );
  IVA U4511 ( .A(n4707), .Z(n4519) );
  IVA U4512 ( .A(n4707), .Z(n4520) );
  IVA U4513 ( .A(n4708), .Z(n4521) );
  IVA U4514 ( .A(n4708), .Z(n4522) );
  IVA U4515 ( .A(n4708), .Z(n4523) );
  IVA U4516 ( .A(n4709), .Z(n4524) );
  IVA U4517 ( .A(n4709), .Z(n4525) );
  IVA U4518 ( .A(n4709), .Z(n4526) );
  IVA U4519 ( .A(n4710), .Z(n4527) );
  IVA U4520 ( .A(n4710), .Z(n4528) );
  IVA U4521 ( .A(n4710), .Z(n4529) );
  IVA U4522 ( .A(n4711), .Z(n4530) );
  IVA U4523 ( .A(n4711), .Z(n4531) );
  IVA U4524 ( .A(n4711), .Z(n4532) );
  IVA U4525 ( .A(n4712), .Z(n4533) );
  IVA U4526 ( .A(n4712), .Z(n4534) );
  IVA U4527 ( .A(n4712), .Z(n4535) );
  IVA U4528 ( .A(n4713), .Z(n4536) );
  IVA U4529 ( .A(n4713), .Z(n4537) );
  IVA U4530 ( .A(n4713), .Z(n4538) );
  IVA U4531 ( .A(n4714), .Z(n4539) );
  IVA U4532 ( .A(n4714), .Z(n4540) );
  IVA U4533 ( .A(n4714), .Z(n4541) );
  IVA U4534 ( .A(n4715), .Z(n4542) );
  IVA U4535 ( .A(n4715), .Z(n4543) );
  IVA U4536 ( .A(n4715), .Z(n4544) );
  IVA U4537 ( .A(n4716), .Z(n4545) );
  IVA U4538 ( .A(n4716), .Z(n4546) );
  IVA U4539 ( .A(n4716), .Z(n4547) );
  IVA U4540 ( .A(n4717), .Z(n4548) );
  IVA U4541 ( .A(n4717), .Z(n4549) );
  IVA U4542 ( .A(n4717), .Z(n4550) );
  IVA U4543 ( .A(n4718), .Z(n4551) );
  IVA U4544 ( .A(n4718), .Z(n4552) );
  IVA U4545 ( .A(n4718), .Z(n4553) );
  IVA U4546 ( .A(n4719), .Z(n4554) );
  IVA U4547 ( .A(n4719), .Z(n4555) );
  IVA U4548 ( .A(n4719), .Z(n4556) );
  IVA U4549 ( .A(n4720), .Z(n4557) );
  IVA U4550 ( .A(n4720), .Z(n4558) );
  IVA U4551 ( .A(n4720), .Z(n4559) );
  IVA U4552 ( .A(n4706), .Z(n4642) );
  IVA U4553 ( .A(LogIn2[41]), .Z(n4643) );
  IVA U4554 ( .A(n4669), .Z(n4644) );
  IVA U4555 ( .A(n4667), .Z(n4645) );
  IVA U4556 ( .A(LogIn2[41]), .Z(n4646) );
  IVA U4557 ( .A(LogIn2[41]), .Z(n4647) );
  IVA U4558 ( .A(n4667), .Z(n4648) );
  IVA U4559 ( .A(n4667), .Z(n4649) );
  IVA U4560 ( .A(n4708), .Z(n4650) );
  IVA U4561 ( .A(n4662), .Z(n4651) );
  IVA U4562 ( .A(LogIn2[41]), .Z(n4652) );
  IVA U4563 ( .A(n4712), .Z(n4653) );
  IVA U4564 ( .A(LogIn2[41]), .Z(n4654) );
  IVA U4565 ( .A(LogIn2[41]), .Z(n4655) );
  IVA U4566 ( .A(n4675), .Z(n4656) );
  IVA U4567 ( .A(LogIn2[41]), .Z(n4657) );
  IVA U4568 ( .A(n4720), .Z(n4658) );
  IVA U4569 ( .A(LogIn2[41]), .Z(n4659) );
  IVA U4570 ( .A(LogIn2[41]), .Z(n4660) );
  IVA U4571 ( .A(LogIn2[41]), .Z(n4661) );
  IVA U4572 ( .A(n4661), .Z(n4662) );
  IVA U4573 ( .A(n4661), .Z(n4663) );
  IVA U4574 ( .A(n4661), .Z(n4664) );
  IVA U4575 ( .A(n4660), .Z(n4665) );
  IVA U4576 ( .A(n4660), .Z(n4666) );
  IVA U4577 ( .A(n4660), .Z(n4667) );
  IVA U4578 ( .A(n4659), .Z(n4668) );
  IVA U4579 ( .A(n4659), .Z(n4669) );
  IVA U4580 ( .A(n4659), .Z(n4670) );
  IVA U4581 ( .A(n4658), .Z(n4671) );
  IVA U4582 ( .A(n4658), .Z(n4672) );
  IVA U4583 ( .A(n4658), .Z(n4673) );
  IVA U4584 ( .A(n4657), .Z(n4674) );
  IVA U4585 ( .A(n4657), .Z(n4675) );
  IVA U4586 ( .A(n4657), .Z(n4676) );
  IVA U4587 ( .A(n4656), .Z(n4677) );
  IVA U4588 ( .A(n4656), .Z(n4678) );
  IVA U4589 ( .A(n4656), .Z(n4679) );
  IVA U4590 ( .A(n4655), .Z(n4680) );
  IVA U4591 ( .A(n4655), .Z(n4681) );
  IVA U4592 ( .A(n4655), .Z(n4682) );
  IVA U4593 ( .A(n4654), .Z(n4683) );
  IVA U4594 ( .A(n4654), .Z(n4684) );
  IVA U4595 ( .A(n4654), .Z(n4685) );
  IVA U4596 ( .A(n4653), .Z(n4686) );
  IVA U4597 ( .A(n4653), .Z(n4687) );
  IVA U4598 ( .A(n4653), .Z(n4688) );
  IVA U4599 ( .A(n4652), .Z(n4689) );
  IVA U4600 ( .A(n4652), .Z(n4690) );
  IVA U4601 ( .A(n4652), .Z(n4691) );
  IVA U4602 ( .A(n4651), .Z(n4692) );
  IVA U4603 ( .A(n4651), .Z(n4693) );
  IVA U4604 ( .A(n4651), .Z(n4694) );
  IVA U4605 ( .A(n4650), .Z(n4695) );
  IVA U4606 ( .A(n4650), .Z(n4696) );
  IVA U4607 ( .A(n4650), .Z(n4697) );
  IVA U4608 ( .A(n4649), .Z(n4698) );
  IVA U4609 ( .A(n4649), .Z(n4699) );
  IVA U4610 ( .A(n4649), .Z(n4700) );
  IVA U4611 ( .A(n4648), .Z(n4701) );
  IVA U4612 ( .A(n4648), .Z(n4702) );
  IVA U4613 ( .A(n4648), .Z(n4703) );
  IVA U4614 ( .A(n4647), .Z(n4704) );
  IVA U4615 ( .A(n4647), .Z(n4705) );
  IVA U4616 ( .A(n4647), .Z(n4706) );
  IVA U4617 ( .A(n4646), .Z(n4707) );
  IVA U4618 ( .A(n4646), .Z(n4708) );
  IVA U4619 ( .A(n4646), .Z(n4709) );
  IVA U4620 ( .A(n4645), .Z(n4710) );
  IVA U4621 ( .A(n4645), .Z(n4711) );
  IVA U4622 ( .A(n4645), .Z(n4712) );
  IVA U4623 ( .A(n4644), .Z(n4713) );
  IVA U4624 ( .A(n4644), .Z(n4714) );
  IVA U4625 ( .A(n4644), .Z(n4715) );
  IVA U4626 ( .A(n4643), .Z(n4716) );
  IVA U4627 ( .A(n4643), .Z(n4717) );
  IVA U4628 ( .A(n4643), .Z(n4718) );
  IVA U4629 ( .A(n4642), .Z(n4719) );
  IVA U4630 ( .A(n4642), .Z(n4720) );
  IVA U4631 ( .A(n4970), .Z(n4721) );
  IVA U4632 ( .A(n4971), .Z(n4722) );
  IVA U4633 ( .A(n4971), .Z(n4723) );
  IVA U4634 ( .A(n4971), .Z(n4724) );
  IVA U4635 ( .A(n4972), .Z(n4725) );
  IVA U4636 ( .A(n4972), .Z(n4726) );
  IVA U4637 ( .A(n4972), .Z(n4727) );
  IVA U4638 ( .A(n4973), .Z(n4728) );
  IVA U4639 ( .A(n4973), .Z(n4729) );
  IVA U4640 ( .A(n4973), .Z(n4730) );
  IVA U4641 ( .A(n4974), .Z(n4731) );
  IVA U4642 ( .A(n4974), .Z(n4732) );
  IVA U4643 ( .A(n4974), .Z(n4733) );
  IVA U4644 ( .A(n4975), .Z(n4734) );
  IVA U4645 ( .A(n4975), .Z(n4735) );
  IVA U4646 ( .A(n4975), .Z(n4736) );
  IVA U4647 ( .A(n4976), .Z(n4737) );
  IVA U4648 ( .A(n4976), .Z(n4738) );
  IVA U4649 ( .A(n4976), .Z(n4739) );
  IVA U4650 ( .A(n4977), .Z(n4740) );
  IVA U4651 ( .A(n4977), .Z(n4741) );
  IVA U4652 ( .A(n4977), .Z(n4742) );
  IVA U4653 ( .A(n4978), .Z(n4743) );
  IVA U4654 ( .A(n4978), .Z(n4744) );
  IVA U4655 ( .A(n4978), .Z(n4745) );
  IVA U4656 ( .A(n4979), .Z(n4746) );
  IVA U4657 ( .A(n4979), .Z(n4747) );
  IVA U4658 ( .A(n4979), .Z(n4748) );
  IVA U4659 ( .A(n4980), .Z(n4749) );
  IVA U4660 ( .A(n4980), .Z(n4750) );
  IVA U4661 ( .A(n4980), .Z(n4751) );
  IVA U4662 ( .A(n4981), .Z(n4752) );
  IVA U4663 ( .A(n4981), .Z(n4753) );
  IVA U4664 ( .A(n4981), .Z(n4754) );
  IVA U4665 ( .A(n4982), .Z(n4755) );
  IVA U4666 ( .A(n4982), .Z(n4756) );
  IVA U4667 ( .A(n4982), .Z(n4757) );
  IVA U4668 ( .A(n4983), .Z(n4758) );
  IVA U4669 ( .A(n4983), .Z(n4759) );
  IVA U4670 ( .A(n4983), .Z(n4760) );
  IVA U4671 ( .A(n4984), .Z(n4761) );
  IVA U4672 ( .A(n4984), .Z(n4762) );
  IVA U4673 ( .A(n4984), .Z(n4763) );
  IVA U4674 ( .A(n4985), .Z(n4764) );
  IVA U4675 ( .A(n4985), .Z(n4765) );
  IVA U4676 ( .A(n4985), .Z(n4766) );
  IVA U4677 ( .A(n4986), .Z(n4767) );
  IVA U4678 ( .A(n4986), .Z(n4768) );
  IVA U4679 ( .A(n4986), .Z(n4769) );
  IVA U4680 ( .A(n4987), .Z(n4770) );
  IVA U4681 ( .A(n4987), .Z(n4771) );
  IVA U4682 ( .A(n4987), .Z(n4772) );
  IVA U4683 ( .A(n4988), .Z(n4773) );
  IVA U4684 ( .A(n4988), .Z(n4774) );
  IVA U4685 ( .A(n4988), .Z(n4775) );
  IVA U4686 ( .A(n4989), .Z(n4776) );
  IVA U4687 ( .A(n4989), .Z(n4777) );
  IVA U4688 ( .A(n4989), .Z(n4778) );
  IVA U4689 ( .A(n4990), .Z(n4779) );
  IVA U4690 ( .A(n4990), .Z(n4780) );
  IVA U4691 ( .A(n4990), .Z(n4781) );
  IVA U4692 ( .A(n4991), .Z(n4782) );
  IVA U4693 ( .A(n4991), .Z(n4783) );
  IVA U4694 ( .A(n4991), .Z(n4784) );
  IVA U4695 ( .A(n4992), .Z(n4785) );
  IVA U4696 ( .A(n4992), .Z(n4786) );
  IVA U4697 ( .A(n4992), .Z(n4787) );
  IVA U4698 ( .A(n4993), .Z(n4788) );
  IVA U4699 ( .A(n4993), .Z(n4789) );
  IVA U4700 ( .A(n4993), .Z(n4790) );
  IVA U4701 ( .A(n4994), .Z(n4791) );
  IVA U4702 ( .A(n4994), .Z(n4792) );
  IVA U4703 ( .A(n4994), .Z(n4793) );
  IVA U4704 ( .A(n4995), .Z(n4794) );
  IVA U4705 ( .A(n4995), .Z(n4795) );
  IVA U4706 ( .A(n4995), .Z(n4796) );
  IVA U4707 ( .A(n4996), .Z(n4797) );
  IVA U4708 ( .A(n4996), .Z(n4798) );
  IVA U4709 ( .A(n4996), .Z(n4799) );
  IVA U4710 ( .A(n4997), .Z(n4800) );
  IVA U4711 ( .A(n4997), .Z(n4801) );
  IVA U4712 ( .A(n4997), .Z(n4802) );
  IVA U4713 ( .A(n4998), .Z(n4803) );
  IVA U4714 ( .A(n4998), .Z(n4804) );
  IVA U4715 ( .A(n4998), .Z(n4805) );
  IVA U4716 ( .A(n4999), .Z(n4806) );
  IVA U4717 ( .A(n4999), .Z(n4807) );
  IVA U4718 ( .A(n4999), .Z(n4808) );
  IVA U4719 ( .A(n5000), .Z(n4809) );
  IVA U4720 ( .A(n5000), .Z(n4810) );
  IVA U4721 ( .A(n5000), .Z(n4811) );
  IVA U4722 ( .A(n5001), .Z(n4812) );
  IVA U4723 ( .A(n5001), .Z(n4813) );
  IVA U4724 ( .A(n5001), .Z(n4814) );
  IVA U4725 ( .A(n5002), .Z(n4815) );
  IVA U4726 ( .A(n5002), .Z(n4816) );
  IVA U4727 ( .A(n5002), .Z(n4817) );
  IVA U4728 ( .A(n5003), .Z(n4818) );
  IVA U4729 ( .A(n5003), .Z(n4819) );
  IVA U4730 ( .A(n5003), .Z(n4820) );
  IVA U4731 ( .A(n5004), .Z(n4821) );
  IVA U4732 ( .A(n5004), .Z(n4822) );
  IVA U4733 ( .A(n5004), .Z(n4823) );
  IVA U4734 ( .A(n5005), .Z(n4824) );
  IVA U4735 ( .A(n5005), .Z(n4825) );
  IVA U4736 ( .A(n5005), .Z(n4826) );
  IVA U4737 ( .A(n5006), .Z(n4827) );
  IVA U4738 ( .A(n5006), .Z(n4828) );
  IVA U4739 ( .A(n5006), .Z(n4829) );
  IVA U4740 ( .A(n5007), .Z(n4830) );
  IVA U4741 ( .A(n5007), .Z(n4831) );
  IVA U4742 ( .A(n5007), .Z(n4832) );
  IVA U4743 ( .A(n5008), .Z(n4833) );
  IVA U4744 ( .A(n5008), .Z(n4834) );
  IVA U4745 ( .A(n5008), .Z(n4835) );
  IVA U4746 ( .A(n5009), .Z(n4836) );
  IVA U4747 ( .A(n5009), .Z(n4837) );
  IVA U4748 ( .A(n5009), .Z(n4838) );
  IVA U4749 ( .A(n5010), .Z(n4839) );
  IVA U4750 ( .A(n5010), .Z(n4840) );
  IVA U4751 ( .A(n5010), .Z(n4841) );
  IVA U4752 ( .A(n5011), .Z(n4842) );
  IVA U4753 ( .A(n5011), .Z(n4843) );
  IVA U4754 ( .A(n5011), .Z(n4844) );
  IVA U4755 ( .A(n5012), .Z(n4845) );
  IVA U4756 ( .A(n5012), .Z(n4846) );
  IVA U4757 ( .A(n5012), .Z(n4847) );
  IVA U4758 ( .A(n5013), .Z(n4848) );
  IVA U4759 ( .A(n5013), .Z(n4849) );
  IVA U4760 ( .A(n5013), .Z(n4850) );
  IVA U4761 ( .A(n5014), .Z(n4851) );
  IVA U4762 ( .A(n5014), .Z(n4852) );
  IVA U4763 ( .A(n5014), .Z(n4853) );
  IVA U4764 ( .A(n5015), .Z(n4854) );
  IVA U4765 ( .A(n5015), .Z(n4855) );
  IVA U4766 ( .A(n5015), .Z(n4856) );
  IVA U4767 ( .A(n5016), .Z(n4857) );
  IVA U4768 ( .A(n5016), .Z(n4858) );
  IVA U4769 ( .A(n5016), .Z(n4859) );
  IVA U4770 ( .A(n5017), .Z(n4860) );
  IVA U4771 ( .A(n5017), .Z(n4861) );
  IVA U4772 ( .A(n5017), .Z(n4862) );
  IVA U4773 ( .A(n5018), .Z(n4863) );
  IVA U4774 ( .A(n5018), .Z(n4864) );
  IVA U4775 ( .A(n5018), .Z(n4865) );
  IVA U4776 ( .A(n5019), .Z(n4866) );
  IVA U4777 ( .A(n5019), .Z(n4867) );
  IVA U4778 ( .A(n5019), .Z(n4868) );
  IVA U4779 ( .A(n5020), .Z(n4869) );
  IVA U4780 ( .A(n5020), .Z(n4870) );
  IVA U4781 ( .A(n5020), .Z(n4871) );
  IVA U4782 ( .A(n5021), .Z(n4872) );
  IVA U4783 ( .A(n5021), .Z(n4873) );
  IVA U4784 ( .A(n5021), .Z(n4874) );
  IVA U4785 ( .A(n5022), .Z(n4875) );
  IVA U4786 ( .A(n5022), .Z(n4876) );
  IVA U4787 ( .A(n5022), .Z(n4877) );
  IVA U4788 ( .A(n5023), .Z(n4878) );
  IVA U4789 ( .A(n5023), .Z(n4879) );
  IVA U4790 ( .A(n5023), .Z(n4880) );
  IVA U4791 ( .A(n5024), .Z(n4881) );
  IVA U4792 ( .A(n5024), .Z(n4882) );
  IVA U4793 ( .A(n5024), .Z(n4883) );
  IVA U4794 ( .A(n4768), .Z(n4970) );
  IVA U4795 ( .A(n25), .Z(n4971) );
  IVA U4796 ( .A(n4776), .Z(n4972) );
  IVA U4797 ( .A(n25), .Z(n4973) );
  IVA U4798 ( .A(n25), .Z(n4974) );
  IVA U4799 ( .A(n4969), .Z(n4975) );
  IVA U4800 ( .A(n4969), .Z(n4976) );
  IVA U4801 ( .A(n4969), .Z(n4977) );
  IVA U4802 ( .A(n4969), .Z(n4978) );
  IVA U4803 ( .A(n4969), .Z(n4979) );
  IVA U4804 ( .A(n4770), .Z(n4980) );
  IVA U4805 ( .A(n4766), .Z(n4981) );
  IVA U4806 ( .A(n4764), .Z(n4982) );
  IVA U4807 ( .A(n4773), .Z(n4983) );
  IVA U4808 ( .A(n4778), .Z(n4984) );
  IVA U4809 ( .A(n4968), .Z(n4985) );
  IVA U4810 ( .A(n4968), .Z(n4986) );
  IVA U4811 ( .A(n4968), .Z(n4987) );
  IVA U4812 ( .A(n4968), .Z(n4988) );
  IVA U4813 ( .A(n4968), .Z(n4989) );
  IVA U4814 ( .A(n4967), .Z(n4990) );
  IVA U4815 ( .A(n4967), .Z(n4991) );
  IVA U4816 ( .A(n4967), .Z(n4992) );
  IVA U4817 ( .A(n4967), .Z(n4993) );
  IVA U4818 ( .A(n4967), .Z(n4994) );
  IVA U4819 ( .A(n4966), .Z(n4995) );
  IVA U4820 ( .A(n4966), .Z(n4996) );
  IVA U4821 ( .A(n4966), .Z(n4997) );
  IVA U4822 ( .A(n4966), .Z(n4998) );
  IVA U4823 ( .A(n4966), .Z(n4999) );
  IVA U4824 ( .A(n4965), .Z(n5000) );
  IVA U4825 ( .A(n4965), .Z(n5001) );
  IVA U4826 ( .A(n4965), .Z(n5002) );
  IVA U4827 ( .A(n4965), .Z(n5003) );
  IVA U4828 ( .A(n4965), .Z(n5004) );
  IVA U4829 ( .A(n4964), .Z(n5005) );
  IVA U4830 ( .A(n4964), .Z(n5006) );
  IVA U4831 ( .A(n4964), .Z(n5007) );
  IVA U4832 ( .A(n4964), .Z(n5008) );
  IVA U4833 ( .A(n4964), .Z(n5009) );
  IVA U4834 ( .A(n4963), .Z(n5010) );
  IVA U4835 ( .A(n4963), .Z(n5011) );
  IVA U4836 ( .A(n4963), .Z(n5012) );
  IVA U4837 ( .A(n4963), .Z(n5013) );
  IVA U4838 ( .A(n4963), .Z(n5014) );
  IVA U4839 ( .A(n4962), .Z(n5015) );
  IVA U4840 ( .A(n4962), .Z(n5016) );
  IVA U4841 ( .A(n4962), .Z(n5017) );
  IVA U4842 ( .A(n4962), .Z(n5018) );
  IVA U4843 ( .A(n4962), .Z(n5019) );
  IVA U4844 ( .A(n4961), .Z(n5020) );
  IVA U4845 ( .A(n4961), .Z(n5021) );
  IVA U4846 ( .A(n4961), .Z(n5022) );
  IVA U4847 ( .A(n4961), .Z(n5023) );
  IVA U4848 ( .A(n4961), .Z(n5024) );
  IVA U4849 ( .A(n5071), .Z(n5049) );
  IVA U4850 ( .A(n5071), .Z(n5050) );
  IVA U4851 ( .A(n5071), .Z(n5051) );
  IVA U4852 ( .A(n5071), .Z(n5052) );
  IVA U4853 ( .A(n5071), .Z(n5053) );
  IVA U4854 ( .A(n5071), .Z(n5054) );
  IVA U4855 ( .A(reset), .Z(n5071) );
  AO5 U4856 ( .A(Term1[103]), .B(Term3[15]), .C(n118), .Z(n5069) );
  IVA U4857 ( .A(n5069), .Z(n5055) );
  AO5 U4858 ( .A(Term1[104]), .B(Term3[16]), .C(n5055), .Z(n5068) );
  IVA U4859 ( .A(n5068), .Z(n5056) );
  AO5 U4860 ( .A(Term1[105]), .B(Term3[17]), .C(n5056), .Z(n5067) );
  IVA U4861 ( .A(n5067), .Z(n5057) );
  AO5 U4862 ( .A(Term1[106]), .B(Term3[18]), .C(n5057), .Z(n5066) );
  IVA U4863 ( .A(n5066), .Z(n5058) );
  AO5 U4864 ( .A(Term1[107]), .B(Term3[19]), .C(n5058), .Z(n5065) );
  IVA U4865 ( .A(n5065), .Z(n5059) );
  AO5 U4866 ( .A(Term1[108]), .B(Term3[20]), .C(n5059), .Z(n5064) );
  IVA U4867 ( .A(n5064), .Z(n5060) );
  AO5 U4868 ( .A(Term1[109]), .B(Term3[21]), .C(n5060), .Z(n5063) );
  IVA U4869 ( .A(n5063), .Z(n5061) );
  AO5 U4870 ( .A(Term1[110]), .B(Term3[22]), .C(n5061), .Z(n5062) );
  EN3P U4871 ( .A(Term1[111]), .B(Term3[23]), .C(n5062), .Z(N252) );
  EN3P U4872 ( .A(Term1[110]), .B(Term3[22]), .C(n5063), .Z(N251) );
  EN3P U4873 ( .A(Term1[109]), .B(Term3[21]), .C(n5064), .Z(N250) );
  EN3P U4874 ( .A(Term1[108]), .B(Term3[20]), .C(n5065), .Z(N249) );
  EN3P U4875 ( .A(Term1[107]), .B(Term3[19]), .C(n5066), .Z(N248) );
  EN3P U4876 ( .A(Term1[106]), .B(Term3[18]), .C(n5067), .Z(N247) );
  EN3P U4877 ( .A(Term1[105]), .B(Term3[17]), .C(n5068), .Z(N246) );
  EN3P U4878 ( .A(Term1[104]), .B(Term3[16]), .C(n5069), .Z(N245) );
  EO U4879 ( .A(Term3[15]), .B(Term1[103]), .Z(n5070) );
  EO U4880 ( .A(n118), .B(n5070), .Z(N244) );
  EO U4881 ( .A(Term3[14]), .B(Term1[102]), .Z(N243) );
  EO U4882 ( .A(Term11[118]), .B(\add_1_root_sub_1_root_add_225_2/carry[6] ), 
        .Z(N284) );
  AN2 U4883 ( .A(\add_1_root_sub_1_root_add_225_2/carry[5] ), .B(Term11[117]), 
        .Z(\add_1_root_sub_1_root_add_225_2/carry[6] ) );
  EO U4884 ( .A(Term11[117]), .B(\add_1_root_sub_1_root_add_225_2/carry[5] ), 
        .Z(N283) );
  AN2 U4885 ( .A(\add_1_root_sub_1_root_add_225_2/carry[4] ), .B(Term11[116]), 
        .Z(\add_1_root_sub_1_root_add_225_2/carry[5] ) );
  EO U4886 ( .A(Term11[116]), .B(\add_1_root_sub_1_root_add_225_2/carry[4] ), 
        .Z(N282) );
  AN2 U4887 ( .A(\add_1_root_sub_1_root_add_225_2/carry[3] ), .B(Term11[115]), 
        .Z(\add_1_root_sub_1_root_add_225_2/carry[4] ) );
  EO U4888 ( .A(Term11[115]), .B(\add_1_root_sub_1_root_add_225_2/carry[3] ), 
        .Z(N281) );
endmodule


module SQRT_POLY_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;

  wire   [13:1] carry;

  FA1A U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(SUM[13]), .S(SUM[12])
         );
  FA1A U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA1A U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA1A U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  FA1A U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA1A U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA1A U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA1A U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA1A U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA1A U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA1A U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA1A U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  EO U1 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
  AN2P U2 ( .A(A[0]), .B(B[0]), .Z(carry[1]) );
endmodule


module SQRT_POLY_DW01_add_1 ( A, B, CI, SUM, CO );
  input [40:0] A;
  input [40:0] B;
  output [40:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128;

  AN2P U2 ( .A(A[11]), .B(B[11]), .Z(n1) );
  IVP U3 ( .A(n90), .Z(n20) );
  IVP U4 ( .A(n59), .Z(n12) );
  IVP U5 ( .A(n46), .Z(n5) );
  IVP U6 ( .A(n38), .Z(n3) );
  IVP U7 ( .A(n50), .Z(n7) );
  IVP U8 ( .A(n65), .Z(n21) );
  IVP U9 ( .A(n32), .Z(n2) );
  IVP U10 ( .A(n40), .Z(n4) );
  IVP U11 ( .A(n108), .Z(n26) );
  IVP U12 ( .A(n78), .Z(n11) );
  IVP U13 ( .A(n54), .Z(n8) );
  IVP U14 ( .A(n107), .Z(n24) );
  IVP U15 ( .A(n48), .Z(n6) );
  IVP U16 ( .A(n106), .Z(n22) );
  IVP U17 ( .A(n85), .Z(n15) );
  IVP U18 ( .A(n86), .Z(n17) );
  IVP U19 ( .A(n83), .Z(n14) );
  IVP U20 ( .A(n58), .Z(n10) );
  IVP U21 ( .A(n112), .Z(n23) );
  IVP U22 ( .A(n62), .Z(n13) );
  IVP U23 ( .A(n87), .Z(n19) );
  IVP U24 ( .A(n94), .Z(n16) );
  IVP U25 ( .A(n75), .Z(n9) );
  IVP U26 ( .A(n102), .Z(n25) );
  IVP U27 ( .A(n88), .Z(n18) );
  IVP U28 ( .A(A[16]), .Z(n27) );
  IVP U29 ( .A(n128), .Z(n29) );
  IVP U30 ( .A(A[13]), .Z(n28) );
  EO U31 ( .A(n30), .B(n31), .Z(SUM[37]) );
  EO U32 ( .A(B[37]), .B(A[37]), .Z(n31) );
  AO7 U33 ( .A(n32), .B(n33), .C(n34), .Z(n30) );
  EO U34 ( .A(n35), .B(n33), .Z(SUM[36]) );
  AO6 U35 ( .A(n3), .B(n36), .C(n37), .Z(n33) );
  ND2 U36 ( .A(n2), .B(n34), .Z(n35) );
  ND2 U37 ( .A(B[36]), .B(A[36]), .Z(n34) );
  NR2 U38 ( .A(B[36]), .B(A[36]), .Z(n32) );
  EO U39 ( .A(n36), .B(n39), .Z(SUM[35]) );
  NR2 U40 ( .A(n37), .B(n38), .Z(n39) );
  NR2 U41 ( .A(B[35]), .B(A[35]), .Z(n38) );
  AN2 U42 ( .A(B[35]), .B(A[35]), .Z(n37) );
  AO7 U43 ( .A(n40), .B(n41), .C(n42), .Z(n36) );
  EO U44 ( .A(n43), .B(n41), .Z(SUM[34]) );
  AO6 U45 ( .A(n5), .B(n44), .C(n45), .Z(n41) );
  ND2 U46 ( .A(n4), .B(n42), .Z(n43) );
  ND2 U47 ( .A(B[34]), .B(A[34]), .Z(n42) );
  NR2 U48 ( .A(B[34]), .B(A[34]), .Z(n40) );
  EO U49 ( .A(n44), .B(n47), .Z(SUM[33]) );
  NR2 U50 ( .A(n45), .B(n46), .Z(n47) );
  NR2 U51 ( .A(B[33]), .B(A[33]), .Z(n46) );
  AN2 U52 ( .A(B[33]), .B(A[33]), .Z(n45) );
  AO7 U53 ( .A(n48), .B(n7), .C(n49), .Z(n44) );
  EN U54 ( .A(n51), .B(n50), .Z(SUM[32]) );
  AO7 U55 ( .A(n52), .B(n53), .C(n54), .Z(n50) );
  AO6 U56 ( .A(n55), .B(n9), .C(n56), .Z(n53) );
  AO7 U57 ( .A(n57), .B(n12), .C(n58), .Z(n55) );
  AO7 U58 ( .A(n60), .B(n61), .C(n62), .Z(n59) );
  AO6 U59 ( .A(n21), .B(n63), .C(n64), .Z(n60) );
  AO1 U60 ( .A(n66), .B(n67), .C(n68), .D(n69), .Z(n65) );
  AN3 U61 ( .A(n66), .B(n70), .C(n71), .Z(n69) );
  ND2 U62 ( .A(n6), .B(n49), .Z(n51) );
  ND2 U63 ( .A(B[32]), .B(A[32]), .Z(n49) );
  NR2 U64 ( .A(B[32]), .B(A[32]), .Z(n48) );
  EN U65 ( .A(n72), .B(n73), .Z(SUM[31]) );
  NR2 U66 ( .A(n8), .B(n52), .Z(n73) );
  NR2 U67 ( .A(B[31]), .B(A[31]), .Z(n52) );
  ND2 U68 ( .A(B[31]), .B(A[31]), .Z(n54) );
  AO6 U69 ( .A(n9), .B(n74), .C(n56), .Z(n72) );
  EO U70 ( .A(n74), .B(n76), .Z(SUM[30]) );
  NR2 U71 ( .A(n56), .B(n75), .Z(n76) );
  NR2 U72 ( .A(B[30]), .B(A[30]), .Z(n75) );
  AN2 U73 ( .A(B[30]), .B(A[30]), .Z(n56) );
  AO7 U74 ( .A(n57), .B(n11), .C(n58), .Z(n74) );
  EN U75 ( .A(n11), .B(n77), .Z(SUM[29]) );
  NR2 U76 ( .A(n10), .B(n57), .Z(n77) );
  NR2 U77 ( .A(B[29]), .B(A[29]), .Z(n57) );
  ND2 U78 ( .A(B[29]), .B(A[29]), .Z(n58) );
  AO7 U79 ( .A(n61), .B(n79), .C(n62), .Z(n78) );
  EN U80 ( .A(n79), .B(n80), .Z(SUM[28]) );
  NR2 U81 ( .A(n13), .B(n61), .Z(n80) );
  NR2 U82 ( .A(B[28]), .B(A[28]), .Z(n61) );
  ND2 U83 ( .A(B[28]), .B(A[28]), .Z(n62) );
  AO6 U84 ( .A(n20), .B(n63), .C(n64), .Z(n79) );
  AO7 U85 ( .A(n81), .B(n82), .C(n83), .Z(n64) );
  AO6 U86 ( .A(n84), .B(n15), .C(n16), .Z(n82) );
  AO7 U87 ( .A(n86), .B(n87), .C(n88), .Z(n84) );
  NR4 U88 ( .A(n81), .B(n85), .C(n86), .D(n89), .Z(n63) );
  EO U89 ( .A(n91), .B(n92), .Z(SUM[27]) );
  NR2 U90 ( .A(n14), .B(n81), .Z(n92) );
  NR2 U91 ( .A(B[27]), .B(A[27]), .Z(n81) );
  ND2 U92 ( .A(B[27]), .B(A[27]), .Z(n83) );
  AO7 U93 ( .A(n85), .B(n93), .C(n94), .Z(n91) );
  EN U94 ( .A(n93), .B(n95), .Z(SUM[26]) );
  NR2 U95 ( .A(n16), .B(n85), .Z(n95) );
  NR2 U96 ( .A(B[26]), .B(A[26]), .Z(n85) );
  ND2 U97 ( .A(B[26]), .B(A[26]), .Z(n94) );
  AO6 U98 ( .A(n17), .B(n96), .C(n18), .Z(n93) );
  EO U99 ( .A(n96), .B(n97), .Z(SUM[25]) );
  NR2 U100 ( .A(n18), .B(n86), .Z(n97) );
  NR2 U101 ( .A(B[25]), .B(A[25]), .Z(n86) );
  ND2 U102 ( .A(B[25]), .B(A[25]), .Z(n88) );
  AO7 U103 ( .A(n89), .B(n90), .C(n87), .Z(n96) );
  EN U104 ( .A(n90), .B(n98), .Z(SUM[24]) );
  NR2 U105 ( .A(n19), .B(n89), .Z(n98) );
  NR2 U106 ( .A(B[24]), .B(A[24]), .Z(n89) );
  ND2 U107 ( .A(B[24]), .B(A[24]), .Z(n87) );
  AO6 U108 ( .A(n26), .B(n66), .C(n68), .Z(n90) );
  ND2 U109 ( .A(n99), .B(n100), .Z(n68) );
  AO7 U110 ( .A(n101), .B(n23), .C(n22), .Z(n100) );
  AO6 U111 ( .A(n102), .B(n103), .C(n104), .Z(n101) );
  ND3 U112 ( .A(A[20]), .B(n24), .C(B[20]), .Z(n103) );
  NR4 U113 ( .A(n105), .B(n106), .C(n104), .D(n107), .Z(n66) );
  EN U114 ( .A(n109), .B(n110), .Z(SUM[23]) );
  ND2 U115 ( .A(n99), .B(n22), .Z(n110) );
  NR2 U116 ( .A(B[23]), .B(A[23]), .Z(n106) );
  ND2 U117 ( .A(B[23]), .B(A[23]), .Z(n99) );
  AO7 U118 ( .A(n104), .B(n111), .C(n112), .Z(n109) );
  EN U119 ( .A(n111), .B(n113), .Z(SUM[22]) );
  NR2 U120 ( .A(n23), .B(n104), .Z(n113) );
  NR2 U121 ( .A(B[22]), .B(A[22]), .Z(n104) );
  ND2 U122 ( .A(B[22]), .B(A[22]), .Z(n112) );
  AO6 U123 ( .A(n24), .B(n114), .C(n25), .Z(n111) );
  EO U124 ( .A(n114), .B(n115), .Z(SUM[21]) );
  NR2 U125 ( .A(n25), .B(n107), .Z(n115) );
  NR2 U126 ( .A(B[21]), .B(A[21]), .Z(n107) );
  ND2 U127 ( .A(B[21]), .B(A[21]), .Z(n102) );
  EON1 U128 ( .A(n105), .B(n108), .C(A[20]), .D(B[20]), .Z(n114) );
  AO6 U129 ( .A(n70), .B(n71), .C(n67), .Z(n108) );
  EON1 U130 ( .A(n116), .B(n117), .C(A[19]), .D(B[19]), .Z(n67) );
  EO1 U131 ( .A(B[18]), .B(A[18]), .C(n118), .D(n119), .Z(n117) );
  AO2 U132 ( .A(A[17]), .B(B[17]), .C(B[16]), .D(n120), .Z(n118) );
  NR2 U133 ( .A(n27), .B(n121), .Z(n120) );
  NR4 U134 ( .A(n122), .B(n116), .C(n119), .D(n121), .Z(n71) );
  NR2 U135 ( .A(B[17]), .B(A[17]), .Z(n121) );
  NR2 U136 ( .A(B[18]), .B(A[18]), .Z(n119) );
  NR2 U137 ( .A(B[19]), .B(A[19]), .Z(n116) );
  NR2 U138 ( .A(B[16]), .B(A[16]), .Z(n122) );
  EON1 U139 ( .A(n123), .B(n124), .C(A[15]), .D(B[15]), .Z(n70) );
  AO5 U140 ( .A(A[14]), .B(B[14]), .C(n125), .Z(n124) );
  EON1 U141 ( .A(n126), .B(n28), .C(B[13]), .D(n127), .Z(n125) );
  ND2 U142 ( .A(n126), .B(n28), .Z(n127) );
  AO6 U143 ( .A(n1), .B(A[12]), .C(n29), .Z(n126) );
  AO7 U144 ( .A(A[12]), .B(n1), .C(B[12]), .Z(n128) );
  NR2 U145 ( .A(A[15]), .B(B[15]), .Z(n123) );
  NR2 U146 ( .A(B[20]), .B(A[20]), .Z(n105) );
endmodule


module SQRT_POLY_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [11:0] A;
  input [30:0] B;
  output [42:0] PRODUCT;
  input TC;
  wire   \ab[11][30] , \ab[11][29] , \ab[11][28] , \ab[11][27] , \ab[11][26] ,
         \ab[11][25] , \ab[11][24] , \ab[11][23] , \ab[11][22] , \ab[11][21] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][30] , \ab[10][29] , \ab[10][28] , \ab[10][27] ,
         \ab[10][26] , \ab[10][25] , \ab[10][24] , \ab[10][23] , \ab[10][22] ,
         \ab[10][21] , \ab[10][20] , \ab[10][19] , \ab[10][18] , \ab[10][17] ,
         \ab[10][16] , \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] ,
         \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] ,
         \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] ,
         \ab[10][1] , \ab[10][0] , \ab[9][30] , \ab[9][29] , \ab[9][28] ,
         \ab[9][27] , \ab[9][26] , \ab[9][25] , \ab[9][24] , \ab[9][23] ,
         \ab[9][22] , \ab[9][21] , \ab[9][20] , \ab[9][19] , \ab[9][18] ,
         \ab[9][17] , \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] ,
         \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] ,
         \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] ,
         \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][30] , \ab[8][29] ,
         \ab[8][28] , \ab[8][27] , \ab[8][26] , \ab[8][25] , \ab[8][24] ,
         \ab[8][23] , \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] ,
         \ab[8][18] , \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][30] ,
         \ab[7][29] , \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][30] , \ab[6][29] , \ab[6][28] , \ab[6][27] , \ab[6][26] ,
         \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] , \ab[6][21] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] ,
         \ab[5][26] , \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] ,
         \ab[5][21] , \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] ,
         \ab[5][16] , \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] ,
         \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] ,
         \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] ,
         \ab[5][1] , \ab[5][0] , \ab[4][30] , \ab[4][29] , \ab[4][28] ,
         \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] , \ab[4][23] ,
         \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][30] , \ab[3][29] ,
         \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] , \ab[3][24] ,
         \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] ,
         \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][30] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] , \ab[1][26] ,
         \ab[1][25] , \ab[1][24] , \ab[1][23] , \ab[1][22] , \ab[1][21] ,
         \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] , \ab[1][16] ,
         \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] ,
         \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[0][30] , \ab[0][29] , \ab[0][28] , \ab[0][27] , \ab[0][26] ,
         \ab[0][25] , \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] ,
         \ab[0][20] , \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \CARRYB[11][29] ,
         \CARRYB[11][28] , \CARRYB[11][27] , \CARRYB[11][26] ,
         \CARRYB[11][25] , \CARRYB[11][24] , \CARRYB[11][23] ,
         \CARRYB[11][22] , \CARRYB[11][21] , \CARRYB[11][20] ,
         \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \CARRYB[11][15] , \CARRYB[11][14] ,
         \CARRYB[11][13] , \CARRYB[11][12] , \CARRYB[11][11] ,
         \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] , \CARRYB[11][7] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][29] ,
         \CARRYB[10][28] , \CARRYB[10][27] , \CARRYB[10][26] ,
         \CARRYB[10][25] , \CARRYB[10][24] , \CARRYB[10][23] ,
         \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][29] ,
         \CARRYB[9][28] , \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][25] ,
         \CARRYB[9][24] , \CARRYB[9][23] , \CARRYB[9][22] , \CARRYB[9][21] ,
         \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] ,
         \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][29] , \CARRYB[8][28] , \CARRYB[8][27] ,
         \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] , \CARRYB[8][23] ,
         \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] , \CARRYB[8][19] ,
         \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] ,
         \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] ,
         \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] ,
         \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][29] ,
         \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] ,
         \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] ,
         \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] ,
         \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] ,
         \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][29] ,
         \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] ,
         \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] ,
         \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] ,
         \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][29] , \CARRYB[4][28] , \CARRYB[4][27] ,
         \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] , \CARRYB[4][23] ,
         \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] ,
         \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] ,
         \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] ,
         \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] ,
         \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] ,
         \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][29] ,
         \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] ,
         \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] ,
         \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] ,
         \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][29] ,
         \CARRYB[1][28] , \CARRYB[1][27] , \CARRYB[1][26] , \CARRYB[1][25] ,
         \CARRYB[1][24] , \CARRYB[1][23] , \CARRYB[1][22] , \CARRYB[1][21] ,
         \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] , \CARRYB[1][17] ,
         \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[11][29] , \SUMB[11][28] , \SUMB[11][27] ,
         \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] , \SUMB[11][23] ,
         \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] , \SUMB[11][19] ,
         \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[11][0] , \SUMB[10][29] ,
         \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] , \SUMB[10][25] ,
         \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] , \SUMB[10][21] ,
         \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] ,
         \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] , \SUMB[9][26] ,
         \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] , \SUMB[9][22] ,
         \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] ,
         \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][29] ,
         \SUMB[8][28] , \SUMB[8][27] , \SUMB[8][26] , \SUMB[8][25] ,
         \SUMB[8][24] , \SUMB[8][23] , \SUMB[8][22] , \SUMB[8][21] ,
         \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] , \SUMB[8][17] ,
         \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][29] ,
         \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] , \SUMB[7][25] ,
         \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] , \SUMB[7][21] ,
         \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] , \SUMB[7][17] ,
         \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] ,
         \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] ,
         \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][29] ,
         \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] , \SUMB[6][25] ,
         \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] , \SUMB[6][21] ,
         \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] ,
         \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] ,
         \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] ,
         \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][29] ,
         \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] , \SUMB[4][25] ,
         \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] , \SUMB[4][21] ,
         \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] , \SUMB[4][17] ,
         \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] ,
         \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] ,
         \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][29] ,
         \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] , \SUMB[3][25] ,
         \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] , \SUMB[3][21] ,
         \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] , \SUMB[3][17] ,
         \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][29] ,
         \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] , \SUMB[2][25] ,
         \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] , \SUMB[2][21] ,
         \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] , \SUMB[2][17] ,
         \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] ,
         \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] ,
         \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][29] ,
         \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] , \SUMB[1][25] ,
         \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] , \SUMB[1][21] ,
         \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] , \SUMB[1][17] ,
         \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] , \SUMB[1][13] ,
         \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] , \SUMB[1][9] ,
         \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[39] , \A1[38] ,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] ,
         \A1[1] , \A1[0] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] ,
         \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , \A2[29] ,
         \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] ,
         \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] ,
         \A2[14] , \A2[13] , \A2[12] , \A2[11] , n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  SQRT_POLY_DW01_add_1 FS_1 ( .A({1'b0, \A1[39] , \A1[38] , \A1[37] , \A1[36] , 
        \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , 
        \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , 
        \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \SUMB[11][0] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , 
        \A1[0] }), .B({\A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , 
        \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , \A2[29] , 
        \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] , 
        \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , 
        \A2[14] , \A2[13] , \A2[12] , \A2[11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, PRODUCT[39:23], SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}) );
  FA1A S5_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\ab[10][30] ), .CO(
        \CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1A S3_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\ab[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1A S3_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\ab[8][30] ), .CO(
        \CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1A S3_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\ab[7][30] ), .CO(
        \CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1A S3_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\ab[6][30] ), .CO(
        \CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1A S3_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\ab[5][30] ), .CO(
        \CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA1A S3_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\ab[4][30] ), .CO(
        \CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA1A S3_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\ab[3][30] ), .CO(
        \CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1A S3_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\ab[2][30] ), .CO(
        \CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1A S3_2_29 ( .A(\ab[2][29] ), .B(\CARRYB[1][29] ), .CI(\ab[1][30] ), .CO(
        \CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1A S4_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA1A S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA1A S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1A S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1A S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA1A S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA1A S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1A S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1A S2_2_27 ( .A(\ab[2][27] ), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1A S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA1A S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1A S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1A S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA1A S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA1A S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1A S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1A S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1A S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1A S4_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1A S4_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1A S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1A S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1A S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1A S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA1A S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA1A S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1A S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1A S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA1A S2_2_25 ( .A(\ab[2][25] ), .B(\CARRYB[1][25] ), .CI(\SUMB[1][26] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1A S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1A S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA1A S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1A S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1A S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1A S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1A S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA1A S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA1A S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1A S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1A S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1A S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1A S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA1A S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA1A S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), 
        .CO(\CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA1A S4_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1A S4_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1A S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA1A S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA1A S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1A S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA1A S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA1A S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1A S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA1A S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1A S4_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1A S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA1A S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA1A S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA1A S4_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1A S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1A S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1A S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1A S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA1A S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA1A S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA1A S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA1A S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA1A S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1A S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA1A S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA1A S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1A S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA1A S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), 
        .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA1A S4_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA1A S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1A S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1A S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1A S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1A S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1A S4_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1A S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1A S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA1A S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1A S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1A S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA1A S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1A S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA1A S4_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1A S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1A S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1A S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1A S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1A S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1A S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1A S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1A S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1A S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1A S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1A S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1A S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1A S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1A S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1A S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1A S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1A S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1A S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1A S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1A S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1A S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA1A S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1A S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1A S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1A S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1A S4_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1A S4_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1A S4_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S4_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S4_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(
        \CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S4_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S4_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), .CO(
        \CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S4_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S4_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(
        \CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S4_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(
        \CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S4_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(
        \CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S4_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S4_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(
        \CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S4_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(
        \CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S4_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(
        \CARRYB[11][0] ), .S(\SUMB[11][0] ) );
  FA1A S4_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(
        \CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(
        \CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1A S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1A S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA1A S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA1A S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1A S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA1A S4_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1A S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1A S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA1A S2_2_28 ( .A(\ab[2][28] ), .B(\CARRYB[1][28] ), .CI(\SUMB[1][29] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  IVP U2 ( .A(A[0]), .Z(n17) );
  IVP U3 ( .A(A[1]), .Z(n12) );
  IVP U4 ( .A(A[2]), .Z(n11) );
  IVP U5 ( .A(A[3]), .Z(n10) );
  IVP U6 ( .A(A[4]), .Z(n9) );
  IVP U7 ( .A(A[7]), .Z(n20) );
  IVP U8 ( .A(A[8]), .Z(n13) );
  EO U9 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  EO U10 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A1[11] ) );
  EO U11 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A1[12] ) );
  EO U12 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A1[13] ) );
  EO U13 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A1[16] ) );
  EO U14 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A1[21] ) );
  EO U15 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A1[17] ) );
  EO U16 ( .A(\CARRYB[11][13] ), .B(\SUMB[11][14] ), .Z(\A1[23] ) );
  EO U17 ( .A(\CARRYB[11][12] ), .B(\SUMB[11][13] ), .Z(\A1[22] ) );
  EO U18 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A1[14] ) );
  EO U19 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A1[15] ) );
  EO U20 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A1[18] ) );
  EO U21 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A1[20] ) );
  EO U22 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A1[19] ) );
  EO U23 ( .A(\CARRYB[11][15] ), .B(\SUMB[11][16] ), .Z(\A1[25] ) );
  EO U24 ( .A(\CARRYB[11][14] ), .B(\SUMB[11][15] ), .Z(\A1[24] ) );
  EO U25 ( .A(\CARRYB[11][16] ), .B(\SUMB[11][17] ), .Z(\A1[26] ) );
  IVP U26 ( .A(A[5]), .Z(n18) );
  EO U27 ( .A(\CARRYB[11][17] ), .B(\SUMB[11][18] ), .Z(\A1[27] ) );
  EO U28 ( .A(\CARRYB[11][18] ), .B(\SUMB[11][19] ), .Z(\A1[28] ) );
  IVP U29 ( .A(A[6]), .Z(n19) );
  EO U30 ( .A(\CARRYB[11][19] ), .B(\SUMB[11][20] ), .Z(\A1[29] ) );
  EO U31 ( .A(\CARRYB[11][20] ), .B(\SUMB[11][21] ), .Z(\A1[30] ) );
  EO U32 ( .A(\CARRYB[11][21] ), .B(\SUMB[11][22] ), .Z(\A1[31] ) );
  EO U33 ( .A(\CARRYB[11][22] ), .B(\SUMB[11][23] ), .Z(\A1[32] ) );
  EO U34 ( .A(\CARRYB[11][23] ), .B(\SUMB[11][24] ), .Z(\A1[33] ) );
  EO U35 ( .A(\CARRYB[11][24] ), .B(\SUMB[11][25] ), .Z(\A1[34] ) );
  EO U36 ( .A(\CARRYB[11][25] ), .B(\SUMB[11][26] ), .Z(\A1[35] ) );
  EO U37 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Z(\SUMB[1][29] ) );
  EO U38 ( .A(\CARRYB[11][26] ), .B(\SUMB[11][27] ), .Z(\A1[36] ) );
  EO U39 ( .A(\CARRYB[11][27] ), .B(\SUMB[11][28] ), .Z(\A1[37] ) );
  IVP U40 ( .A(A[9]), .Z(n14) );
  IVP U41 ( .A(A[10]), .Z(n15) );
  IVP U42 ( .A(A[11]), .Z(n16) );
  EO U43 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A1[10] ) );
  EO U44 ( .A(\CARRYB[11][28] ), .B(\SUMB[11][29] ), .Z(\A1[38] ) );
  EO U45 ( .A(\CARRYB[11][29] ), .B(\ab[11][30] ), .Z(\A1[39] ) );
  EO U46 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U47 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U48 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U49 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U50 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U51 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U52 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U53 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U54 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U55 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U56 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U57 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U58 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U59 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U60 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Z(\SUMB[1][16] ) );
  EO U61 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Z(\SUMB[1][17] ) );
  EO U62 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Z(\SUMB[1][18] ) );
  EO U63 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Z(\SUMB[1][19] ) );
  EO U64 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Z(\SUMB[1][20] ) );
  EO U65 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Z(\SUMB[1][21] ) );
  EO U66 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Z(\SUMB[1][22] ) );
  EO U67 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Z(\SUMB[1][23] ) );
  EO U68 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Z(\SUMB[1][24] ) );
  EO U69 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Z(\SUMB[1][25] ) );
  EO U70 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Z(\SUMB[1][26] ) );
  EO U71 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Z(\SUMB[1][27] ) );
  EO U72 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Z(\SUMB[1][28] ) );
  IVP U73 ( .A(B[28]), .Z(n6) );
  IVP U74 ( .A(B[29]), .Z(n7) );
  IVP U75 ( .A(B[2]), .Z(n43) );
  IVP U76 ( .A(B[3]), .Z(n42) );
  IVP U77 ( .A(B[4]), .Z(n41) );
  IVP U78 ( .A(B[1]), .Z(n44) );
  IVP U79 ( .A(B[5]), .Z(n40) );
  IVP U80 ( .A(B[0]), .Z(n45) );
  IVP U81 ( .A(B[6]), .Z(n39) );
  IVP U82 ( .A(B[10]), .Z(n35) );
  IVP U83 ( .A(B[11]), .Z(n34) );
  IVP U84 ( .A(B[12]), .Z(n33) );
  IVP U85 ( .A(B[13]), .Z(n32) );
  IVP U86 ( .A(B[7]), .Z(n38) );
  IVP U87 ( .A(B[8]), .Z(n37) );
  IVP U88 ( .A(B[9]), .Z(n36) );
  IVP U89 ( .A(B[14]), .Z(n31) );
  IVP U90 ( .A(B[15]), .Z(n30) );
  IVP U91 ( .A(B[16]), .Z(n29) );
  IVP U92 ( .A(B[17]), .Z(n28) );
  IVP U93 ( .A(B[18]), .Z(n27) );
  IVP U94 ( .A(B[19]), .Z(n26) );
  IVP U95 ( .A(B[20]), .Z(n25) );
  IVP U96 ( .A(B[21]), .Z(n24) );
  IVP U97 ( .A(B[22]), .Z(n23) );
  IVP U98 ( .A(B[23]), .Z(n22) );
  IVP U99 ( .A(B[24]), .Z(n21) );
  IVP U100 ( .A(B[25]), .Z(n3) );
  IVP U101 ( .A(B[26]), .Z(n4) );
  IVP U102 ( .A(B[27]), .Z(n5) );
  IVP U103 ( .A(B[30]), .Z(n8) );
  AN2P U104 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A2[11] ) );
  AN2P U105 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A2[12] ) );
  AN2P U106 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A2[13] ) );
  AN2P U107 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A2[14] ) );
  AN2P U108 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A2[15] ) );
  AN2P U109 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A2[16] ) );
  AN2P U110 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A2[17] ) );
  AN2P U111 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A2[18] ) );
  AN2P U112 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A2[19] ) );
  AN2P U113 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A2[20] ) );
  AN2P U114 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A2[21] ) );
  AN2P U115 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A2[22] ) );
  AN2P U116 ( .A(\CARRYB[11][12] ), .B(\SUMB[11][13] ), .Z(\A2[23] ) );
  AN2P U117 ( .A(\CARRYB[11][13] ), .B(\SUMB[11][14] ), .Z(\A2[24] ) );
  AN2P U118 ( .A(\CARRYB[11][14] ), .B(\SUMB[11][15] ), .Z(\A2[25] ) );
  AN2P U119 ( .A(\CARRYB[11][15] ), .B(\SUMB[11][16] ), .Z(\A2[26] ) );
  AN2P U120 ( .A(\CARRYB[11][16] ), .B(\SUMB[11][17] ), .Z(\A2[27] ) );
  AN2P U121 ( .A(\CARRYB[11][17] ), .B(\SUMB[11][18] ), .Z(\A2[28] ) );
  AN2P U122 ( .A(\CARRYB[11][19] ), .B(\SUMB[11][20] ), .Z(\A2[30] ) );
  AN2P U123 ( .A(\CARRYB[11][20] ), .B(\SUMB[11][21] ), .Z(\A2[31] ) );
  AN2P U124 ( .A(\CARRYB[11][21] ), .B(\SUMB[11][22] ), .Z(\A2[32] ) );
  AN2P U125 ( .A(\CARRYB[11][22] ), .B(\SUMB[11][23] ), .Z(\A2[33] ) );
  AN2P U126 ( .A(\CARRYB[11][23] ), .B(\SUMB[11][24] ), .Z(\A2[34] ) );
  AN2P U127 ( .A(\CARRYB[11][24] ), .B(\SUMB[11][25] ), .Z(\A2[35] ) );
  AN2P U128 ( .A(\CARRYB[11][25] ), .B(\SUMB[11][26] ), .Z(\A2[36] ) );
  AN2P U129 ( .A(\CARRYB[11][26] ), .B(\SUMB[11][27] ), .Z(\A2[37] ) );
  AN2P U130 ( .A(\CARRYB[11][27] ), .B(\SUMB[11][28] ), .Z(\A2[38] ) );
  AN2P U131 ( .A(\CARRYB[11][28] ), .B(\SUMB[11][29] ), .Z(\A2[39] ) );
  AN2P U132 ( .A(\CARRYB[11][29] ), .B(\ab[11][30] ), .Z(\A2[40] ) );
  AN2P U133 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U134 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U135 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U136 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U137 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U138 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U139 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U140 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U141 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U142 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U143 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U144 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U145 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U146 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U147 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U148 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\CARRYB[1][16] ) );
  AN2P U149 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\CARRYB[1][17] ) );
  AN2P U150 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\CARRYB[1][18] ) );
  AN2P U151 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\CARRYB[1][19] ) );
  AN2P U152 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\CARRYB[1][20] ) );
  AN2P U153 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\CARRYB[1][21] ) );
  AN2P U154 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(\CARRYB[1][22] ) );
  AN2P U155 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(\CARRYB[1][23] ) );
  AN2P U156 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(\CARRYB[1][24] ) );
  AN2P U157 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(\CARRYB[1][25] ) );
  AN2P U158 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\CARRYB[1][26] ) );
  AN2P U159 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(\CARRYB[1][27] ) );
  AN2P U160 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(\CARRYB[1][28] ) );
  AN2P U161 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(\CARRYB[1][29] ) );
  AN2P U162 ( .A(\CARRYB[11][18] ), .B(\SUMB[11][19] ), .Z(\A2[29] ) );
  NR2 U164 ( .A(n14), .B(n36), .Z(\ab[9][9] ) );
  NR2 U165 ( .A(n14), .B(n37), .Z(\ab[9][8] ) );
  NR2 U166 ( .A(n14), .B(n38), .Z(\ab[9][7] ) );
  NR2 U167 ( .A(n14), .B(n39), .Z(\ab[9][6] ) );
  NR2 U168 ( .A(n14), .B(n40), .Z(\ab[9][5] ) );
  NR2 U169 ( .A(n14), .B(n41), .Z(\ab[9][4] ) );
  NR2 U170 ( .A(n14), .B(n42), .Z(\ab[9][3] ) );
  NR2 U171 ( .A(n14), .B(n8), .Z(\ab[9][30] ) );
  NR2 U172 ( .A(n14), .B(n43), .Z(\ab[9][2] ) );
  NR2 U173 ( .A(n14), .B(n7), .Z(\ab[9][29] ) );
  NR2 U174 ( .A(n14), .B(n6), .Z(\ab[9][28] ) );
  NR2 U175 ( .A(n14), .B(n5), .Z(\ab[9][27] ) );
  NR2 U176 ( .A(n14), .B(n4), .Z(\ab[9][26] ) );
  NR2 U177 ( .A(n14), .B(n3), .Z(\ab[9][25] ) );
  NR2 U178 ( .A(n14), .B(n21), .Z(\ab[9][24] ) );
  NR2 U179 ( .A(n14), .B(n22), .Z(\ab[9][23] ) );
  NR2 U180 ( .A(n14), .B(n23), .Z(\ab[9][22] ) );
  NR2 U181 ( .A(n14), .B(n24), .Z(\ab[9][21] ) );
  NR2 U182 ( .A(n14), .B(n25), .Z(\ab[9][20] ) );
  NR2 U183 ( .A(n14), .B(n44), .Z(\ab[9][1] ) );
  NR2 U184 ( .A(n14), .B(n26), .Z(\ab[9][19] ) );
  NR2 U185 ( .A(n14), .B(n27), .Z(\ab[9][18] ) );
  NR2 U186 ( .A(n14), .B(n28), .Z(\ab[9][17] ) );
  NR2 U187 ( .A(n14), .B(n29), .Z(\ab[9][16] ) );
  NR2 U188 ( .A(n14), .B(n30), .Z(\ab[9][15] ) );
  NR2 U189 ( .A(n14), .B(n31), .Z(\ab[9][14] ) );
  NR2 U190 ( .A(n14), .B(n32), .Z(\ab[9][13] ) );
  NR2 U191 ( .A(n14), .B(n33), .Z(\ab[9][12] ) );
  NR2 U192 ( .A(n14), .B(n34), .Z(\ab[9][11] ) );
  NR2 U193 ( .A(n14), .B(n35), .Z(\ab[9][10] ) );
  NR2 U194 ( .A(n14), .B(n45), .Z(\ab[9][0] ) );
  NR2 U195 ( .A(n36), .B(n13), .Z(\ab[8][9] ) );
  NR2 U196 ( .A(n37), .B(n13), .Z(\ab[8][8] ) );
  NR2 U197 ( .A(n38), .B(n13), .Z(\ab[8][7] ) );
  NR2 U198 ( .A(n39), .B(n13), .Z(\ab[8][6] ) );
  NR2 U199 ( .A(n40), .B(n13), .Z(\ab[8][5] ) );
  NR2 U200 ( .A(n41), .B(n13), .Z(\ab[8][4] ) );
  NR2 U201 ( .A(n42), .B(n13), .Z(\ab[8][3] ) );
  NR2 U202 ( .A(n8), .B(n13), .Z(\ab[8][30] ) );
  NR2 U203 ( .A(n43), .B(n13), .Z(\ab[8][2] ) );
  NR2 U204 ( .A(n7), .B(n13), .Z(\ab[8][29] ) );
  NR2 U205 ( .A(n6), .B(n13), .Z(\ab[8][28] ) );
  NR2 U206 ( .A(n5), .B(n13), .Z(\ab[8][27] ) );
  NR2 U207 ( .A(n4), .B(n13), .Z(\ab[8][26] ) );
  NR2 U208 ( .A(n3), .B(n13), .Z(\ab[8][25] ) );
  NR2 U209 ( .A(n21), .B(n13), .Z(\ab[8][24] ) );
  NR2 U210 ( .A(n22), .B(n13), .Z(\ab[8][23] ) );
  NR2 U211 ( .A(n23), .B(n13), .Z(\ab[8][22] ) );
  NR2 U212 ( .A(n24), .B(n13), .Z(\ab[8][21] ) );
  NR2 U213 ( .A(n25), .B(n13), .Z(\ab[8][20] ) );
  NR2 U214 ( .A(n44), .B(n13), .Z(\ab[8][1] ) );
  NR2 U215 ( .A(n26), .B(n13), .Z(\ab[8][19] ) );
  NR2 U216 ( .A(n27), .B(n13), .Z(\ab[8][18] ) );
  NR2 U217 ( .A(n28), .B(n13), .Z(\ab[8][17] ) );
  NR2 U218 ( .A(n29), .B(n13), .Z(\ab[8][16] ) );
  NR2 U219 ( .A(n30), .B(n13), .Z(\ab[8][15] ) );
  NR2 U220 ( .A(n31), .B(n13), .Z(\ab[8][14] ) );
  NR2 U221 ( .A(n32), .B(n13), .Z(\ab[8][13] ) );
  NR2 U222 ( .A(n33), .B(n13), .Z(\ab[8][12] ) );
  NR2 U223 ( .A(n34), .B(n13), .Z(\ab[8][11] ) );
  NR2 U224 ( .A(n35), .B(n13), .Z(\ab[8][10] ) );
  NR2 U225 ( .A(n45), .B(n13), .Z(\ab[8][0] ) );
  NR2 U226 ( .A(n36), .B(n20), .Z(\ab[7][9] ) );
  NR2 U227 ( .A(n37), .B(n20), .Z(\ab[7][8] ) );
  NR2 U228 ( .A(n38), .B(n20), .Z(\ab[7][7] ) );
  NR2 U229 ( .A(n39), .B(n20), .Z(\ab[7][6] ) );
  NR2 U230 ( .A(n40), .B(n20), .Z(\ab[7][5] ) );
  NR2 U231 ( .A(n41), .B(n20), .Z(\ab[7][4] ) );
  NR2 U232 ( .A(n42), .B(n20), .Z(\ab[7][3] ) );
  NR2 U233 ( .A(n8), .B(n20), .Z(\ab[7][30] ) );
  NR2 U234 ( .A(n43), .B(n20), .Z(\ab[7][2] ) );
  NR2 U235 ( .A(n7), .B(n20), .Z(\ab[7][29] ) );
  NR2 U236 ( .A(n6), .B(n20), .Z(\ab[7][28] ) );
  NR2 U237 ( .A(n5), .B(n20), .Z(\ab[7][27] ) );
  NR2 U238 ( .A(n4), .B(n20), .Z(\ab[7][26] ) );
  NR2 U239 ( .A(n3), .B(n20), .Z(\ab[7][25] ) );
  NR2 U240 ( .A(n21), .B(n20), .Z(\ab[7][24] ) );
  NR2 U241 ( .A(n22), .B(n20), .Z(\ab[7][23] ) );
  NR2 U242 ( .A(n23), .B(n20), .Z(\ab[7][22] ) );
  NR2 U243 ( .A(n24), .B(n20), .Z(\ab[7][21] ) );
  NR2 U244 ( .A(n25), .B(n20), .Z(\ab[7][20] ) );
  NR2 U245 ( .A(n44), .B(n20), .Z(\ab[7][1] ) );
  NR2 U246 ( .A(n26), .B(n20), .Z(\ab[7][19] ) );
  NR2 U247 ( .A(n27), .B(n20), .Z(\ab[7][18] ) );
  NR2 U248 ( .A(n28), .B(n20), .Z(\ab[7][17] ) );
  NR2 U249 ( .A(n29), .B(n20), .Z(\ab[7][16] ) );
  NR2 U250 ( .A(n30), .B(n20), .Z(\ab[7][15] ) );
  NR2 U251 ( .A(n31), .B(n20), .Z(\ab[7][14] ) );
  NR2 U252 ( .A(n32), .B(n20), .Z(\ab[7][13] ) );
  NR2 U253 ( .A(n33), .B(n20), .Z(\ab[7][12] ) );
  NR2 U254 ( .A(n34), .B(n20), .Z(\ab[7][11] ) );
  NR2 U255 ( .A(n35), .B(n20), .Z(\ab[7][10] ) );
  NR2 U256 ( .A(n45), .B(n20), .Z(\ab[7][0] ) );
  NR2 U257 ( .A(n36), .B(n19), .Z(\ab[6][9] ) );
  NR2 U258 ( .A(n37), .B(n19), .Z(\ab[6][8] ) );
  NR2 U259 ( .A(n38), .B(n19), .Z(\ab[6][7] ) );
  NR2 U260 ( .A(n39), .B(n19), .Z(\ab[6][6] ) );
  NR2 U261 ( .A(n40), .B(n19), .Z(\ab[6][5] ) );
  NR2 U262 ( .A(n41), .B(n19), .Z(\ab[6][4] ) );
  NR2 U263 ( .A(n42), .B(n19), .Z(\ab[6][3] ) );
  NR2 U264 ( .A(n8), .B(n19), .Z(\ab[6][30] ) );
  NR2 U265 ( .A(n43), .B(n19), .Z(\ab[6][2] ) );
  NR2 U266 ( .A(n7), .B(n19), .Z(\ab[6][29] ) );
  NR2 U267 ( .A(n6), .B(n19), .Z(\ab[6][28] ) );
  NR2 U268 ( .A(n5), .B(n19), .Z(\ab[6][27] ) );
  NR2 U269 ( .A(n4), .B(n19), .Z(\ab[6][26] ) );
  NR2 U270 ( .A(n3), .B(n19), .Z(\ab[6][25] ) );
  NR2 U271 ( .A(n21), .B(n19), .Z(\ab[6][24] ) );
  NR2 U272 ( .A(n22), .B(n19), .Z(\ab[6][23] ) );
  NR2 U273 ( .A(n23), .B(n19), .Z(\ab[6][22] ) );
  NR2 U274 ( .A(n24), .B(n19), .Z(\ab[6][21] ) );
  NR2 U275 ( .A(n25), .B(n19), .Z(\ab[6][20] ) );
  NR2 U276 ( .A(n44), .B(n19), .Z(\ab[6][1] ) );
  NR2 U277 ( .A(n26), .B(n19), .Z(\ab[6][19] ) );
  NR2 U278 ( .A(n27), .B(n19), .Z(\ab[6][18] ) );
  NR2 U279 ( .A(n28), .B(n19), .Z(\ab[6][17] ) );
  NR2 U280 ( .A(n29), .B(n19), .Z(\ab[6][16] ) );
  NR2 U281 ( .A(n30), .B(n19), .Z(\ab[6][15] ) );
  NR2 U282 ( .A(n31), .B(n19), .Z(\ab[6][14] ) );
  NR2 U283 ( .A(n32), .B(n19), .Z(\ab[6][13] ) );
  NR2 U284 ( .A(n33), .B(n19), .Z(\ab[6][12] ) );
  NR2 U285 ( .A(n34), .B(n19), .Z(\ab[6][11] ) );
  NR2 U286 ( .A(n35), .B(n19), .Z(\ab[6][10] ) );
  NR2 U287 ( .A(n45), .B(n19), .Z(\ab[6][0] ) );
  NR2 U288 ( .A(n36), .B(n18), .Z(\ab[5][9] ) );
  NR2 U289 ( .A(n37), .B(n18), .Z(\ab[5][8] ) );
  NR2 U290 ( .A(n38), .B(n18), .Z(\ab[5][7] ) );
  NR2 U291 ( .A(n39), .B(n18), .Z(\ab[5][6] ) );
  NR2 U292 ( .A(n40), .B(n18), .Z(\ab[5][5] ) );
  NR2 U293 ( .A(n41), .B(n18), .Z(\ab[5][4] ) );
  NR2 U294 ( .A(n42), .B(n18), .Z(\ab[5][3] ) );
  NR2 U295 ( .A(n8), .B(n18), .Z(\ab[5][30] ) );
  NR2 U296 ( .A(n43), .B(n18), .Z(\ab[5][2] ) );
  NR2 U297 ( .A(n7), .B(n18), .Z(\ab[5][29] ) );
  NR2 U298 ( .A(n6), .B(n18), .Z(\ab[5][28] ) );
  NR2 U299 ( .A(n5), .B(n18), .Z(\ab[5][27] ) );
  NR2 U300 ( .A(n4), .B(n18), .Z(\ab[5][26] ) );
  NR2 U301 ( .A(n3), .B(n18), .Z(\ab[5][25] ) );
  NR2 U302 ( .A(n21), .B(n18), .Z(\ab[5][24] ) );
  NR2 U303 ( .A(n22), .B(n18), .Z(\ab[5][23] ) );
  NR2 U304 ( .A(n23), .B(n18), .Z(\ab[5][22] ) );
  NR2 U305 ( .A(n24), .B(n18), .Z(\ab[5][21] ) );
  NR2 U306 ( .A(n25), .B(n18), .Z(\ab[5][20] ) );
  NR2 U307 ( .A(n44), .B(n18), .Z(\ab[5][1] ) );
  NR2 U308 ( .A(n26), .B(n18), .Z(\ab[5][19] ) );
  NR2 U309 ( .A(n27), .B(n18), .Z(\ab[5][18] ) );
  NR2 U310 ( .A(n28), .B(n18), .Z(\ab[5][17] ) );
  NR2 U311 ( .A(n29), .B(n18), .Z(\ab[5][16] ) );
  NR2 U312 ( .A(n30), .B(n18), .Z(\ab[5][15] ) );
  NR2 U313 ( .A(n31), .B(n18), .Z(\ab[5][14] ) );
  NR2 U314 ( .A(n32), .B(n18), .Z(\ab[5][13] ) );
  NR2 U315 ( .A(n33), .B(n18), .Z(\ab[5][12] ) );
  NR2 U316 ( .A(n34), .B(n18), .Z(\ab[5][11] ) );
  NR2 U317 ( .A(n35), .B(n18), .Z(\ab[5][10] ) );
  NR2 U318 ( .A(n45), .B(n18), .Z(\ab[5][0] ) );
  NR2 U319 ( .A(n36), .B(n9), .Z(\ab[4][9] ) );
  NR2 U320 ( .A(n37), .B(n9), .Z(\ab[4][8] ) );
  NR2 U321 ( .A(n38), .B(n9), .Z(\ab[4][7] ) );
  NR2 U322 ( .A(n39), .B(n9), .Z(\ab[4][6] ) );
  NR2 U323 ( .A(n40), .B(n9), .Z(\ab[4][5] ) );
  NR2 U324 ( .A(n41), .B(n9), .Z(\ab[4][4] ) );
  NR2 U325 ( .A(n42), .B(n9), .Z(\ab[4][3] ) );
  NR2 U326 ( .A(n8), .B(n9), .Z(\ab[4][30] ) );
  NR2 U327 ( .A(n43), .B(n9), .Z(\ab[4][2] ) );
  NR2 U328 ( .A(n7), .B(n9), .Z(\ab[4][29] ) );
  NR2 U329 ( .A(n6), .B(n9), .Z(\ab[4][28] ) );
  NR2 U330 ( .A(n5), .B(n9), .Z(\ab[4][27] ) );
  NR2 U331 ( .A(n4), .B(n9), .Z(\ab[4][26] ) );
  NR2 U332 ( .A(n3), .B(n9), .Z(\ab[4][25] ) );
  NR2 U333 ( .A(n21), .B(n9), .Z(\ab[4][24] ) );
  NR2 U334 ( .A(n22), .B(n9), .Z(\ab[4][23] ) );
  NR2 U335 ( .A(n23), .B(n9), .Z(\ab[4][22] ) );
  NR2 U336 ( .A(n24), .B(n9), .Z(\ab[4][21] ) );
  NR2 U337 ( .A(n25), .B(n9), .Z(\ab[4][20] ) );
  NR2 U338 ( .A(n44), .B(n9), .Z(\ab[4][1] ) );
  NR2 U339 ( .A(n26), .B(n9), .Z(\ab[4][19] ) );
  NR2 U340 ( .A(n27), .B(n9), .Z(\ab[4][18] ) );
  NR2 U341 ( .A(n28), .B(n9), .Z(\ab[4][17] ) );
  NR2 U342 ( .A(n29), .B(n9), .Z(\ab[4][16] ) );
  NR2 U343 ( .A(n30), .B(n9), .Z(\ab[4][15] ) );
  NR2 U344 ( .A(n31), .B(n9), .Z(\ab[4][14] ) );
  NR2 U345 ( .A(n32), .B(n9), .Z(\ab[4][13] ) );
  NR2 U346 ( .A(n33), .B(n9), .Z(\ab[4][12] ) );
  NR2 U347 ( .A(n34), .B(n9), .Z(\ab[4][11] ) );
  NR2 U348 ( .A(n35), .B(n9), .Z(\ab[4][10] ) );
  NR2 U349 ( .A(n45), .B(n9), .Z(\ab[4][0] ) );
  NR2 U350 ( .A(n36), .B(n10), .Z(\ab[3][9] ) );
  NR2 U351 ( .A(n37), .B(n10), .Z(\ab[3][8] ) );
  NR2 U352 ( .A(n38), .B(n10), .Z(\ab[3][7] ) );
  NR2 U353 ( .A(n39), .B(n10), .Z(\ab[3][6] ) );
  NR2 U354 ( .A(n40), .B(n10), .Z(\ab[3][5] ) );
  NR2 U355 ( .A(n41), .B(n10), .Z(\ab[3][4] ) );
  NR2 U356 ( .A(n42), .B(n10), .Z(\ab[3][3] ) );
  NR2 U357 ( .A(n8), .B(n10), .Z(\ab[3][30] ) );
  NR2 U358 ( .A(n43), .B(n10), .Z(\ab[3][2] ) );
  NR2 U359 ( .A(n7), .B(n10), .Z(\ab[3][29] ) );
  NR2 U360 ( .A(n6), .B(n10), .Z(\ab[3][28] ) );
  NR2 U361 ( .A(n5), .B(n10), .Z(\ab[3][27] ) );
  NR2 U362 ( .A(n4), .B(n10), .Z(\ab[3][26] ) );
  NR2 U363 ( .A(n3), .B(n10), .Z(\ab[3][25] ) );
  NR2 U364 ( .A(n21), .B(n10), .Z(\ab[3][24] ) );
  NR2 U365 ( .A(n22), .B(n10), .Z(\ab[3][23] ) );
  NR2 U366 ( .A(n23), .B(n10), .Z(\ab[3][22] ) );
  NR2 U367 ( .A(n24), .B(n10), .Z(\ab[3][21] ) );
  NR2 U368 ( .A(n25), .B(n10), .Z(\ab[3][20] ) );
  NR2 U369 ( .A(n44), .B(n10), .Z(\ab[3][1] ) );
  NR2 U370 ( .A(n26), .B(n10), .Z(\ab[3][19] ) );
  NR2 U371 ( .A(n27), .B(n10), .Z(\ab[3][18] ) );
  NR2 U372 ( .A(n28), .B(n10), .Z(\ab[3][17] ) );
  NR2 U373 ( .A(n29), .B(n10), .Z(\ab[3][16] ) );
  NR2 U374 ( .A(n30), .B(n10), .Z(\ab[3][15] ) );
  NR2 U375 ( .A(n31), .B(n10), .Z(\ab[3][14] ) );
  NR2 U376 ( .A(n32), .B(n10), .Z(\ab[3][13] ) );
  NR2 U377 ( .A(n33), .B(n10), .Z(\ab[3][12] ) );
  NR2 U378 ( .A(n34), .B(n10), .Z(\ab[3][11] ) );
  NR2 U379 ( .A(n35), .B(n10), .Z(\ab[3][10] ) );
  NR2 U380 ( .A(n45), .B(n10), .Z(\ab[3][0] ) );
  NR2 U381 ( .A(n36), .B(n11), .Z(\ab[2][9] ) );
  NR2 U382 ( .A(n37), .B(n11), .Z(\ab[2][8] ) );
  NR2 U383 ( .A(n38), .B(n11), .Z(\ab[2][7] ) );
  NR2 U384 ( .A(n39), .B(n11), .Z(\ab[2][6] ) );
  NR2 U385 ( .A(n40), .B(n11), .Z(\ab[2][5] ) );
  NR2 U386 ( .A(n41), .B(n11), .Z(\ab[2][4] ) );
  NR2 U387 ( .A(n42), .B(n11), .Z(\ab[2][3] ) );
  NR2 U388 ( .A(n8), .B(n11), .Z(\ab[2][30] ) );
  NR2 U389 ( .A(n43), .B(n11), .Z(\ab[2][2] ) );
  NR2 U390 ( .A(n7), .B(n11), .Z(\ab[2][29] ) );
  NR2 U391 ( .A(n6), .B(n11), .Z(\ab[2][28] ) );
  NR2 U392 ( .A(n5), .B(n11), .Z(\ab[2][27] ) );
  NR2 U393 ( .A(n4), .B(n11), .Z(\ab[2][26] ) );
  NR2 U394 ( .A(n3), .B(n11), .Z(\ab[2][25] ) );
  NR2 U395 ( .A(n21), .B(n11), .Z(\ab[2][24] ) );
  NR2 U396 ( .A(n22), .B(n11), .Z(\ab[2][23] ) );
  NR2 U397 ( .A(n23), .B(n11), .Z(\ab[2][22] ) );
  NR2 U398 ( .A(n24), .B(n11), .Z(\ab[2][21] ) );
  NR2 U399 ( .A(n25), .B(n11), .Z(\ab[2][20] ) );
  NR2 U400 ( .A(n44), .B(n11), .Z(\ab[2][1] ) );
  NR2 U401 ( .A(n26), .B(n11), .Z(\ab[2][19] ) );
  NR2 U402 ( .A(n27), .B(n11), .Z(\ab[2][18] ) );
  NR2 U403 ( .A(n28), .B(n11), .Z(\ab[2][17] ) );
  NR2 U404 ( .A(n29), .B(n11), .Z(\ab[2][16] ) );
  NR2 U405 ( .A(n30), .B(n11), .Z(\ab[2][15] ) );
  NR2 U406 ( .A(n31), .B(n11), .Z(\ab[2][14] ) );
  NR2 U407 ( .A(n32), .B(n11), .Z(\ab[2][13] ) );
  NR2 U408 ( .A(n33), .B(n11), .Z(\ab[2][12] ) );
  NR2 U409 ( .A(n34), .B(n11), .Z(\ab[2][11] ) );
  NR2 U410 ( .A(n35), .B(n11), .Z(\ab[2][10] ) );
  NR2 U411 ( .A(n45), .B(n11), .Z(\ab[2][0] ) );
  NR2 U412 ( .A(n36), .B(n12), .Z(\ab[1][9] ) );
  NR2 U413 ( .A(n37), .B(n12), .Z(\ab[1][8] ) );
  NR2 U414 ( .A(n38), .B(n12), .Z(\ab[1][7] ) );
  NR2 U415 ( .A(n39), .B(n12), .Z(\ab[1][6] ) );
  NR2 U416 ( .A(n40), .B(n12), .Z(\ab[1][5] ) );
  NR2 U417 ( .A(n41), .B(n12), .Z(\ab[1][4] ) );
  NR2 U418 ( .A(n42), .B(n12), .Z(\ab[1][3] ) );
  NR2 U419 ( .A(n8), .B(n12), .Z(\ab[1][30] ) );
  NR2 U420 ( .A(n43), .B(n12), .Z(\ab[1][2] ) );
  NR2 U421 ( .A(n7), .B(n12), .Z(\ab[1][29] ) );
  NR2 U422 ( .A(n6), .B(n12), .Z(\ab[1][28] ) );
  NR2 U423 ( .A(n5), .B(n12), .Z(\ab[1][27] ) );
  NR2 U424 ( .A(n4), .B(n12), .Z(\ab[1][26] ) );
  NR2 U425 ( .A(n3), .B(n12), .Z(\ab[1][25] ) );
  NR2 U426 ( .A(n21), .B(n12), .Z(\ab[1][24] ) );
  NR2 U427 ( .A(n22), .B(n12), .Z(\ab[1][23] ) );
  NR2 U428 ( .A(n23), .B(n12), .Z(\ab[1][22] ) );
  NR2 U429 ( .A(n24), .B(n12), .Z(\ab[1][21] ) );
  NR2 U430 ( .A(n25), .B(n12), .Z(\ab[1][20] ) );
  NR2 U431 ( .A(n26), .B(n12), .Z(\ab[1][19] ) );
  NR2 U432 ( .A(n27), .B(n12), .Z(\ab[1][18] ) );
  NR2 U433 ( .A(n28), .B(n12), .Z(\ab[1][17] ) );
  NR2 U434 ( .A(n29), .B(n12), .Z(\ab[1][16] ) );
  NR2 U435 ( .A(n30), .B(n12), .Z(\ab[1][15] ) );
  NR2 U436 ( .A(n31), .B(n12), .Z(\ab[1][14] ) );
  NR2 U437 ( .A(n32), .B(n12), .Z(\ab[1][13] ) );
  NR2 U438 ( .A(n33), .B(n12), .Z(\ab[1][12] ) );
  NR2 U439 ( .A(n34), .B(n12), .Z(\ab[1][11] ) );
  NR2 U440 ( .A(n35), .B(n12), .Z(\ab[1][10] ) );
  NR2 U441 ( .A(n36), .B(n16), .Z(\ab[11][9] ) );
  NR2 U442 ( .A(n37), .B(n16), .Z(\ab[11][8] ) );
  NR2 U443 ( .A(n38), .B(n16), .Z(\ab[11][7] ) );
  NR2 U444 ( .A(n39), .B(n16), .Z(\ab[11][6] ) );
  NR2 U445 ( .A(n40), .B(n16), .Z(\ab[11][5] ) );
  NR2 U446 ( .A(n41), .B(n16), .Z(\ab[11][4] ) );
  NR2 U447 ( .A(n42), .B(n16), .Z(\ab[11][3] ) );
  NR2 U448 ( .A(n8), .B(n16), .Z(\ab[11][30] ) );
  NR2 U449 ( .A(n43), .B(n16), .Z(\ab[11][2] ) );
  NR2 U450 ( .A(n7), .B(n16), .Z(\ab[11][29] ) );
  NR2 U451 ( .A(n6), .B(n16), .Z(\ab[11][28] ) );
  NR2 U452 ( .A(n5), .B(n16), .Z(\ab[11][27] ) );
  NR2 U453 ( .A(n4), .B(n16), .Z(\ab[11][26] ) );
  NR2 U454 ( .A(n3), .B(n16), .Z(\ab[11][25] ) );
  NR2 U455 ( .A(n21), .B(n16), .Z(\ab[11][24] ) );
  NR2 U456 ( .A(n22), .B(n16), .Z(\ab[11][23] ) );
  NR2 U457 ( .A(n23), .B(n16), .Z(\ab[11][22] ) );
  NR2 U458 ( .A(n24), .B(n16), .Z(\ab[11][21] ) );
  NR2 U459 ( .A(n25), .B(n16), .Z(\ab[11][20] ) );
  NR2 U460 ( .A(n44), .B(n16), .Z(\ab[11][1] ) );
  NR2 U461 ( .A(n26), .B(n16), .Z(\ab[11][19] ) );
  NR2 U462 ( .A(n27), .B(n16), .Z(\ab[11][18] ) );
  NR2 U463 ( .A(n28), .B(n16), .Z(\ab[11][17] ) );
  NR2 U464 ( .A(n29), .B(n16), .Z(\ab[11][16] ) );
  NR2 U465 ( .A(n30), .B(n16), .Z(\ab[11][15] ) );
  NR2 U466 ( .A(n31), .B(n16), .Z(\ab[11][14] ) );
  NR2 U467 ( .A(n32), .B(n16), .Z(\ab[11][13] ) );
  NR2 U468 ( .A(n33), .B(n16), .Z(\ab[11][12] ) );
  NR2 U469 ( .A(n34), .B(n16), .Z(\ab[11][11] ) );
  NR2 U470 ( .A(n35), .B(n16), .Z(\ab[11][10] ) );
  NR2 U471 ( .A(n45), .B(n16), .Z(\ab[11][0] ) );
  NR2 U472 ( .A(n36), .B(n15), .Z(\ab[10][9] ) );
  NR2 U473 ( .A(n37), .B(n15), .Z(\ab[10][8] ) );
  NR2 U474 ( .A(n38), .B(n15), .Z(\ab[10][7] ) );
  NR2 U475 ( .A(n39), .B(n15), .Z(\ab[10][6] ) );
  NR2 U476 ( .A(n40), .B(n15), .Z(\ab[10][5] ) );
  NR2 U477 ( .A(n41), .B(n15), .Z(\ab[10][4] ) );
  NR2 U478 ( .A(n42), .B(n15), .Z(\ab[10][3] ) );
  NR2 U479 ( .A(n8), .B(n15), .Z(\ab[10][30] ) );
  NR2 U480 ( .A(n43), .B(n15), .Z(\ab[10][2] ) );
  NR2 U481 ( .A(n7), .B(n15), .Z(\ab[10][29] ) );
  NR2 U482 ( .A(n6), .B(n15), .Z(\ab[10][28] ) );
  NR2 U483 ( .A(n5), .B(n15), .Z(\ab[10][27] ) );
  NR2 U484 ( .A(n4), .B(n15), .Z(\ab[10][26] ) );
  NR2 U485 ( .A(n3), .B(n15), .Z(\ab[10][25] ) );
  NR2 U486 ( .A(n21), .B(n15), .Z(\ab[10][24] ) );
  NR2 U487 ( .A(n22), .B(n15), .Z(\ab[10][23] ) );
  NR2 U488 ( .A(n23), .B(n15), .Z(\ab[10][22] ) );
  NR2 U489 ( .A(n24), .B(n15), .Z(\ab[10][21] ) );
  NR2 U490 ( .A(n25), .B(n15), .Z(\ab[10][20] ) );
  NR2 U491 ( .A(n44), .B(n15), .Z(\ab[10][1] ) );
  NR2 U492 ( .A(n26), .B(n15), .Z(\ab[10][19] ) );
  NR2 U493 ( .A(n27), .B(n15), .Z(\ab[10][18] ) );
  NR2 U494 ( .A(n28), .B(n15), .Z(\ab[10][17] ) );
  NR2 U495 ( .A(n29), .B(n15), .Z(\ab[10][16] ) );
  NR2 U496 ( .A(n30), .B(n15), .Z(\ab[10][15] ) );
  NR2 U497 ( .A(n31), .B(n15), .Z(\ab[10][14] ) );
  NR2 U498 ( .A(n32), .B(n15), .Z(\ab[10][13] ) );
  NR2 U499 ( .A(n33), .B(n15), .Z(\ab[10][12] ) );
  NR2 U500 ( .A(n34), .B(n15), .Z(\ab[10][11] ) );
  NR2 U501 ( .A(n35), .B(n15), .Z(\ab[10][10] ) );
  NR2 U502 ( .A(n45), .B(n15), .Z(\ab[10][0] ) );
  NR2 U503 ( .A(n36), .B(n17), .Z(\ab[0][9] ) );
  NR2 U504 ( .A(n37), .B(n17), .Z(\ab[0][8] ) );
  NR2 U505 ( .A(n38), .B(n17), .Z(\ab[0][7] ) );
  NR2 U506 ( .A(n39), .B(n17), .Z(\ab[0][6] ) );
  NR2 U507 ( .A(n40), .B(n17), .Z(\ab[0][5] ) );
  NR2 U508 ( .A(n41), .B(n17), .Z(\ab[0][4] ) );
  NR2 U509 ( .A(n42), .B(n17), .Z(\ab[0][3] ) );
  NR2 U510 ( .A(n8), .B(n17), .Z(\ab[0][30] ) );
  NR2 U511 ( .A(n43), .B(n17), .Z(\ab[0][2] ) );
  NR2 U512 ( .A(n7), .B(n17), .Z(\ab[0][29] ) );
  NR2 U513 ( .A(n6), .B(n17), .Z(\ab[0][28] ) );
  NR2 U514 ( .A(n5), .B(n17), .Z(\ab[0][27] ) );
  NR2 U515 ( .A(n4), .B(n17), .Z(\ab[0][26] ) );
  NR2 U516 ( .A(n3), .B(n17), .Z(\ab[0][25] ) );
  NR2 U517 ( .A(n21), .B(n17), .Z(\ab[0][24] ) );
  NR2 U518 ( .A(n22), .B(n17), .Z(\ab[0][23] ) );
  NR2 U519 ( .A(n23), .B(n17), .Z(\ab[0][22] ) );
  NR2 U520 ( .A(n24), .B(n17), .Z(\ab[0][21] ) );
  NR2 U521 ( .A(n25), .B(n17), .Z(\ab[0][20] ) );
  NR2 U522 ( .A(n26), .B(n17), .Z(\ab[0][19] ) );
  NR2 U523 ( .A(n27), .B(n17), .Z(\ab[0][18] ) );
  NR2 U524 ( .A(n28), .B(n17), .Z(\ab[0][17] ) );
  NR2 U525 ( .A(n29), .B(n17), .Z(\ab[0][16] ) );
  NR2 U526 ( .A(n30), .B(n17), .Z(\ab[0][15] ) );
  NR2 U527 ( .A(n31), .B(n17), .Z(\ab[0][14] ) );
  NR2 U528 ( .A(n32), .B(n17), .Z(\ab[0][13] ) );
  NR2 U529 ( .A(n33), .B(n17), .Z(\ab[0][12] ) );
  NR2 U530 ( .A(n34), .B(n17), .Z(\ab[0][11] ) );
  NR2 U531 ( .A(n35), .B(n17), .Z(\ab[0][10] ) );
  AN3 U532 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U533 ( .A(n12), .B(n44), .Z(\ab[1][1] ) );
endmodule


module SQRT_POLY ( clk, reset, RootIn, RootOut );
  input [30:0] RootIn;
  output [16:0] RootOut;
  input clk, reset;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N70, N71, N72, N73, n90, n91, n92, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n1, n2, n3, n4, n5, n6, n7, n8, n9, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651;
  wire   [39:23] Term1;
  wire   [19:4] Term2;
  wire   [13:0] FractionBit;
  wire   [39:36] Term11;
  wire   [19:17] Term21;
  wire   [3:0] IntegerBits;
  wire   [12:0] Root;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25;

  AN2P U1886 ( .A(Term11[37]), .B(n97), .Z(n96) );
  SQRT_POLY_DW01_add_0 add_1060 ( .A({1'b0, Term1[35:23]}), .B({1'b0, 
        Term2[16:4]}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52}) );
  SQRT_POLY_DW02_mult_0 mult_1055 ( .A({n7, n6, n5, N10, N11, N12, N13, N14, 
        N15, N16, N17, N18}), .B({RootIn[30], n648, n646, RootIn[27:0]}), .TC(
        1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25}) );
  FDS2L \Term1_reg[35]  ( .CR(1'b1), .D(N31), .LD(n643), .CP(clk), .Q(
        Term1[35]) );
  FDS2L \Term2_reg[16]  ( .CR(1'b1), .D(N39), .LD(n642), .CP(clk), .Q(
        Term2[16]) );
  FDS2L \Term1_reg[34]  ( .CR(1'b1), .D(N30), .LD(n643), .CP(clk), .Q(
        Term1[34]) );
  FDS2L \Term2_reg[15]  ( .CR(1'b1), .D(N40), .LD(n642), .CP(clk), .Q(
        Term2[15]) );
  FDS2L \Term1_reg[33]  ( .CR(1'b1), .D(N29), .LD(n643), .CP(clk), .Q(
        Term1[33]) );
  FDS2L \Term2_reg[14]  ( .CR(1'b1), .D(N41), .LD(n642), .CP(clk), .Q(
        Term2[14]) );
  FDS2L \Term1_reg[32]  ( .CR(1'b1), .D(N28), .LD(n643), .CP(clk), .Q(
        Term1[32]) );
  FDS2L \Term2_reg[13]  ( .CR(1'b1), .D(N42), .LD(n642), .CP(clk), .Q(
        Term2[13]) );
  FDS2L \Term21_reg[17]  ( .CR(1'b1), .D(Term2[17]), .LD(n639), .CP(clk), .Q(
        Term21[17]), .QN(n92) );
  FDS2L \FractionBit_reg[13]  ( .CR(1'b1), .D(N65), .LD(n641), .CP(clk), .Q(
        FractionBit[13]), .QN(n90) );
  FDS2L \Term11_reg[36]  ( .CR(1'b1), .D(Term1[36]), .LD(n640), .CP(clk), .Q(
        Term11[36]), .QN(n91) );
  FDS2L \Term1_reg[31]  ( .CR(1'b1), .D(N27), .LD(n643), .CP(clk), .Q(
        Term1[31]) );
  FDS2L \Term2_reg[12]  ( .CR(1'b1), .D(N43), .LD(n642), .CP(clk), .Q(
        Term2[12]) );
  FDS2L \Term1_reg[30]  ( .CR(1'b1), .D(N26), .LD(n643), .CP(clk), .Q(
        Term1[30]) );
  FDS2L \Term2_reg[11]  ( .CR(1'b1), .D(N44), .LD(n642), .CP(clk), .Q(
        Term2[11]) );
  FDS2L \Term1_reg[29]  ( .CR(1'b1), .D(N25), .LD(n643), .CP(clk), .Q(
        Term1[29]) );
  FDS2L \Term2_reg[10]  ( .CR(1'b1), .D(N45), .LD(n642), .CP(clk), .Q(
        Term2[10]) );
  FDS2L \Term1_reg[28]  ( .CR(1'b1), .D(N24), .LD(n643), .CP(clk), .Q(
        Term1[28]) );
  FDS2L \Term2_reg[9]  ( .CR(1'b1), .D(N46), .LD(n642), .CP(clk), .Q(Term2[9])
         );
  FDS2L \Term1_reg[27]  ( .CR(1'b1), .D(N23), .LD(n643), .CP(clk), .Q(
        Term1[27]) );
  FDS2L \Term2_reg[8]  ( .CR(1'b1), .D(N47), .LD(n641), .CP(clk), .Q(Term2[8])
         );
  FDS2L \Term1_reg[26]  ( .CR(1'b1), .D(N22), .LD(n643), .CP(clk), .Q(
        Term1[26]) );
  FDS2L \Term2_reg[7]  ( .CR(1'b1), .D(N48), .LD(n641), .CP(clk), .Q(Term2[7])
         );
  FDS2L \Term1_reg[25]  ( .CR(1'b1), .D(N21), .LD(n643), .CP(clk), .Q(
        Term1[25]) );
  FDS2L \Term2_reg[6]  ( .CR(1'b1), .D(N49), .LD(n641), .CP(clk), .Q(Term2[6])
         );
  FDS2L \Term1_reg[24]  ( .CR(1'b1), .D(N20), .LD(n643), .CP(clk), .Q(
        Term1[24]) );
  FDS2L \Term1_reg[23]  ( .CR(1'b1), .D(N19), .LD(n642), .CP(clk), .Q(
        Term1[23]) );
  FDS2L \Term2_reg[5]  ( .CR(1'b1), .D(N50), .LD(n641), .CP(clk), .Q(Term2[5])
         );
  FDS2L \Term2_reg[4]  ( .CR(1'b1), .D(N51), .LD(n641), .CP(clk), .Q(Term2[4])
         );
  FDS2L \FractionBit_reg[12]  ( .CR(1'b1), .D(N64), .LD(n641), .CP(clk), .Q(
        FractionBit[12]) );
  FDS2L \FractionBit_reg[11]  ( .CR(1'b1), .D(N63), .LD(n641), .CP(clk), .Q(
        FractionBit[11]) );
  FDS2L \FractionBit_reg[10]  ( .CR(1'b1), .D(N62), .LD(n641), .CP(clk), .Q(
        FractionBit[10]) );
  FDS2L \FractionBit_reg[9]  ( .CR(1'b1), .D(N61), .LD(n641), .CP(clk), .Q(
        FractionBit[9]) );
  FDS2L \FractionBit_reg[8]  ( .CR(1'b1), .D(N60), .LD(n641), .CP(clk), .Q(
        FractionBit[8]) );
  FDS2L \FractionBit_reg[7]  ( .CR(1'b1), .D(N59), .LD(n641), .CP(clk), .Q(
        FractionBit[7]) );
  FDS2L \FractionBit_reg[6]  ( .CR(1'b1), .D(N58), .LD(n640), .CP(clk), .Q(
        FractionBit[6]) );
  FDS2L \FractionBit_reg[5]  ( .CR(1'b1), .D(N57), .LD(n640), .CP(clk), .Q(
        FractionBit[5]) );
  FDS2L \FractionBit_reg[4]  ( .CR(1'b1), .D(N56), .LD(n640), .CP(clk), .Q(
        FractionBit[4]) );
  FDS2L \FractionBit_reg[3]  ( .CR(1'b1), .D(N55), .LD(n640), .CP(clk), .Q(
        FractionBit[3]) );
  FDS2L \FractionBit_reg[2]  ( .CR(1'b1), .D(N54), .LD(n640), .CP(clk), .Q(
        FractionBit[2]) );
  FDS2L \FractionBit_reg[1]  ( .CR(1'b1), .D(N53), .LD(n640), .CP(clk), .Q(
        FractionBit[1]) );
  FDS2L \IntegerBits_reg[3]  ( .CR(1'b1), .D(N73), .LD(n639), .CP(clk), .Q(
        IntegerBits[3]) );
  FDS2L \IntegerBits_reg[2]  ( .CR(1'b1), .D(N72), .LD(n639), .CP(clk), .Q(
        IntegerBits[2]) );
  FDS2L \IntegerBits_reg[1]  ( .CR(1'b1), .D(N71), .LD(n639), .CP(clk), .Q(
        IntegerBits[1]) );
  FDS2L \IntegerBits_reg[0]  ( .CR(1'b1), .D(N70), .LD(n639), .CP(clk), .Q(
        IntegerBits[0]) );
  FDS2L \Term1_reg[39]  ( .CR(1'b1), .D(N35), .LD(n644), .CP(clk), .Q(
        Term1[39]) );
  FDS2L \Term1_reg[38]  ( .CR(1'b1), .D(N34), .LD(n644), .CP(clk), .Q(
        Term1[38]) );
  FDS2L \Term1_reg[37]  ( .CR(1'b1), .D(N33), .LD(n644), .CP(clk), .Q(
        Term1[37]) );
  FDS2L \Term1_reg[36]  ( .CR(1'b1), .D(N32), .LD(n644), .CP(clk), .Q(
        Term1[36]) );
  FDS2L \Term2_reg[19]  ( .CR(1'b1), .D(N36), .LD(n642), .CP(clk), .Q(
        Term2[19]) );
  FDS2L \Term2_reg[18]  ( .CR(1'b1), .D(N37), .LD(n642), .CP(clk), .Q(
        Term2[18]) );
  FDS2L \Term2_reg[17]  ( .CR(1'b1), .D(N38), .LD(n642), .CP(clk), .Q(
        Term2[17]) );
  FDS2L \Term21_reg[19]  ( .CR(1'b1), .D(Term2[19]), .LD(n640), .CP(clk), .Q(
        Term21[19]) );
  FDS2L \Term21_reg[18]  ( .CR(1'b1), .D(Term2[18]), .LD(n639), .CP(clk), .Q(
        Term21[18]) );
  FDS2L \Term11_reg[39]  ( .CR(1'b1), .D(Term1[39]), .LD(n640), .CP(clk), .Q(
        Term11[39]) );
  FDS2L \Term11_reg[38]  ( .CR(1'b1), .D(Term1[38]), .LD(n640), .CP(clk), .Q(
        Term11[38]) );
  FDS2L \Term11_reg[37]  ( .CR(1'b1), .D(Term1[37]), .LD(n640), .CP(clk), .Q(
        Term11[37]) );
  FDS2L \Root_reg[12]  ( .CR(1'b1), .D(FractionBit[12]), .LD(n639), .CP(clk), 
        .Q(Root[12]) );
  FDS2L \Root_reg[11]  ( .CR(1'b1), .D(FractionBit[11]), .LD(n639), .CP(clk), 
        .Q(Root[11]) );
  FDS2L \Root_reg[10]  ( .CR(1'b1), .D(FractionBit[10]), .LD(n639), .CP(clk), 
        .Q(Root[10]) );
  FDS2L \Root_reg[9]  ( .CR(1'b1), .D(FractionBit[9]), .LD(n639), .CP(clk), 
        .Q(Root[9]) );
  FDS2L \Root_reg[8]  ( .CR(1'b1), .D(FractionBit[8]), .LD(n639), .CP(clk), 
        .Q(Root[8]) );
  FDS2L \Root_reg[7]  ( .CR(1'b1), .D(FractionBit[7]), .LD(n639), .CP(clk), 
        .Q(Root[7]) );
  FDS2L \Root_reg[6]  ( .CR(1'b1), .D(FractionBit[6]), .LD(n638), .CP(clk), 
        .Q(Root[6]) );
  FDS2L \Root_reg[5]  ( .CR(1'b1), .D(FractionBit[5]), .LD(n638), .CP(clk), 
        .Q(Root[5]) );
  FDS2L \Root_reg[4]  ( .CR(1'b1), .D(FractionBit[4]), .LD(n638), .CP(clk), 
        .Q(Root[4]) );
  FDS2L \Root_reg[3]  ( .CR(1'b1), .D(FractionBit[3]), .LD(n638), .CP(clk), 
        .Q(Root[3]) );
  FDS2L \Root_reg[2]  ( .CR(1'b1), .D(FractionBit[2]), .LD(n638), .CP(clk), 
        .Q(Root[2]) );
  FDS2L \Root_reg[1]  ( .CR(1'b1), .D(FractionBit[1]), .LD(n638), .CP(clk), 
        .Q(Root[1]) );
  FDS2L \Root_reg[0]  ( .CR(1'b1), .D(FractionBit[0]), .LD(n638), .CP(clk), 
        .Q(Root[0]) );
  FDS2L \RootOut_reg[16]  ( .CR(1'b1), .D(IntegerBits[3]), .LD(n638), .CP(clk), 
        .Q(RootOut[16]) );
  FDS2L \RootOut_reg[15]  ( .CR(1'b1), .D(IntegerBits[2]), .LD(n638), .CP(clk), 
        .Q(RootOut[15]) );
  FDS2L \RootOut_reg[14]  ( .CR(1'b1), .D(IntegerBits[1]), .LD(n638), .CP(clk), 
        .Q(RootOut[14]) );
  FDS2L \RootOut_reg[13]  ( .CR(1'b1), .D(IntegerBits[0]), .LD(n638), .CP(clk), 
        .Q(RootOut[13]) );
  FDS2L \RootOut_reg[12]  ( .CR(1'b1), .D(Root[12]), .LD(n638), .CP(clk), .Q(
        RootOut[12]) );
  FDS2L \RootOut_reg[11]  ( .CR(1'b1), .D(Root[11]), .LD(n637), .CP(clk), .Q(
        RootOut[11]) );
  FDS2L \RootOut_reg[10]  ( .CR(1'b1), .D(Root[10]), .LD(n637), .CP(clk), .Q(
        RootOut[10]) );
  FDS2L \RootOut_reg[9]  ( .CR(1'b1), .D(Root[9]), .LD(n637), .CP(clk), .Q(
        RootOut[9]) );
  FDS2L \RootOut_reg[8]  ( .CR(1'b1), .D(Root[8]), .LD(n637), .CP(clk), .Q(
        RootOut[8]) );
  FDS2L \RootOut_reg[7]  ( .CR(1'b1), .D(Root[7]), .LD(n637), .CP(clk), .Q(
        RootOut[7]) );
  FDS2L \RootOut_reg[6]  ( .CR(1'b1), .D(Root[6]), .LD(n637), .CP(clk), .Q(
        RootOut[6]) );
  FDS2L \RootOut_reg[5]  ( .CR(1'b1), .D(Root[5]), .LD(n637), .CP(clk), .Q(
        RootOut[5]) );
  FDS2L \RootOut_reg[4]  ( .CR(1'b1), .D(Root[4]), .LD(n637), .CP(clk), .Q(
        RootOut[4]) );
  FDS2L \RootOut_reg[3]  ( .CR(1'b1), .D(Root[3]), .LD(n637), .CP(clk), .Q(
        RootOut[3]) );
  FDS2L \RootOut_reg[2]  ( .CR(1'b1), .D(Root[2]), .LD(n637), .CP(clk), .Q(
        RootOut[2]) );
  FDS2L \RootOut_reg[1]  ( .CR(1'b1), .D(Root[1]), .LD(n637), .CP(clk), .Q(
        RootOut[1]) );
  FDS2L \RootOut_reg[0]  ( .CR(1'b1), .D(Root[0]), .LD(n637), .CP(clk), .Q(
        RootOut[0]) );
  FDS2L \FractionBit_reg[0]  ( .CR(1'b1), .D(N52), .LD(n640), .CP(clk), .Q(
        FractionBit[0]) );
  AN3 U3 ( .A(n518), .B(n563), .C(n622), .Z(n1) );
  AN2P U4 ( .A(n417), .B(n538), .Z(n2) );
  OR2P U5 ( .A(n586), .B(n546), .Z(n3) );
  AN2P U6 ( .A(n406), .B(n405), .Z(n4) );
  AN4P U7 ( .A(n210), .B(n491), .C(n500), .D(n506), .Z(n5) );
  AN4P U8 ( .A(n1), .B(n491), .C(n499), .D(n507), .Z(n6) );
  AN4P U9 ( .A(n209), .B(n492), .C(n498), .D(n507), .Z(n7) );
  AN2P U10 ( .A(n425), .B(n424), .Z(n8) );
  AN2P U11 ( .A(n513), .B(n561), .Z(n9) );
  ND2 U48 ( .A(n548), .B(n336), .Z(n244) );
  ND2 U49 ( .A(n626), .B(n585), .Z(n336) );
  NR2 U50 ( .A(n628), .B(n546), .Z(n300) );
  EO U51 ( .A(n620), .B(n588), .Z(n235) );
  NR3 U52 ( .A(n542), .B(n625), .C(n590), .Z(n239) );
  EN U53 ( .A(n621), .B(n548), .Z(n237) );
  NR3 U54 ( .A(n545), .B(n628), .C(n587), .Z(n220) );
  AO7 U55 ( .A(n627), .B(n587), .C(n548), .Z(n222) );
  EO U56 ( .A(n621), .B(n590), .Z(n224) );
  ND2 U57 ( .A(n398), .B(n622), .Z(n225) );
  EO U58 ( .A(n583), .B(n539), .Z(n398) );
  ND2 U59 ( .A(n376), .B(n375), .Z(n216) );
  ND2 U60 ( .A(n591), .B(n540), .Z(n375) );
  MUX21L U61 ( .A(n374), .B(n540), .S(n624), .Z(n376) );
  NR2 U62 ( .A(n591), .B(n540), .Z(n374) );
  IVP U63 ( .A(n213), .Z(n488) );
  AO7 U64 ( .A(n625), .B(n590), .C(n542), .Z(n213) );
  NR3 U65 ( .A(n543), .B(n629), .C(n589), .Z(n212) );
  NR2 U66 ( .A(n584), .B(n538), .Z(n402) );
  AN2P U67 ( .A(n592), .B(n540), .Z(n112) );
  MUX21L U68 ( .A(n629), .B(n261), .S(n589), .Z(n263) );
  NR2 U69 ( .A(n629), .B(n544), .Z(n261) );
  NR2 U70 ( .A(n592), .B(n540), .Z(n387) );
  ND2 U71 ( .A(n394), .B(n592), .Z(n148) );
  EO U72 ( .A(n621), .B(n539), .Z(n394) );
  ND2 U73 ( .A(n360), .B(n624), .Z(n161) );
  EN U74 ( .A(n583), .B(n541), .Z(n360) );
  ND2 U75 ( .A(n378), .B(n377), .Z(n126) );
  ND2 U76 ( .A(n623), .B(n540), .Z(n377) );
  EO U77 ( .A(n583), .B(n540), .Z(n378) );
  ND2 U78 ( .A(n355), .B(n354), .Z(n192) );
  AO2 U79 ( .A(n625), .B(n542), .C(n625), .D(n590), .Z(n355) );
  MUX21L U80 ( .A(n353), .B(n542), .S(n590), .Z(n354) );
  NR2 U81 ( .A(n625), .B(n542), .Z(n353) );
  ND2 U82 ( .A(n372), .B(n371), .Z(n133) );
  ND2 U83 ( .A(n368), .B(n624), .Z(n371) );
  MUX21L U84 ( .A(n369), .B(n370), .S(n624), .Z(n372) );
  NR2 U85 ( .A(n591), .B(n541), .Z(n368) );
  NR3 U86 ( .A(n545), .B(n628), .C(n587), .Z(n189) );
  AO7 U87 ( .A(n629), .B(n543), .C(n589), .Z(n172) );
  AO4 U88 ( .A(n622), .B(n539), .C(n623), .D(n592), .Z(n162) );
  NR2 U89 ( .A(n587), .B(n545), .Z(n117) );
  EO U90 ( .A(n620), .B(n544), .Z(n149) );
  EO U91 ( .A(n620), .B(n539), .Z(n134) );
  ND2 U92 ( .A(n624), .B(n541), .Z(n365) );
  ND2 U93 ( .A(n341), .B(n340), .Z(n191) );
  EO U94 ( .A(n620), .B(n548), .Z(n341) );
  EO U95 ( .A(n583), .B(n548), .Z(n340) );
  ND2 U96 ( .A(n367), .B(n366), .Z(n185) );
  ND2 U97 ( .A(n624), .B(n541), .Z(n366) );
  ND2 U98 ( .A(n591), .B(n624), .Z(n367) );
  ND2 U99 ( .A(n339), .B(n626), .Z(n167) );
  EO U100 ( .A(n583), .B(n548), .Z(n339) );
  ND2 U101 ( .A(n316), .B(n586), .Z(n151) );
  EO U102 ( .A(n621), .B(n547), .Z(n316) );
  ND2 U103 ( .A(n427), .B(n426), .Z(n128) );
  EN U104 ( .A(n620), .B(n538), .Z(n427) );
  EO U105 ( .A(n583), .B(n548), .Z(n426) );
  MUX21L U106 ( .A(n623), .B(n592), .S(n539), .Z(n186) );
  ND2 U107 ( .A(n325), .B(n324), .Z(n124) );
  ND2 U108 ( .A(n585), .B(n547), .Z(n324) );
  MUX21L U109 ( .A(n323), .B(n547), .S(n627), .Z(n325) );
  NR2 U110 ( .A(n586), .B(n547), .Z(n323) );
  EO U111 ( .A(n620), .B(n538), .Z(n418) );
  ND2 U112 ( .A(n622), .B(n537), .Z(n420) );
  ND2 U113 ( .A(n586), .B(n547), .Z(n322) );
  ND2 U114 ( .A(n628), .B(n546), .Z(n296) );
  IVP U115 ( .A(n560), .Z(n589) );
  IVP U116 ( .A(n559), .Z(n584) );
  IVP U117 ( .A(n560), .Z(n588) );
  EO U118 ( .A(n583), .B(n538), .Z(n248) );
  AO7 U119 ( .A(n590), .B(n609), .C(n527), .Z(n245) );
  NR3 U120 ( .A(n493), .B(n509), .C(n2), .Z(n438) );
  EO U121 ( .A(n620), .B(n584), .Z(n417) );
  ND2 U122 ( .A(n276), .B(n275), .Z(n242) );
  ND2 U123 ( .A(n588), .B(n544), .Z(n275) );
  MUX21L U124 ( .A(n274), .B(n617), .S(n544), .Z(n276) );
  NR2 U125 ( .A(n588), .B(n617), .Z(n274) );
  MUX21L U126 ( .A(n435), .B(n436), .S(n502), .Z(n441) );
  AN3 U127 ( .A(n254), .B(n492), .C(n508), .Z(n435) );
  AN3 U128 ( .A(n249), .B(n508), .C(N36), .Z(n436) );
  ND2 U129 ( .A(n380), .B(n379), .Z(n254) );
  ND2 U130 ( .A(n256), .B(n255), .Z(n249) );
  ND2 U131 ( .A(n528), .B(n577), .Z(n255) );
  EN U132 ( .A(n620), .B(n589), .Z(n256) );
  IVP U133 ( .A(n602), .Z(n620) );
  IVP U134 ( .A(n512), .Z(n540) );
  IVP U135 ( .A(n603), .Z(n624) );
  IVP U136 ( .A(n512), .Z(n541) );
  IVP U137 ( .A(n603), .Z(n626) );
  IVP U138 ( .A(n603), .Z(n627) );
  IVP U139 ( .A(n513), .Z(n546) );
  IVP U140 ( .A(n603), .Z(n625) );
  IVP U141 ( .A(n560), .Z(n590) );
  IVP U142 ( .A(n603), .Z(n628) );
  IVP U143 ( .A(n560), .Z(n591) );
  IVP U144 ( .A(n512), .Z(n544) );
  IVP U145 ( .A(n512), .Z(n543) );
  AN3 U146 ( .A(n252), .B(n490), .C(n508), .Z(n437) );
  AO7 U147 ( .A(n626), .B(n543), .C(n589), .Z(n252) );
  ND2 U148 ( .A(n591), .B(n522), .Z(n379) );
  ND2 U149 ( .A(n382), .B(n381), .Z(n247) );
  ND2 U150 ( .A(n623), .B(n522), .Z(n381) );
  EN U151 ( .A(n583), .B(n540), .Z(n382) );
  MUX21L U152 ( .A(n624), .B(n581), .S(n541), .Z(n253) );
  MUX21L U153 ( .A(n364), .B(n363), .S(n591), .Z(n246) );
  ND2 U154 ( .A(n624), .B(n524), .Z(n364) );
  ND2 U155 ( .A(n625), .B(n541), .Z(n363) );
  MUX21L U156 ( .A(n313), .B(n534), .S(n627), .Z(n243) );
  ND2 U157 ( .A(n586), .B(n534), .Z(n313) );
  IVP U158 ( .A(n559), .Z(n583) );
  IVP U159 ( .A(n559), .Z(n586) );
  IVP U160 ( .A(n560), .Z(n587) );
  IVP U161 ( .A(n559), .Z(n585) );
  NR2 U162 ( .A(n538), .B(n564), .Z(n241) );
  AO7 U163 ( .A(n544), .B(n617), .C(n575), .Z(n234) );
  ND2 U164 ( .A(n302), .B(n301), .Z(n236) );
  MUX21L U165 ( .A(n299), .B(n613), .S(n587), .Z(n301) );
  AO6 U166 ( .A(n587), .B(n532), .C(n300), .Z(n302) );
  ND2 U167 ( .A(n343), .B(n342), .Z(n238) );
  ND2 U168 ( .A(n528), .B(n577), .Z(n342) );
  EN U169 ( .A(n621), .B(n543), .Z(n343) );
  MUX21L U170 ( .A(n383), .B(n623), .S(n591), .Z(n240) );
  ND2 U171 ( .A(n624), .B(n522), .Z(n383) );
  IVP U172 ( .A(n511), .Z(n538) );
  IVP U173 ( .A(n602), .Z(n623) );
  IVP U174 ( .A(n513), .Z(n548) );
  IVP U175 ( .A(n512), .Z(n542) );
  IVP U176 ( .A(n602), .Z(n621) );
  IVP U177 ( .A(n490), .Z(N36) );
  ND2 U178 ( .A(n523), .B(n607), .Z(n380) );
  MUX21L U179 ( .A(n519), .B(n585), .S(n622), .Z(n233) );
  MUX21L U180 ( .A(n569), .B(n303), .S(n546), .Z(n229) );
  IVP U181 ( .A(n490), .Z(n493) );
  ND2 U182 ( .A(n346), .B(n345), .Z(n231) );
  ND2 U183 ( .A(n543), .B(n578), .Z(n345) );
  MUX21L U184 ( .A(n626), .B(n344), .S(n589), .Z(n346) );
  NR2 U185 ( .A(n626), .B(n543), .Z(n344) );
  ND2 U186 ( .A(n385), .B(n384), .Z(n232) );
  ND2 U187 ( .A(n540), .B(n607), .Z(n384) );
  EN U188 ( .A(n583), .B(n540), .Z(n385) );
  ND2 U189 ( .A(n258), .B(n257), .Z(n227) );
  ND2 U190 ( .A(n629), .B(n529), .Z(n257) );
  EN U191 ( .A(n583), .B(n543), .Z(n258) );
  IVP U192 ( .A(n513), .Z(n547) );
  IVP U193 ( .A(n603), .Z(n629) );
  ND2 U194 ( .A(n281), .B(n280), .Z(n228) );
  ND2 U195 ( .A(n588), .B(n531), .Z(n280) );
  MUX21L U196 ( .A(n279), .B(n531), .S(n628), .Z(n281) );
  NR2 U197 ( .A(n588), .B(n531), .Z(n279) );
  ND2 U198 ( .A(n330), .B(n329), .Z(n230) );
  ND2 U199 ( .A(n627), .B(n567), .Z(n329) );
  MUX21L U200 ( .A(n567), .B(n328), .S(n547), .Z(n330) );
  NR2 U201 ( .A(n627), .B(n566), .Z(n328) );
  IVP U202 ( .A(n602), .Z(n622) );
  IVP U203 ( .A(n512), .Z(n539) );
  ND2 U204 ( .A(n535), .B(n568), .Z(n221) );
  ND3 U205 ( .A(n575), .B(n616), .C(n530), .Z(n219) );
  ND2 U206 ( .A(n569), .B(n613), .Z(n303) );
  ND2 U207 ( .A(n348), .B(n347), .Z(n223) );
  ND2 U208 ( .A(n626), .B(n528), .Z(n348) );
  ND2 U209 ( .A(n589), .B(n527), .Z(n347) );
  IVP U210 ( .A(n513), .Z(n545) );
  MUX21L U211 ( .A(n622), .B(n562), .S(n537), .Z(n226) );
  AN3 U212 ( .A(n217), .B(n491), .C(n508), .Z(n445) );
  AO7 U213 ( .A(n622), .B(n539), .C(n582), .Z(n217) );
  MUX21L U214 ( .A(n447), .B(n448), .S(n493), .Z(n450) );
  NR2 U215 ( .A(n509), .B(n502), .Z(n448) );
  AN3 U216 ( .A(n501), .B(n215), .C(n508), .Z(n447) );
  NR3 U217 ( .A(n543), .B(n626), .C(n589), .Z(n215) );
  MUX21L U218 ( .A(n479), .B(n478), .S(n501), .Z(n484) );
  NR2 U219 ( .A(n509), .B(n401), .Z(n479) );
  NR2 U220 ( .A(n508), .B(n488), .Z(n478) );
  ND3 U221 ( .A(n538), .B(n564), .C(n621), .Z(n401) );
  AN3 U222 ( .A(n214), .B(N36), .C(n508), .Z(n446) );
  ND3 U223 ( .A(n574), .B(n616), .C(n530), .Z(n214) );
  MUX21L U224 ( .A(n519), .B(n584), .S(n623), .Z(n218) );
  MUX21L U225 ( .A(n493), .B(n480), .S(n508), .Z(n483) );
  NR2 U226 ( .A(n501), .B(n340), .Z(n480) );
  NR2 U227 ( .A(n502), .B(n4), .Z(n486) );
  ND2 U228 ( .A(n402), .B(n621), .Z(n405) );
  MUX21L U229 ( .A(n403), .B(n404), .S(n539), .Z(n406) );
  NR2 U230 ( .A(n622), .B(n564), .Z(n403) );
  NR2 U231 ( .A(n621), .B(n585), .Z(n404) );
  ND2 U232 ( .A(n487), .B(n491), .Z(N11) );
  MUX21L U233 ( .A(n486), .B(n485), .S(n510), .Z(n487) );
  NR2 U234 ( .A(n502), .B(n112), .Z(n485) );
  IVP U235 ( .A(n560), .Z(n592) );
  ND3 U236 ( .A(n430), .B(n429), .C(n428), .Z(N10) );
  ND2 U237 ( .A(n509), .B(n490), .Z(n429) );
  ND2 U238 ( .A(n502), .B(n491), .Z(n428) );
  ND2 U239 ( .A(n211), .B(n490), .Z(n430) );
  ND2 U240 ( .A(n408), .B(n407), .Z(n211) );
  ND2 U241 ( .A(n519), .B(n606), .Z(n408) );
  ND2 U242 ( .A(n585), .B(n518), .Z(n407) );
  NR2 U243 ( .A(n627), .B(n568), .Z(n309) );
  NR2 U244 ( .A(n591), .B(n524), .Z(n369) );
  AN3 U245 ( .A(n146), .B(n489), .C(n508), .Z(n462) );
  NR3 U246 ( .A(n542), .B(n626), .C(n589), .Z(n146) );
  ND2 U247 ( .A(n356), .B(n579), .Z(n168) );
  EO U248 ( .A(n620), .B(n542), .Z(n356) );
  ND2 U249 ( .A(n391), .B(n390), .Z(n170) );
  ND2 U250 ( .A(n521), .B(n582), .Z(n390) );
  EN U251 ( .A(n621), .B(n539), .Z(n391) );
  ND2 U252 ( .A(n362), .B(n361), .Z(n140) );
  ND2 U253 ( .A(n525), .B(n580), .Z(n361) );
  EN U254 ( .A(n620), .B(n541), .Z(n362) );
  ND2 U255 ( .A(n333), .B(n332), .Z(n198) );
  ND2 U256 ( .A(n548), .B(n566), .Z(n332) );
  MUX21L U257 ( .A(n627), .B(n331), .S(n585), .Z(n333) );
  NR2 U258 ( .A(n627), .B(n548), .Z(n331) );
  ND2 U259 ( .A(n389), .B(n388), .Z(n194) );
  MUX21L U260 ( .A(n623), .B(n386), .S(n592), .Z(n388) );
  AO6 U261 ( .A(n623), .B(n521), .C(n387), .Z(n389) );
  NR2 U262 ( .A(n623), .B(n521), .Z(n386) );
  ND2 U263 ( .A(n311), .B(n310), .Z(n182) );
  ND2 U264 ( .A(n307), .B(n612), .Z(n310) );
  MUX21L U265 ( .A(n308), .B(n309), .S(n546), .Z(n311) );
  NR2 U266 ( .A(n547), .B(n586), .Z(n307) );
  ND2 U267 ( .A(n357), .B(n526), .Z(n153) );
  EO U268 ( .A(n621), .B(n590), .Z(n357) );
  ND2 U269 ( .A(n265), .B(n264), .Z(n136) );
  ND2 U270 ( .A(n529), .B(n576), .Z(n264) );
  EN U271 ( .A(n620), .B(n544), .Z(n265) );
  ND3 U272 ( .A(n411), .B(n410), .C(n409), .Z(n202) );
  AO7 U273 ( .A(n624), .B(n540), .C(n592), .Z(n201) );
  MUX21L U274 ( .A(n589), .B(n349), .S(n626), .Z(n199) );
  ND2 U275 ( .A(n418), .B(n584), .Z(n195) );
  MUX21L U276 ( .A(n306), .B(n305), .S(n628), .Z(n190) );
  MUX21L U277 ( .A(n541), .B(n365), .S(n591), .Z(n193) );
  MUX21L U278 ( .A(n419), .B(n516), .S(n622), .Z(n187) );
  NR2 U279 ( .A(n628), .B(n574), .Z(n181) );
  MUX21L U280 ( .A(n335), .B(n334), .S(n627), .Z(n183) );
  ND2 U281 ( .A(n514), .B(n604), .Z(n171) );
  MUX21L U282 ( .A(n614), .B(n285), .S(n545), .Z(n165) );
  ND2 U283 ( .A(n591), .B(n608), .Z(n169) );
  AO7 U284 ( .A(n584), .B(n516), .C(n420), .Z(n163) );
  MUX21L U285 ( .A(n573), .B(n286), .S(n545), .Z(n157) );
  AO7 U286 ( .A(n626), .B(n565), .C(n548), .Z(n159) );
  ND2 U287 ( .A(n585), .B(n548), .Z(n152) );
  AO7 U288 ( .A(n629), .B(n561), .C(n514), .Z(n156) );
  MUX21L U289 ( .A(n592), .B(n539), .S(n623), .Z(n155) );
  EO U290 ( .A(n620), .B(n545), .Z(n137) );
  ND2 U291 ( .A(n627), .B(n322), .Z(n138) );
  ND2 U292 ( .A(n416), .B(n415), .Z(n142) );
  MUX21L U293 ( .A(n584), .B(n515), .S(n621), .Z(n135) );
  AO7 U294 ( .A(n625), .B(n542), .C(n579), .Z(n132) );
  MUX21L U295 ( .A(n586), .B(n312), .S(n627), .Z(n131) );
  AO7 U296 ( .A(n625), .B(n590), .C(n526), .Z(n125) );
  AO7 U297 ( .A(n629), .B(n588), .C(n544), .Z(n122) );
  MUX21L U298 ( .A(n546), .B(n296), .S(n587), .Z(n123) );
  MUX21H U299 ( .A(n604), .B(n515), .S(n592), .Z(n113) );
  MUX21L U300 ( .A(n460), .B(n461), .S(n502), .Z(n466) );
  AN3 U301 ( .A(n143), .B(n508), .C(N36), .Z(n461) );
  AN3 U302 ( .A(n148), .B(n490), .C(n508), .Z(n460) );
  ND2 U303 ( .A(n263), .B(n262), .Z(n143) );
  MUX21L U304 ( .A(n473), .B(n472), .S(n501), .Z(n475) );
  AN3 U305 ( .A(n119), .B(n489), .C(n508), .Z(n472) );
  NR3 U306 ( .A(n493), .B(n508), .C(n113), .Z(n473) );
  ND3 U307 ( .A(n580), .B(n609), .C(n525), .Z(n119) );
  NR3 U308 ( .A(n493), .B(n509), .C(n8), .Z(n463) );
  NR2 U309 ( .A(n423), .B(n422), .Z(n425) );
  AO7 U310 ( .A(n628), .B(n532), .C(n587), .Z(n144) );
  AO7 U311 ( .A(n545), .B(n572), .C(n290), .Z(n204) );
  ND2 U312 ( .A(n628), .B(n587), .Z(n290) );
  AO7 U313 ( .A(n626), .B(n589), .C(n536), .Z(n206) );
  AO7 U314 ( .A(n591), .B(n541), .C(n608), .Z(n154) );
  AO7 U315 ( .A(n590), .B(n542), .C(n610), .Z(n139) );
  NR2 U316 ( .A(n622), .B(n562), .Z(n422) );
  NR2 U317 ( .A(n621), .B(n515), .Z(n423) );
  AN3 U318 ( .A(n147), .B(n489), .C(n501), .Z(n458) );
  AO7 U319 ( .A(n624), .B(n541), .C(n581), .Z(n147) );
  AN3 U320 ( .A(n116), .B(n508), .C(N36), .Z(n471) );
  ND2 U321 ( .A(n278), .B(n277), .Z(n116) );
  ND2 U322 ( .A(n629), .B(n544), .Z(n278) );
  ND2 U323 ( .A(n588), .B(n545), .Z(n277) );
  AN3 U324 ( .A(n121), .B(n489), .C(n508), .Z(n470) );
  ND2 U325 ( .A(n400), .B(n399), .Z(n121) );
  ND2 U326 ( .A(n584), .B(n538), .Z(n399) );
  ND2 U327 ( .A(n622), .B(n539), .Z(n400) );
  AN3 U328 ( .A(n120), .B(n489), .C(n501), .Z(n468) );
  NR2 U329 ( .A(n590), .B(n541), .Z(n120) );
  ND2 U330 ( .A(n293), .B(n292), .Z(n173) );
  ND2 U331 ( .A(n571), .B(n614), .Z(n292) );
  MUX21L U332 ( .A(n571), .B(n291), .S(n546), .Z(n293) );
  ND3 U333 ( .A(n590), .B(n526), .C(n625), .Z(n160) );
  ND2 U334 ( .A(n544), .B(n576), .Z(n262) );
  ND2 U335 ( .A(n589), .B(n527), .Z(n349) );
  ND2 U336 ( .A(n284), .B(n283), .Z(n196) );
  ND2 U337 ( .A(n545), .B(n615), .Z(n283) );
  MUX21L U338 ( .A(n282), .B(n616), .S(n587), .Z(n284) );
  NR2 U339 ( .A(n545), .B(n615), .Z(n282) );
  ND2 U340 ( .A(n319), .B(n318), .Z(n197) );
  ND2 U341 ( .A(n534), .B(n612), .Z(n318) );
  EO U342 ( .A(n583), .B(n547), .Z(n319) );
  ND2 U343 ( .A(n359), .B(n358), .Z(n177) );
  ND2 U344 ( .A(n541), .B(n608), .Z(n358) );
  ND2 U345 ( .A(n590), .B(n609), .Z(n359) );
  ND2 U346 ( .A(n338), .B(n337), .Z(n175) );
  ND2 U347 ( .A(n536), .B(n565), .Z(n337) );
  EO U348 ( .A(n620), .B(n586), .Z(n338) );
  ND2 U349 ( .A(n260), .B(n259), .Z(n164) );
  ND2 U350 ( .A(n543), .B(n577), .Z(n260) );
  ND2 U351 ( .A(n543), .B(n619), .Z(n259) );
  ND2 U352 ( .A(n315), .B(n314), .Z(n166) );
  ND2 U353 ( .A(n547), .B(n568), .Z(n314) );
  EO U354 ( .A(n620), .B(n586), .Z(n315) );
  ND2 U355 ( .A(n321), .B(n320), .Z(n158) );
  ND2 U356 ( .A(n547), .B(n612), .Z(n320) );
  EO U357 ( .A(n583), .B(n547), .Z(n321) );
  ND2 U358 ( .A(n295), .B(n294), .Z(n150) );
  ND2 U359 ( .A(n546), .B(n571), .Z(n294) );
  EO U360 ( .A(n621), .B(n546), .Z(n295) );
  ND2 U361 ( .A(n393), .B(n392), .Z(n141) );
  ND2 U362 ( .A(n540), .B(n582), .Z(n393) );
  ND2 U363 ( .A(n539), .B(n606), .Z(n392) );
  ND2 U364 ( .A(n397), .B(n396), .Z(n127) );
  ND2 U365 ( .A(n625), .B(n592), .Z(n396) );
  MUX21L U366 ( .A(n395), .B(n520), .S(n592), .Z(n397) );
  NR2 U367 ( .A(n623), .B(n520), .Z(n395) );
  MUX21L U368 ( .A(n605), .B(n584), .S(n538), .Z(n208) );
  AO7 U369 ( .A(n542), .B(n610), .C(n578), .Z(n207) );
  ND2 U370 ( .A(n413), .B(n412), .Z(n179) );
  EN U371 ( .A(n621), .B(n586), .Z(n174) );
  AO7 U372 ( .A(n592), .B(n520), .C(n606), .Z(n178) );
  MUX21L U373 ( .A(n421), .B(n537), .S(n584), .Z(n424) );
  NR2 U374 ( .A(n537), .B(n604), .Z(n421) );
  MUX21L U375 ( .A(n546), .B(n304), .S(n587), .Z(n205) );
  ND2 U376 ( .A(n546), .B(n613), .Z(n304) );
  MUX21L U377 ( .A(n266), .B(n619), .S(n588), .Z(n203) );
  ND2 U378 ( .A(n544), .B(n619), .Z(n266) );
  MUX21L U379 ( .A(n373), .B(n523), .S(n591), .Z(n200) );
  ND2 U380 ( .A(n524), .B(n607), .Z(n373) );
  ND2 U381 ( .A(n269), .B(n268), .Z(n188) );
  ND2 U382 ( .A(n575), .B(n618), .Z(n268) );
  MUX21L U383 ( .A(n576), .B(n267), .S(n544), .Z(n269) );
  ND2 U384 ( .A(n352), .B(n351), .Z(n184) );
  ND2 U385 ( .A(n578), .B(n610), .Z(n351) );
  MUX21L U386 ( .A(n611), .B(n350), .S(n542), .Z(n352) );
  MUX21L U387 ( .A(n270), .B(n618), .S(n588), .Z(n180) );
  ND2 U388 ( .A(n544), .B(n618), .Z(n270) );
  MUX21L U389 ( .A(n626), .B(n579), .S(n542), .Z(n176) );
  ND2 U390 ( .A(n273), .B(n272), .Z(n129) );
  ND2 U391 ( .A(n629), .B(n588), .Z(n272) );
  MUX21L U392 ( .A(n271), .B(n530), .S(n588), .Z(n273) );
  NR2 U393 ( .A(n629), .B(n529), .Z(n271) );
  ND2 U394 ( .A(n289), .B(n288), .Z(n130) );
  ND2 U395 ( .A(n628), .B(n572), .Z(n288) );
  MUX21L U396 ( .A(n573), .B(n287), .S(n545), .Z(n289) );
  NR2 U397 ( .A(n628), .B(n572), .Z(n287) );
  NR3 U398 ( .A(n502), .B(n9), .C(n493), .Z(n455) );
  ND2 U399 ( .A(n586), .B(n533), .Z(n305) );
  ND2 U400 ( .A(n548), .B(n565), .Z(n334) );
  ND2 U401 ( .A(n584), .B(n516), .Z(n419) );
  ND2 U402 ( .A(n585), .B(n517), .Z(n415) );
  ND2 U403 ( .A(n586), .B(n533), .Z(n312) );
  MUX21L U404 ( .A(n414), .B(n517), .S(n621), .Z(n416) );
  NR2 U405 ( .A(n584), .B(n517), .Z(n414) );
  ND2 U406 ( .A(n457), .B(n456), .Z(N38) );
  MUX21L U407 ( .A(n454), .B(n453), .S(n493), .Z(n457) );
  MUX21L U408 ( .A(n455), .B(n502), .S(n508), .Z(n456) );
  ND2 U409 ( .A(n538), .B(n563), .Z(n409) );
  ND2 U410 ( .A(n538), .B(n605), .Z(n411) );
  ND2 U411 ( .A(n622), .B(n562), .Z(n412) );
  ND2 U412 ( .A(n623), .B(n518), .Z(n413) );
  ND2 U413 ( .A(n532), .B(n570), .Z(n114) );
  ND2 U414 ( .A(n563), .B(n605), .Z(n410) );
  ND2 U415 ( .A(n533), .B(n569), .Z(n306) );
  ND2 U416 ( .A(n536), .B(n566), .Z(n335) );
  ND2 U417 ( .A(n574), .B(n615), .Z(n285) );
  ND2 U418 ( .A(n573), .B(n614), .Z(n286) );
  ND2 U419 ( .A(n523), .B(n581), .Z(n115) );
  ND2 U420 ( .A(n432), .B(n431), .Z(N37) );
  ND2 U421 ( .A(n509), .B(n492), .Z(n432) );
  ND2 U422 ( .A(n502), .B(n492), .Z(n431) );
  ND4 U423 ( .A(n442), .B(n441), .C(n440), .D(n439), .Z(N18) );
  ND4 U424 ( .A(n253), .B(n502), .C(n492), .D(n506), .Z(n439) );
  MUX21L U425 ( .A(n433), .B(n434), .S(n509), .Z(n442) );
  MUX21L U426 ( .A(n438), .B(n437), .S(n502), .Z(n440) );
  AN3 U427 ( .A(n250), .B(n498), .C(N36), .Z(n434) );
  ND2 U428 ( .A(n298), .B(n297), .Z(n250) );
  ND2 U429 ( .A(n546), .B(n570), .Z(n297) );
  ND2 U430 ( .A(n628), .B(n570), .Z(n298) );
  AN3 U431 ( .A(n251), .B(n498), .C(N36), .Z(n433) );
  ND2 U432 ( .A(n327), .B(n326), .Z(n251) );
  ND2 U433 ( .A(n585), .B(n535), .Z(n327) );
  ND2 U434 ( .A(n585), .B(n611), .Z(n326) );
  IVP U435 ( .A(n495), .Z(n490) );
  IVP U436 ( .A(n505), .Z(n508) );
  IVP U437 ( .A(n500), .Z(n502) );
  IVP U438 ( .A(n506), .Z(n509) );
  IVP U439 ( .A(n496), .Z(n492) );
  ND4 U440 ( .A(n452), .B(n451), .C(n450), .D(n449), .Z(N13) );
  ND3 U441 ( .A(n218), .B(n505), .C(n499), .Z(n449) );
  MUX21L U442 ( .A(n445), .B(n446), .S(n502), .Z(n451) );
  MUX21L U443 ( .A(n443), .B(n444), .S(n493), .Z(n452) );
  NR2 U444 ( .A(n502), .B(n3), .Z(n444) );
  AN3 U445 ( .A(n216), .B(n504), .C(n501), .Z(n443) );
  IVP U446 ( .A(n498), .Z(n503) );
  ND4 U447 ( .A(n484), .B(n483), .C(n482), .D(n481), .Z(N12) );
  ND2 U448 ( .A(n493), .B(n500), .Z(n482) );
  ND2 U449 ( .A(n212), .B(n493), .Z(n481) );
  IVP U450 ( .A(n499), .Z(n501) );
  IVP U451 ( .A(n507), .Z(n510) );
  IVP U452 ( .A(n496), .Z(n491) );
  ND2 U453 ( .A(n514), .B(n561), .Z(n210) );
  NR3 U454 ( .A(n538), .B(n621), .C(n585), .Z(n209) );
  ND4 U455 ( .A(n467), .B(n466), .C(n465), .D(n464), .Z(N43) );
  ND4 U456 ( .A(n144), .B(n493), .C(n501), .D(n505), .Z(n464) );
  MUX21L U457 ( .A(n458), .B(n459), .S(n509), .Z(n467) );
  MUX21L U458 ( .A(n463), .B(n462), .S(n501), .Z(n465) );
  ND4 U459 ( .A(n477), .B(n476), .C(n475), .D(n474), .Z(N39) );
  ND4 U460 ( .A(n117), .B(n493), .C(n502), .D(n504), .Z(n474) );
  MUX21L U461 ( .A(n468), .B(n469), .S(n508), .Z(n477) );
  MUX21L U462 ( .A(n470), .B(n471), .S(n501), .Z(n476) );
  AN3 U463 ( .A(n145), .B(n497), .C(N36), .Z(n459) );
  ND2 U464 ( .A(n547), .B(n317), .Z(n145) );
  ND2 U465 ( .A(n627), .B(n587), .Z(n317) );
  AN3 U466 ( .A(n118), .B(n497), .C(N36), .Z(n469) );
  ND3 U467 ( .A(n567), .B(n611), .C(n535), .Z(n118) );
  IVP U468 ( .A(n495), .Z(n489) );
  IVP U469 ( .A(n645), .Z(n637) );
  IVP U470 ( .A(n645), .Z(n638) );
  IVP U471 ( .A(n645), .Z(n639) );
  IVP U472 ( .A(n645), .Z(n640) );
  IVP U473 ( .A(n645), .Z(n641) );
  IVP U474 ( .A(n645), .Z(n642) );
  IVP U475 ( .A(n645), .Z(n643) );
  AO5 U476 ( .A(n91), .B(n90), .C(n92), .Z(n97) );
  EN U477 ( .A(Term11[39]), .B(n94), .Z(N73) );
  AO5 U478 ( .A(n650), .B(Term11[38]), .C(Term21[19]), .Z(n94) );
  IVP U479 ( .A(n95), .Z(n650) );
  AO4 U480 ( .A(n96), .B(Term21[18]), .C(n97), .D(Term11[37]), .Z(n95) );
  ND2 U481 ( .A(Term11[36]), .B(FractionBit[13]), .Z(n101) );
  EN U482 ( .A(n97), .B(n102), .Z(N71) );
  EN U483 ( .A(Term11[37]), .B(Term21[18]), .Z(n102) );
  EO U484 ( .A(n98), .B(n99), .Z(N72) );
  EN U485 ( .A(Term11[38]), .B(Term21[19]), .Z(n99) );
  AO5 U486 ( .A(Term11[37]), .B(n100), .C(Term21[18]), .Z(n98) );
  AO2 U487 ( .A(n101), .B(n92), .C(n90), .D(n91), .Z(n100) );
  EO U488 ( .A(FractionBit[13]), .B(n103), .Z(N70) );
  EO U489 ( .A(Term21[17]), .B(Term11[36]), .Z(n103) );
  IVP U490 ( .A(n651), .Z(n645) );
  IVP U491 ( .A(reset), .Z(n651) );
  MUX81P U492 ( .D0(n128), .D1(n543), .D2(n126), .D3(n123), .D4(n127), .D5(
        n124), .D6(n125), .D7(n122), .A(N36), .B(n503), .C(n509), .Z(N40) );
  MUX81P U493 ( .D0(n135), .D1(n585), .D2(n133), .D3(n130), .D4(n134), .D5(
        n131), .D6(n132), .D7(n129), .A(N36), .B(n503), .C(n510), .Z(N41) );
  MUX81P U494 ( .D0(n142), .D1(n629), .D2(n140), .D3(n137), .D4(n141), .D5(
        n138), .D6(n139), .D7(n136), .A(N36), .B(n503), .C(n510), .Z(N42) );
  MUX81P U495 ( .D0(n156), .D1(n152), .D2(n154), .D3(n150), .D4(n155), .D5(
        n151), .D6(n153), .D7(n149), .A(N36), .B(n503), .C(n510), .Z(N44) );
  MUX81P U496 ( .D0(n163), .D1(n159), .D2(n161), .D3(n157), .D4(n162), .D5(
        n158), .D6(n160), .D7(n543), .A(N36), .B(n503), .C(n510), .Z(N45) );
  MUX81P U497 ( .D0(n171), .D1(n167), .D2(n169), .D3(n165), .D4(n170), .D5(
        n166), .D6(n168), .D7(n164), .A(N36), .B(n503), .C(n510), .Z(N46) );
  MUX81P U498 ( .D0(n179), .D1(n175), .D2(n177), .D3(n173), .D4(n178), .D5(
        n174), .D6(n176), .D7(n172), .A(N36), .B(n503), .C(n510), .Z(N47) );
  MUX81P U499 ( .D0(n187), .D1(n183), .D2(n185), .D3(n181), .D4(n186), .D5(
        n182), .D6(n184), .D7(n180), .A(N36), .B(n503), .C(n510), .Z(N48) );
  MUX81P U500 ( .D0(n195), .D1(n191), .D2(n193), .D3(n189), .D4(n194), .D5(
        n190), .D6(n192), .D7(n188), .A(N36), .B(n503), .C(n510), .Z(N49) );
  MUX81P U501 ( .D0(n202), .D1(n198), .D2(n200), .D3(n196), .D4(n201), .D5(
        n197), .D6(n199), .D7(n545), .A(N36), .B(n503), .C(n510), .Z(N50) );
  MUX81P U502 ( .D0(n208), .D1(n206), .D2(n1), .D3(n204), .D4(n588), .D5(n205), 
        .D6(n207), .D7(n203), .A(N36), .B(n503), .C(n510), .Z(N51) );
  MUX81P U503 ( .D0(n226), .D1(n222), .D2(n224), .D3(n220), .D4(n225), .D5(
        n221), .D6(n223), .D7(n219), .A(N36), .B(n503), .C(n510), .Z(N14) );
  MUX81P U504 ( .D0(n233), .D1(n230), .D2(n629), .D3(n228), .D4(n232), .D5(
        n229), .D6(n231), .D7(n227), .A(N36), .B(n502), .C(n509), .Z(N15) );
  MUX81P U505 ( .D0(n241), .D1(n237), .D2(n239), .D3(n235), .D4(n240), .D5(
        n236), .D6(n238), .D7(n234), .A(N36), .B(n502), .C(n509), .Z(N16) );
  MUX81P U506 ( .D0(n248), .D1(n244), .D2(n246), .D3(n625), .D4(n247), .D5(
        n243), .D6(n245), .D7(n242), .A(N36), .B(n502), .C(n509), .Z(N17) );
  AN2P U507 ( .A(n620), .B(n583), .Z(n267) );
  AN2P U508 ( .A(n620), .B(n584), .Z(n291) );
  AN2P U509 ( .A(n620), .B(n537), .Z(n299) );
  AN2P U510 ( .A(n621), .B(n584), .Z(n308) );
  AN2P U511 ( .A(n620), .B(n583), .Z(n350) );
  AN2P U512 ( .A(n583), .B(n537), .Z(n370) );
  AN2P U513 ( .A(n114), .B(n501), .Z(n453) );
  AN2P U514 ( .A(n115), .B(n501), .Z(n454) );
  IVA U515 ( .A(RootIn[30]), .Z(n494) );
  IVP U516 ( .A(n494), .Z(n495) );
  IVP U517 ( .A(n494), .Z(n496) );
  IVA U518 ( .A(n648), .Z(n497) );
  IVA U519 ( .A(n648), .Z(n498) );
  IVA U520 ( .A(n648), .Z(n499) );
  IVA U521 ( .A(n648), .Z(n500) );
  IVA U522 ( .A(n646), .Z(n504) );
  IVA U523 ( .A(n646), .Z(n505) );
  IVA U524 ( .A(n646), .Z(n506) );
  IVA U525 ( .A(n646), .Z(n507) );
  IVA U526 ( .A(n550), .Z(n511) );
  IVA U527 ( .A(n550), .Z(n512) );
  IVA U528 ( .A(n551), .Z(n513) );
  IVA U529 ( .A(n551), .Z(n514) );
  IVA U530 ( .A(n551), .Z(n515) );
  IVA U531 ( .A(n552), .Z(n516) );
  IVA U532 ( .A(n552), .Z(n517) );
  IVA U533 ( .A(n552), .Z(n518) );
  IVA U534 ( .A(n553), .Z(n519) );
  IVA U535 ( .A(n553), .Z(n520) );
  IVA U536 ( .A(n553), .Z(n521) );
  IVA U537 ( .A(n554), .Z(n522) );
  IVA U538 ( .A(n554), .Z(n523) );
  IVA U539 ( .A(n554), .Z(n524) );
  IVA U540 ( .A(n555), .Z(n525) );
  IVA U541 ( .A(n555), .Z(n526) );
  IVA U542 ( .A(n555), .Z(n527) );
  IVA U543 ( .A(n556), .Z(n528) );
  IVA U544 ( .A(n556), .Z(n529) );
  IVA U545 ( .A(n556), .Z(n530) );
  IVA U546 ( .A(n557), .Z(n531) );
  IVA U547 ( .A(n557), .Z(n532) );
  IVA U548 ( .A(n557), .Z(n533) );
  IVA U549 ( .A(n558), .Z(n534) );
  IVA U550 ( .A(n558), .Z(n535) );
  IVA U551 ( .A(n558), .Z(n536) );
  IV U552 ( .A(n511), .Z(n537) );
  IVA U553 ( .A(RootIn[27]), .Z(n549) );
  IVA U554 ( .A(n549), .Z(n550) );
  IVA U555 ( .A(n549), .Z(n551) );
  IVA U556 ( .A(n549), .Z(n552) );
  IVA U557 ( .A(n517), .Z(n553) );
  IVA U558 ( .A(n511), .Z(n554) );
  IVA U559 ( .A(n515), .Z(n555) );
  IVA U560 ( .A(n511), .Z(n556) );
  IVA U561 ( .A(n518), .Z(n557) );
  IVA U562 ( .A(n514), .Z(n558) );
  IVA U563 ( .A(n594), .Z(n559) );
  IVA U564 ( .A(n594), .Z(n560) );
  IVA U565 ( .A(n594), .Z(n561) );
  IVA U566 ( .A(n595), .Z(n562) );
  IVA U567 ( .A(n595), .Z(n563) );
  IVA U568 ( .A(n595), .Z(n564) );
  IVA U569 ( .A(n596), .Z(n565) );
  IVA U570 ( .A(n596), .Z(n566) );
  IVA U571 ( .A(n596), .Z(n567) );
  IVA U572 ( .A(n597), .Z(n568) );
  IVA U573 ( .A(n597), .Z(n569) );
  IVA U574 ( .A(n597), .Z(n570) );
  IVA U575 ( .A(n598), .Z(n571) );
  IVA U576 ( .A(n598), .Z(n572) );
  IVA U577 ( .A(n598), .Z(n573) );
  IVA U578 ( .A(n599), .Z(n574) );
  IVA U579 ( .A(n599), .Z(n575) );
  IVA U580 ( .A(n599), .Z(n576) );
  IVA U581 ( .A(n600), .Z(n577) );
  IVA U582 ( .A(n600), .Z(n578) );
  IVA U583 ( .A(n600), .Z(n579) );
  IVA U584 ( .A(n601), .Z(n580) );
  IVA U585 ( .A(n601), .Z(n581) );
  IVA U586 ( .A(n601), .Z(n582) );
  IVA U587 ( .A(RootIn[26]), .Z(n593) );
  IVA U588 ( .A(n593), .Z(n594) );
  IVA U589 ( .A(n593), .Z(n595) );
  IVA U590 ( .A(n593), .Z(n596) );
  IVA U591 ( .A(n561), .Z(n597) );
  IVA U592 ( .A(n565), .Z(n598) );
  IVA U593 ( .A(n563), .Z(n599) );
  IVA U594 ( .A(n566), .Z(n600) );
  IVA U595 ( .A(n564), .Z(n601) );
  IVA U596 ( .A(n631), .Z(n602) );
  IVA U597 ( .A(n631), .Z(n603) );
  IVA U598 ( .A(n631), .Z(n604) );
  IVA U599 ( .A(n632), .Z(n605) );
  IVA U600 ( .A(n632), .Z(n606) );
  IVA U601 ( .A(n632), .Z(n607) );
  IVA U602 ( .A(n633), .Z(n608) );
  IVA U603 ( .A(n633), .Z(n609) );
  IVA U604 ( .A(n633), .Z(n610) );
  IVA U605 ( .A(n634), .Z(n611) );
  IVA U606 ( .A(n634), .Z(n612) );
  IVA U607 ( .A(n634), .Z(n613) );
  IVA U608 ( .A(n635), .Z(n614) );
  IVA U609 ( .A(n635), .Z(n615) );
  IVA U610 ( .A(n635), .Z(n616) );
  IVA U611 ( .A(n636), .Z(n617) );
  IVA U612 ( .A(n636), .Z(n618) );
  IVA U613 ( .A(n636), .Z(n619) );
  IVA U614 ( .A(RootIn[25]), .Z(n630) );
  IVA U615 ( .A(n630), .Z(n631) );
  IVA U616 ( .A(n630), .Z(n632) );
  IVA U617 ( .A(n630), .Z(n633) );
  IVA U618 ( .A(n607), .Z(n634) );
  IVA U619 ( .A(n606), .Z(n635) );
  IVA U620 ( .A(n609), .Z(n636) );
  IV U621 ( .A(n645), .Z(n644) );
  IVA U622 ( .A(n647), .Z(n646) );
  IV U623 ( .A(RootIn[28]), .Z(n647) );
  IVA U624 ( .A(n649), .Z(n648) );
  IV U625 ( .A(RootIn[29]), .Z(n649) );
endmodule


module SinBlock_0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   \A[9] , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59;
  assign SUM[10] = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];

  OR2P U2 ( .A(B[11]), .B(A[11]), .Z(n1) );
  AN2P U3 ( .A(n1), .B(n59), .Z(SUM[11]) );
  IVP U4 ( .A(n57), .Z(n13) );
  IVP U5 ( .A(n50), .Z(n11) );
  IVP U6 ( .A(n42), .Z(n9) );
  IVP U7 ( .A(n34), .Z(n7) );
  IVP U8 ( .A(n26), .Z(n5) );
  IVP U9 ( .A(n59), .Z(n14) );
  IVP U10 ( .A(n22), .Z(n4) );
  IVP U11 ( .A(n30), .Z(n6) );
  IVP U12 ( .A(n38), .Z(n8) );
  IVP U13 ( .A(n46), .Z(n10) );
  IVP U14 ( .A(n54), .Z(n12) );
  IVP U15 ( .A(n18), .Z(n3) );
  EN U16 ( .A(B[23]), .B(n15), .Z(SUM[23]) );
  AO6 U17 ( .A(n16), .B(n3), .C(n17), .Z(n15) );
  EO U18 ( .A(n16), .B(n19), .Z(SUM[22]) );
  NR2 U19 ( .A(n17), .B(n18), .Z(n19) );
  NR2 U20 ( .A(B[22]), .B(A[22]), .Z(n18) );
  AN2 U21 ( .A(B[22]), .B(A[22]), .Z(n17) );
  AO7 U22 ( .A(n20), .B(n21), .C(n22), .Z(n16) );
  EN U23 ( .A(n21), .B(n23), .Z(SUM[21]) );
  NR2 U24 ( .A(n4), .B(n20), .Z(n23) );
  NR2 U25 ( .A(B[21]), .B(A[21]), .Z(n20) );
  ND2 U26 ( .A(B[21]), .B(A[21]), .Z(n22) );
  AO6 U27 ( .A(n5), .B(n24), .C(n25), .Z(n21) );
  EO U28 ( .A(n24), .B(n27), .Z(SUM[20]) );
  NR2 U29 ( .A(n25), .B(n26), .Z(n27) );
  NR2 U30 ( .A(B[20]), .B(A[20]), .Z(n26) );
  AN2 U31 ( .A(B[20]), .B(A[20]), .Z(n25) );
  AO7 U32 ( .A(n28), .B(n29), .C(n30), .Z(n24) );
  EN U33 ( .A(n29), .B(n31), .Z(SUM[19]) );
  NR2 U34 ( .A(n6), .B(n28), .Z(n31) );
  NR2 U35 ( .A(B[19]), .B(A[19]), .Z(n28) );
  ND2 U36 ( .A(B[19]), .B(A[19]), .Z(n30) );
  AO6 U37 ( .A(n7), .B(n32), .C(n33), .Z(n29) );
  EO U38 ( .A(n32), .B(n35), .Z(SUM[18]) );
  NR2 U39 ( .A(n33), .B(n34), .Z(n35) );
  NR2 U40 ( .A(B[18]), .B(A[18]), .Z(n34) );
  AN2 U41 ( .A(B[18]), .B(A[18]), .Z(n33) );
  AO7 U42 ( .A(n36), .B(n37), .C(n38), .Z(n32) );
  EN U43 ( .A(n37), .B(n39), .Z(SUM[17]) );
  NR2 U44 ( .A(n8), .B(n36), .Z(n39) );
  NR2 U45 ( .A(B[17]), .B(A[17]), .Z(n36) );
  ND2 U46 ( .A(B[17]), .B(A[17]), .Z(n38) );
  AO6 U47 ( .A(n9), .B(n40), .C(n41), .Z(n37) );
  EO U48 ( .A(n40), .B(n43), .Z(SUM[16]) );
  NR2 U49 ( .A(n41), .B(n42), .Z(n43) );
  NR2 U50 ( .A(B[16]), .B(A[16]), .Z(n42) );
  AN2 U51 ( .A(B[16]), .B(A[16]), .Z(n41) );
  AO7 U52 ( .A(n44), .B(n45), .C(n46), .Z(n40) );
  EN U53 ( .A(n45), .B(n47), .Z(SUM[15]) );
  NR2 U54 ( .A(n10), .B(n44), .Z(n47) );
  NR2 U55 ( .A(B[15]), .B(A[15]), .Z(n44) );
  ND2 U56 ( .A(B[15]), .B(A[15]), .Z(n46) );
  AO6 U57 ( .A(n11), .B(n48), .C(n49), .Z(n45) );
  EO U58 ( .A(n48), .B(n51), .Z(SUM[14]) );
  NR2 U59 ( .A(n49), .B(n50), .Z(n51) );
  NR2 U60 ( .A(B[14]), .B(A[14]), .Z(n50) );
  AN2 U61 ( .A(B[14]), .B(A[14]), .Z(n49) );
  AO7 U62 ( .A(n52), .B(n53), .C(n54), .Z(n48) );
  EN U63 ( .A(n53), .B(n55), .Z(SUM[13]) );
  NR2 U64 ( .A(n12), .B(n52), .Z(n55) );
  NR2 U65 ( .A(B[13]), .B(A[13]), .Z(n52) );
  ND2 U66 ( .A(B[13]), .B(A[13]), .Z(n54) );
  AO6 U67 ( .A(n13), .B(n14), .C(n56), .Z(n53) );
  EO U68 ( .A(n14), .B(n58), .Z(SUM[12]) );
  NR2 U69 ( .A(n56), .B(n57), .Z(n58) );
  NR2 U70 ( .A(B[12]), .B(A[12]), .Z(n57) );
  AN2 U71 ( .A(B[12]), .B(A[12]), .Z(n56) );
  ND2 U72 ( .A(B[11]), .B(A[11]), .Z(n59) );
endmodule


module SinBlock_0_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [11:0] A;
  input [13:0] B;
  output [25:0] PRODUCT;
  input TC;
  wire   \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][13] ,
         \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] ,
         \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] ,
         \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][13] , \ab[8][12] , \ab[8][11] ,
         \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] , \ab[8][6] ,
         \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] ,
         \ab[8][0] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][13] ,
         \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] ,
         \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] ,
         \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][13] , \ab[3][12] , \ab[3][11] ,
         \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[0][13] , \ab[0][12] ,
         \ab[0][11] , \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] ,
         \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] ,
         \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] ,
         \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] ,
         \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] ,
         \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] ,
         \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][12] , \CARRYB[1][11] ,
         \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] ,
         \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[11][0] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][12] ,
         \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] ,
         \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] ,
         \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][12] ,
         \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] ,
         \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] ,
         \A2[17] , \A2[16] , \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] ,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8;

  SinBlock_0_DW01_add_1 FS_1 ( .A({1'b0, \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \SUMB[11][0] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[23] , 
        \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , 
        \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        PRODUCT[25:11], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8}) );
  FA1A S5_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\ab[10][13] ), .CO(
        \CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S3_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\ab[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S3_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\ab[8][13] ), .CO(
        \CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S3_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\ab[7][13] ), .CO(
        \CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S3_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\ab[6][13] ), .CO(
        \CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S3_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\ab[5][13] ), .CO(
        \CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S3_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\ab[4][13] ), .CO(
        \CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S3_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\ab[3][13] ), .CO(
        \CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S3_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\ab[2][13] ), .CO(
        \CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S3_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\ab[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S4_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(
        \CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S4_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), .CO(
        \CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S4_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(
        \CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S4_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(
        \CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S4_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(
        \CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S4_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(
        \CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S4_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(
        \CARRYB[11][0] ), .S(\SUMB[11][0] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S4_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(
        \CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S4_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(
        \CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(
        \CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  IVP U2 ( .A(A[0]), .Z(n10) );
  EO U3 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A1[12] ) );
  EO U4 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  EO U5 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A1[11] ) );
  EO U6 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A1[13] ) );
  EO U7 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A1[14] ) );
  EO U8 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A1[15] ) );
  EO U9 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A1[16] ) );
  EO U10 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A1[17] ) );
  EO U11 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A1[18] ) );
  EO U12 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A1[19] ) );
  EO U13 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A1[20] ) );
  EO U14 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A1[21] ) );
  EO U15 ( .A(\CARRYB[11][12] ), .B(\ab[11][13] ), .Z(\A1[22] ) );
  EO U16 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A1[10] ) );
  IVP U17 ( .A(A[1]), .Z(n11) );
  EO U18 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U19 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  IVP U20 ( .A(A[2]), .Z(n12) );
  EO U21 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U22 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U23 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  IVP U24 ( .A(A[3]), .Z(n13) );
  EO U25 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U26 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U27 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  IVP U28 ( .A(A[4]), .Z(n14) );
  EO U29 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U30 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  IVP U31 ( .A(A[5]), .Z(n15) );
  EO U32 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  IVP U33 ( .A(A[6]), .Z(n16) );
  IVP U34 ( .A(A[7]), .Z(n17) );
  IVP U35 ( .A(A[8]), .Z(n18) );
  IVP U36 ( .A(B[13]), .Z(n8) );
  IVP U37 ( .A(A[9]), .Z(n19) );
  IVP U38 ( .A(A[10]), .Z(n20) );
  IVP U39 ( .A(A[11]), .Z(n9) );
  IVP U40 ( .A(B[2]), .Z(n26) );
  IVP U41 ( .A(B[3]), .Z(n25) );
  IVP U42 ( .A(B[4]), .Z(n24) );
  IVP U43 ( .A(B[1]), .Z(n27) );
  IVP U44 ( .A(B[5]), .Z(n23) );
  IVP U45 ( .A(B[6]), .Z(n22) );
  IVP U46 ( .A(B[7]), .Z(n21) );
  IVP U47 ( .A(B[0]), .Z(n28) );
  IVP U48 ( .A(B[8]), .Z(n3) );
  IVP U49 ( .A(B[9]), .Z(n4) );
  IVP U50 ( .A(B[10]), .Z(n5) );
  IVP U51 ( .A(B[11]), .Z(n6) );
  IVP U52 ( .A(B[12]), .Z(n7) );
  AN2P U53 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A2[11] ) );
  AN2P U54 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A2[13] ) );
  AN2P U55 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A2[14] ) );
  AN2P U56 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A2[15] ) );
  AN2P U57 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A2[16] ) );
  AN2P U58 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A2[17] ) );
  AN2P U59 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A2[18] ) );
  AN2P U60 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A2[19] ) );
  AN2P U61 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A2[20] ) );
  AN2P U62 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A2[21] ) );
  AN2P U63 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A2[22] ) );
  AN2P U64 ( .A(\CARRYB[11][12] ), .B(\ab[11][13] ), .Z(\A2[23] ) );
  AN2P U65 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U66 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U67 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U68 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U69 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U70 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U71 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U72 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U73 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U74 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U75 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U76 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U77 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A2[12] ) );
  NR2 U79 ( .A(n19), .B(n4), .Z(\ab[9][9] ) );
  NR2 U80 ( .A(n19), .B(n3), .Z(\ab[9][8] ) );
  NR2 U81 ( .A(n19), .B(n21), .Z(\ab[9][7] ) );
  NR2 U82 ( .A(n19), .B(n22), .Z(\ab[9][6] ) );
  NR2 U83 ( .A(n19), .B(n23), .Z(\ab[9][5] ) );
  NR2 U84 ( .A(n19), .B(n24), .Z(\ab[9][4] ) );
  NR2 U85 ( .A(n19), .B(n25), .Z(\ab[9][3] ) );
  NR2 U86 ( .A(n19), .B(n26), .Z(\ab[9][2] ) );
  NR2 U87 ( .A(n19), .B(n27), .Z(\ab[9][1] ) );
  NR2 U88 ( .A(n19), .B(n8), .Z(\ab[9][13] ) );
  NR2 U89 ( .A(n19), .B(n7), .Z(\ab[9][12] ) );
  NR2 U90 ( .A(n19), .B(n6), .Z(\ab[9][11] ) );
  NR2 U91 ( .A(n19), .B(n5), .Z(\ab[9][10] ) );
  NR2 U92 ( .A(n19), .B(n28), .Z(\ab[9][0] ) );
  NR2 U93 ( .A(n4), .B(n18), .Z(\ab[8][9] ) );
  NR2 U94 ( .A(n3), .B(n18), .Z(\ab[8][8] ) );
  NR2 U95 ( .A(n21), .B(n18), .Z(\ab[8][7] ) );
  NR2 U96 ( .A(n22), .B(n18), .Z(\ab[8][6] ) );
  NR2 U97 ( .A(n23), .B(n18), .Z(\ab[8][5] ) );
  NR2 U98 ( .A(n24), .B(n18), .Z(\ab[8][4] ) );
  NR2 U99 ( .A(n25), .B(n18), .Z(\ab[8][3] ) );
  NR2 U100 ( .A(n26), .B(n18), .Z(\ab[8][2] ) );
  NR2 U101 ( .A(n27), .B(n18), .Z(\ab[8][1] ) );
  NR2 U102 ( .A(n8), .B(n18), .Z(\ab[8][13] ) );
  NR2 U103 ( .A(n7), .B(n18), .Z(\ab[8][12] ) );
  NR2 U104 ( .A(n6), .B(n18), .Z(\ab[8][11] ) );
  NR2 U105 ( .A(n5), .B(n18), .Z(\ab[8][10] ) );
  NR2 U106 ( .A(n28), .B(n18), .Z(\ab[8][0] ) );
  NR2 U107 ( .A(n4), .B(n17), .Z(\ab[7][9] ) );
  NR2 U108 ( .A(n3), .B(n17), .Z(\ab[7][8] ) );
  NR2 U109 ( .A(n21), .B(n17), .Z(\ab[7][7] ) );
  NR2 U110 ( .A(n22), .B(n17), .Z(\ab[7][6] ) );
  NR2 U111 ( .A(n23), .B(n17), .Z(\ab[7][5] ) );
  NR2 U112 ( .A(n24), .B(n17), .Z(\ab[7][4] ) );
  NR2 U113 ( .A(n25), .B(n17), .Z(\ab[7][3] ) );
  NR2 U114 ( .A(n26), .B(n17), .Z(\ab[7][2] ) );
  NR2 U115 ( .A(n27), .B(n17), .Z(\ab[7][1] ) );
  NR2 U116 ( .A(n8), .B(n17), .Z(\ab[7][13] ) );
  NR2 U117 ( .A(n7), .B(n17), .Z(\ab[7][12] ) );
  NR2 U118 ( .A(n6), .B(n17), .Z(\ab[7][11] ) );
  NR2 U119 ( .A(n5), .B(n17), .Z(\ab[7][10] ) );
  NR2 U120 ( .A(n28), .B(n17), .Z(\ab[7][0] ) );
  NR2 U121 ( .A(n4), .B(n16), .Z(\ab[6][9] ) );
  NR2 U122 ( .A(n3), .B(n16), .Z(\ab[6][8] ) );
  NR2 U123 ( .A(n21), .B(n16), .Z(\ab[6][7] ) );
  NR2 U124 ( .A(n22), .B(n16), .Z(\ab[6][6] ) );
  NR2 U125 ( .A(n23), .B(n16), .Z(\ab[6][5] ) );
  NR2 U126 ( .A(n24), .B(n16), .Z(\ab[6][4] ) );
  NR2 U127 ( .A(n25), .B(n16), .Z(\ab[6][3] ) );
  NR2 U128 ( .A(n26), .B(n16), .Z(\ab[6][2] ) );
  NR2 U129 ( .A(n27), .B(n16), .Z(\ab[6][1] ) );
  NR2 U130 ( .A(n8), .B(n16), .Z(\ab[6][13] ) );
  NR2 U131 ( .A(n7), .B(n16), .Z(\ab[6][12] ) );
  NR2 U132 ( .A(n6), .B(n16), .Z(\ab[6][11] ) );
  NR2 U133 ( .A(n5), .B(n16), .Z(\ab[6][10] ) );
  NR2 U134 ( .A(n28), .B(n16), .Z(\ab[6][0] ) );
  NR2 U135 ( .A(n4), .B(n15), .Z(\ab[5][9] ) );
  NR2 U136 ( .A(n3), .B(n15), .Z(\ab[5][8] ) );
  NR2 U137 ( .A(n21), .B(n15), .Z(\ab[5][7] ) );
  NR2 U138 ( .A(n22), .B(n15), .Z(\ab[5][6] ) );
  NR2 U139 ( .A(n23), .B(n15), .Z(\ab[5][5] ) );
  NR2 U140 ( .A(n24), .B(n15), .Z(\ab[5][4] ) );
  NR2 U141 ( .A(n25), .B(n15), .Z(\ab[5][3] ) );
  NR2 U142 ( .A(n26), .B(n15), .Z(\ab[5][2] ) );
  NR2 U143 ( .A(n27), .B(n15), .Z(\ab[5][1] ) );
  NR2 U144 ( .A(n8), .B(n15), .Z(\ab[5][13] ) );
  NR2 U145 ( .A(n7), .B(n15), .Z(\ab[5][12] ) );
  NR2 U146 ( .A(n6), .B(n15), .Z(\ab[5][11] ) );
  NR2 U147 ( .A(n5), .B(n15), .Z(\ab[5][10] ) );
  NR2 U148 ( .A(n28), .B(n15), .Z(\ab[5][0] ) );
  NR2 U149 ( .A(n4), .B(n14), .Z(\ab[4][9] ) );
  NR2 U150 ( .A(n3), .B(n14), .Z(\ab[4][8] ) );
  NR2 U151 ( .A(n21), .B(n14), .Z(\ab[4][7] ) );
  NR2 U152 ( .A(n22), .B(n14), .Z(\ab[4][6] ) );
  NR2 U153 ( .A(n23), .B(n14), .Z(\ab[4][5] ) );
  NR2 U154 ( .A(n24), .B(n14), .Z(\ab[4][4] ) );
  NR2 U155 ( .A(n25), .B(n14), .Z(\ab[4][3] ) );
  NR2 U156 ( .A(n26), .B(n14), .Z(\ab[4][2] ) );
  NR2 U157 ( .A(n27), .B(n14), .Z(\ab[4][1] ) );
  NR2 U158 ( .A(n8), .B(n14), .Z(\ab[4][13] ) );
  NR2 U159 ( .A(n7), .B(n14), .Z(\ab[4][12] ) );
  NR2 U160 ( .A(n6), .B(n14), .Z(\ab[4][11] ) );
  NR2 U161 ( .A(n5), .B(n14), .Z(\ab[4][10] ) );
  NR2 U162 ( .A(n28), .B(n14), .Z(\ab[4][0] ) );
  NR2 U163 ( .A(n4), .B(n13), .Z(\ab[3][9] ) );
  NR2 U164 ( .A(n3), .B(n13), .Z(\ab[3][8] ) );
  NR2 U165 ( .A(n21), .B(n13), .Z(\ab[3][7] ) );
  NR2 U166 ( .A(n22), .B(n13), .Z(\ab[3][6] ) );
  NR2 U167 ( .A(n23), .B(n13), .Z(\ab[3][5] ) );
  NR2 U168 ( .A(n24), .B(n13), .Z(\ab[3][4] ) );
  NR2 U169 ( .A(n25), .B(n13), .Z(\ab[3][3] ) );
  NR2 U170 ( .A(n26), .B(n13), .Z(\ab[3][2] ) );
  NR2 U171 ( .A(n27), .B(n13), .Z(\ab[3][1] ) );
  NR2 U172 ( .A(n8), .B(n13), .Z(\ab[3][13] ) );
  NR2 U173 ( .A(n7), .B(n13), .Z(\ab[3][12] ) );
  NR2 U174 ( .A(n6), .B(n13), .Z(\ab[3][11] ) );
  NR2 U175 ( .A(n5), .B(n13), .Z(\ab[3][10] ) );
  NR2 U176 ( .A(n28), .B(n13), .Z(\ab[3][0] ) );
  NR2 U177 ( .A(n4), .B(n12), .Z(\ab[2][9] ) );
  NR2 U178 ( .A(n3), .B(n12), .Z(\ab[2][8] ) );
  NR2 U179 ( .A(n21), .B(n12), .Z(\ab[2][7] ) );
  NR2 U180 ( .A(n22), .B(n12), .Z(\ab[2][6] ) );
  NR2 U181 ( .A(n23), .B(n12), .Z(\ab[2][5] ) );
  NR2 U182 ( .A(n24), .B(n12), .Z(\ab[2][4] ) );
  NR2 U183 ( .A(n25), .B(n12), .Z(\ab[2][3] ) );
  NR2 U184 ( .A(n26), .B(n12), .Z(\ab[2][2] ) );
  NR2 U185 ( .A(n27), .B(n12), .Z(\ab[2][1] ) );
  NR2 U186 ( .A(n8), .B(n12), .Z(\ab[2][13] ) );
  NR2 U187 ( .A(n7), .B(n12), .Z(\ab[2][12] ) );
  NR2 U188 ( .A(n6), .B(n12), .Z(\ab[2][11] ) );
  NR2 U189 ( .A(n5), .B(n12), .Z(\ab[2][10] ) );
  NR2 U190 ( .A(n28), .B(n12), .Z(\ab[2][0] ) );
  NR2 U191 ( .A(n4), .B(n11), .Z(\ab[1][9] ) );
  NR2 U192 ( .A(n3), .B(n11), .Z(\ab[1][8] ) );
  NR2 U193 ( .A(n21), .B(n11), .Z(\ab[1][7] ) );
  NR2 U194 ( .A(n22), .B(n11), .Z(\ab[1][6] ) );
  NR2 U195 ( .A(n23), .B(n11), .Z(\ab[1][5] ) );
  NR2 U196 ( .A(n24), .B(n11), .Z(\ab[1][4] ) );
  NR2 U197 ( .A(n25), .B(n11), .Z(\ab[1][3] ) );
  NR2 U198 ( .A(n26), .B(n11), .Z(\ab[1][2] ) );
  NR2 U199 ( .A(n8), .B(n11), .Z(\ab[1][13] ) );
  NR2 U200 ( .A(n7), .B(n11), .Z(\ab[1][12] ) );
  NR2 U201 ( .A(n6), .B(n11), .Z(\ab[1][11] ) );
  NR2 U202 ( .A(n5), .B(n11), .Z(\ab[1][10] ) );
  NR2 U203 ( .A(n4), .B(n9), .Z(\ab[11][9] ) );
  NR2 U204 ( .A(n3), .B(n9), .Z(\ab[11][8] ) );
  NR2 U205 ( .A(n21), .B(n9), .Z(\ab[11][7] ) );
  NR2 U206 ( .A(n22), .B(n9), .Z(\ab[11][6] ) );
  NR2 U207 ( .A(n23), .B(n9), .Z(\ab[11][5] ) );
  NR2 U208 ( .A(n24), .B(n9), .Z(\ab[11][4] ) );
  NR2 U209 ( .A(n25), .B(n9), .Z(\ab[11][3] ) );
  NR2 U210 ( .A(n26), .B(n9), .Z(\ab[11][2] ) );
  NR2 U211 ( .A(n27), .B(n9), .Z(\ab[11][1] ) );
  NR2 U212 ( .A(n8), .B(n9), .Z(\ab[11][13] ) );
  NR2 U213 ( .A(n7), .B(n9), .Z(\ab[11][12] ) );
  NR2 U214 ( .A(n6), .B(n9), .Z(\ab[11][11] ) );
  NR2 U215 ( .A(n5), .B(n9), .Z(\ab[11][10] ) );
  NR2 U216 ( .A(n28), .B(n9), .Z(\ab[11][0] ) );
  NR2 U217 ( .A(n4), .B(n20), .Z(\ab[10][9] ) );
  NR2 U218 ( .A(n3), .B(n20), .Z(\ab[10][8] ) );
  NR2 U219 ( .A(n21), .B(n20), .Z(\ab[10][7] ) );
  NR2 U220 ( .A(n22), .B(n20), .Z(\ab[10][6] ) );
  NR2 U221 ( .A(n23), .B(n20), .Z(\ab[10][5] ) );
  NR2 U222 ( .A(n24), .B(n20), .Z(\ab[10][4] ) );
  NR2 U223 ( .A(n25), .B(n20), .Z(\ab[10][3] ) );
  NR2 U224 ( .A(n26), .B(n20), .Z(\ab[10][2] ) );
  NR2 U225 ( .A(n27), .B(n20), .Z(\ab[10][1] ) );
  NR2 U226 ( .A(n8), .B(n20), .Z(\ab[10][13] ) );
  NR2 U227 ( .A(n7), .B(n20), .Z(\ab[10][12] ) );
  NR2 U228 ( .A(n6), .B(n20), .Z(\ab[10][11] ) );
  NR2 U229 ( .A(n5), .B(n20), .Z(\ab[10][10] ) );
  NR2 U230 ( .A(n28), .B(n20), .Z(\ab[10][0] ) );
  NR2 U231 ( .A(n4), .B(n10), .Z(\ab[0][9] ) );
  NR2 U232 ( .A(n3), .B(n10), .Z(\ab[0][8] ) );
  NR2 U233 ( .A(n21), .B(n10), .Z(\ab[0][7] ) );
  NR2 U234 ( .A(n22), .B(n10), .Z(\ab[0][6] ) );
  NR2 U235 ( .A(n23), .B(n10), .Z(\ab[0][5] ) );
  NR2 U236 ( .A(n24), .B(n10), .Z(\ab[0][4] ) );
  NR2 U237 ( .A(n25), .B(n10), .Z(\ab[0][3] ) );
  NR2 U238 ( .A(n26), .B(n10), .Z(\ab[0][2] ) );
  NR2 U239 ( .A(n8), .B(n10), .Z(\ab[0][13] ) );
  NR2 U240 ( .A(n7), .B(n10), .Z(\ab[0][12] ) );
  NR2 U241 ( .A(n6), .B(n10), .Z(\ab[0][11] ) );
  NR2 U242 ( .A(n5), .B(n10), .Z(\ab[0][10] ) );
  AN3 U243 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U244 ( .A(n11), .B(n27), .Z(\ab[1][1] ) );
endmodule


module SinBlock_0 ( clk, reset, func, x, sinValue );
  input [15:0] x;
  output [15:0] sinValue;
  input clk, reset, func;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         \Term2[18] , N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, sValue, N57, n35, \add_1242/carry[14] ,
         \add_1242/carry[13] , \add_1242/carry[12] , \add_1242/carry[11] ,
         \add_1242/carry[10] , \add_1242/carry[9] , \add_1242/carry[8] ,
         \add_1242/carry[7] , \add_1242/carry[6] , \add_1242/carry[5] ,
         \add_1242/carry[4] , \add_1242/carry[3] , \add_1242/carry[2] ,
         \add_1242/carry[1] , n1, n2, n3, n34, n36, n37, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544;
  wire   [25:11] Term1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10;

  SinBlock_0_DW02_mult_0 mult_1238 ( .A({n37, N9, N10, N11, N12, N13, N14, N15, 
        N16, N17, N18, N19}), .B({n542, x[12:0]}), .TC(1'b0), .PRODUCT({N34, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  FDS2L \Term1_reg[25]  ( .CR(1'b1), .D(N34), .LD(n544), .CP(clk), .Q(
        Term1[25]) );
  FDS2L \Term1_reg[24]  ( .CR(1'b1), .D(N33), .LD(n544), .CP(clk), .Q(
        Term1[24]) );
  FDS2L \Term1_reg[23]  ( .CR(1'b1), .D(N32), .LD(n544), .CP(clk), .Q(
        Term1[23]) );
  FDS2L \Term1_reg[22]  ( .CR(1'b1), .D(N31), .LD(n544), .CP(clk), .Q(
        Term1[22]) );
  FDS2L \Term1_reg[21]  ( .CR(1'b1), .D(N30), .LD(n544), .CP(clk), .Q(
        Term1[21]) );
  FDS2L \Term1_reg[20]  ( .CR(1'b1), .D(N29), .LD(n544), .CP(clk), .Q(
        Term1[20]) );
  FDS2L \Term1_reg[19]  ( .CR(1'b1), .D(N28), .LD(n544), .CP(clk), .Q(
        Term1[19]) );
  FDS2L \Term1_reg[18]  ( .CR(1'b1), .D(N27), .LD(n544), .CP(clk), .Q(
        Term1[18]) );
  FDS2L \Term1_reg[17]  ( .CR(1'b1), .D(N26), .LD(n544), .CP(clk), .Q(
        Term1[17]) );
  FDS2L \Term1_reg[16]  ( .CR(1'b1), .D(N25), .LD(n544), .CP(clk), .Q(
        Term1[16]) );
  FDS2L \Term1_reg[15]  ( .CR(1'b1), .D(N24), .LD(n544), .CP(clk), .Q(
        Term1[15]) );
  FDS2L \Term1_reg[14]  ( .CR(1'b1), .D(N23), .LD(n544), .CP(clk), .Q(
        Term1[14]) );
  FDS2L \Term1_reg[13]  ( .CR(1'b1), .D(N22), .LD(n544), .CP(clk), .Q(
        Term1[13]) );
  FDS2L \Term1_reg[12]  ( .CR(1'b1), .D(N21), .LD(n544), .CP(clk), .Q(
        Term1[12]) );
  FDS2L \Term1_reg[11]  ( .CR(1'b1), .D(N20), .LD(n544), .CP(clk), .Q(
        Term1[11]) );
  FDS2L \Term2_reg[18]  ( .CR(1'b1), .D(1'b1), .LD(n544), .CP(clk), .Q(
        \Term2[18] ) );
  FDS2L \sinValue_reg[14]  ( .CR(1'b1), .D(N50), .LD(n544), .CP(clk), .Q(
        sinValue[14]) );
  FDS2L \sinValue_reg[13]  ( .CR(1'b1), .D(N49), .LD(n544), .CP(clk), .Q(
        sinValue[13]) );
  FDS2L \sinValue_reg[12]  ( .CR(1'b1), .D(N48), .LD(n544), .CP(clk), .Q(
        sinValue[12]) );
  FDS2L \sinValue_reg[11]  ( .CR(1'b1), .D(N47), .LD(n544), .CP(clk), .Q(
        sinValue[11]) );
  FDS2L \sinValue_reg[10]  ( .CR(1'b1), .D(N46), .LD(n544), .CP(clk), .Q(
        sinValue[10]) );
  FDS2L \sinValue_reg[9]  ( .CR(1'b1), .D(N45), .LD(n544), .CP(clk), .Q(
        sinValue[9]) );
  FDS2L \sinValue_reg[8]  ( .CR(1'b1), .D(N44), .LD(n544), .CP(clk), .Q(
        sinValue[8]) );
  FDS2L \sinValue_reg[7]  ( .CR(1'b1), .D(N43), .LD(n544), .CP(clk), .Q(
        sinValue[7]) );
  FDS2L \sinValue_reg[6]  ( .CR(1'b1), .D(N42), .LD(n544), .CP(clk), .Q(
        sinValue[6]) );
  FDS2L \sinValue_reg[5]  ( .CR(1'b1), .D(N41), .LD(n544), .CP(clk), .Q(
        sinValue[5]) );
  FDS2L \sinValue_reg[4]  ( .CR(1'b1), .D(N40), .LD(n544), .CP(clk), .Q(
        sinValue[4]) );
  FDS2L \sinValue_reg[3]  ( .CR(1'b1), .D(N39), .LD(n544), .CP(clk), .Q(
        sinValue[3]) );
  FDS2L \sinValue_reg[2]  ( .CR(1'b1), .D(N38), .LD(n544), .CP(clk), .Q(
        sinValue[2]) );
  FDS2L \sinValue_reg[1]  ( .CR(1'b1), .D(N37), .LD(n544), .CP(clk), .Q(
        sinValue[1]) );
  FDS2L \sinValue_reg[15]  ( .CR(1'b1), .D(sValue), .LD(n544), .CP(clk), .Q(
        sinValue[15]) );
  FDS2L sValue_reg ( .CR(1'b1), .D(N57), .LD(n544), .CP(clk), .Q(sValue) );
  FDS2L \sinValue_reg[0]  ( .CR(1'b1), .D(N36), .LD(n544), .CP(clk), .Q(
        sinValue[0]) );
  AN2P U3 ( .A(n339), .B(n338), .Z(n1) );
  AN2P U4 ( .A(n300), .B(n299), .Z(n2) );
  AN2P U5 ( .A(n243), .B(n242), .Z(n3) );
  AN2P U6 ( .A(n258), .B(n257), .Z(n34) );
  AN2P U7 ( .A(n324), .B(n323), .Z(n36) );
  AN2P U8 ( .A(n425), .B(n44), .Z(n37) );
  NR2 U12 ( .A(n463), .B(n503), .Z(n186) );
  NR2 U13 ( .A(n500), .B(n465), .Z(n229) );
  NR2 U14 ( .A(n532), .B(n500), .Z(n231) );
  EO U15 ( .A(n527), .B(n495), .Z(n163) );
  ND2 U16 ( .A(n529), .B(n332), .Z(n179) );
  ND2 U17 ( .A(n496), .B(n461), .Z(n332) );
  ND2 U18 ( .A(n502), .B(n203), .Z(n150) );
  ND2 U19 ( .A(n534), .B(n462), .Z(n203) );
  ND2 U20 ( .A(n334), .B(n333), .Z(n162) );
  ND2 U21 ( .A(n528), .B(n460), .Z(n333) );
  EN U22 ( .A(n527), .B(n496), .Z(n334) );
  ND2 U23 ( .A(n468), .B(n530), .Z(n289) );
  AN2P U24 ( .A(n530), .B(n468), .Z(n41) );
  MUX21L U25 ( .A(n530), .B(n503), .S(n464), .Z(n148) );
  MUX21L U26 ( .A(n500), .B(n465), .S(n532), .Z(n153) );
  MUX21L U27 ( .A(n530), .B(n288), .S(n497), .Z(n290) );
  NR2 U28 ( .A(n529), .B(n468), .Z(n288) );
  ND2 U29 ( .A(n266), .B(n265), .Z(n144) );
  ND2 U30 ( .A(n466), .B(n498), .Z(n265) );
  MUX21L U31 ( .A(n264), .B(n499), .S(n531), .Z(n266) );
  NR2 U32 ( .A(n499), .B(n466), .Z(n264) );
  AO4 U33 ( .A(n496), .B(n462), .C(n528), .D(n461), .Z(n146) );
  AO4 U34 ( .A(n529), .B(n469), .C(n529), .D(n497), .Z(n176) );
  AO7 U35 ( .A(n528), .B(n496), .C(n470), .Z(n161) );
  AO7 U36 ( .A(n532), .B(n500), .C(n465), .Z(n141) );
  ND2 U37 ( .A(n497), .B(n302), .Z(n160) );
  ND2 U38 ( .A(n529), .B(n469), .Z(n302) );
  ND2 U39 ( .A(n225), .B(n224), .Z(n139) );
  ND2 U40 ( .A(n461), .B(n501), .Z(n224) );
  MUX21L U41 ( .A(n223), .B(n501), .S(n533), .Z(n225) );
  NR2 U42 ( .A(n501), .B(n462), .Z(n223) );
  EO U43 ( .A(n495), .B(n465), .Z(n245) );
  EN U44 ( .A(n527), .B(n498), .Z(n129) );
  EN U45 ( .A(n527), .B(n469), .Z(n131) );
  NR2 U46 ( .A(n530), .B(n467), .Z(n285) );
  ND2 U47 ( .A(n228), .B(n227), .Z(n112) );
  ND2 U48 ( .A(n461), .B(n501), .Z(n227) );
  MUX21L U49 ( .A(n226), .B(n501), .S(n533), .Z(n228) );
  NR2 U50 ( .A(n501), .B(n461), .Z(n226) );
  EO U51 ( .A(n526), .B(n501), .Z(n111) );
  ND2 U52 ( .A(n503), .B(n464), .Z(n108) );
  NR2 U53 ( .A(n531), .B(n467), .Z(n273) );
  AO4 U54 ( .A(n502), .B(n463), .C(n534), .D(n462), .Z(n92) );
  EN U55 ( .A(n527), .B(n499), .Z(n97) );
  EN U56 ( .A(n527), .B(n500), .Z(n96) );
  ND2 U57 ( .A(n307), .B(n306), .Z(n102) );
  EN U58 ( .A(n527), .B(n469), .Z(n307) );
  ND2 U59 ( .A(n496), .B(n469), .Z(n306) );
  ND2 U60 ( .A(n503), .B(n464), .Z(n90) );
  EO U61 ( .A(n527), .B(n470), .Z(n103) );
  EO U62 ( .A(n527), .B(n470), .Z(n104) );
  EO U63 ( .A(n527), .B(n461), .Z(n105) );
  AO4 U64 ( .A(n501), .B(n462), .C(n533), .D(n462), .Z(n78) );
  EO U65 ( .A(n495), .B(n466), .Z(n81) );
  ND2 U66 ( .A(n533), .B(n502), .Z(n209) );
  ND2 U67 ( .A(n280), .B(n279), .Z(n68) );
  EN U68 ( .A(n495), .B(n467), .Z(n280) );
  EN U69 ( .A(n527), .B(n467), .Z(n279) );
  ND2 U70 ( .A(n500), .B(n466), .Z(n254) );
  ND2 U71 ( .A(n532), .B(n465), .Z(n255) );
  AO4 U72 ( .A(n498), .B(n468), .C(n530), .D(n468), .Z(n69) );
  AO7 U73 ( .A(n529), .B(n497), .C(n470), .Z(n72) );
  ND2 U74 ( .A(n351), .B(n350), .Z(n74) );
  ND2 U75 ( .A(n503), .B(n460), .Z(n350) );
  ND2 U76 ( .A(n530), .B(n460), .Z(n351) );
  ND2 U77 ( .A(n309), .B(n308), .Z(n70) );
  ND2 U78 ( .A(n529), .B(n469), .Z(n309) );
  ND2 U79 ( .A(n497), .B(n469), .Z(n308) );
  AN2P U80 ( .A(n498), .B(n467), .Z(n42) );
  MUX21L U81 ( .A(n461), .B(n331), .S(n497), .Z(n73) );
  ND2 U82 ( .A(n527), .B(n461), .Z(n331) );
  AN3 U83 ( .A(n495), .B(n460), .C(n526), .Z(n59) );
  ND2 U84 ( .A(n529), .B(n470), .Z(n324) );
  ND2 U85 ( .A(n498), .B(n470), .Z(n323) );
  AO4 U86 ( .A(n497), .B(n468), .C(n530), .D(n468), .Z(n51) );
  ND2 U87 ( .A(n499), .B(n466), .Z(n260) );
  AN2P U88 ( .A(n503), .B(n464), .Z(n43) );
  IVP U89 ( .A(n442), .Z(n466) );
  IVP U90 ( .A(n442), .Z(n463) );
  IVP U91 ( .A(n442), .Z(n467) );
  ND2 U92 ( .A(n259), .B(n518), .Z(n172) );
  EO U93 ( .A(n495), .B(n466), .Z(n259) );
  ND2 U94 ( .A(n190), .B(n189), .Z(n149) );
  MUX21L U95 ( .A(n187), .B(n188), .S(n503), .Z(n190) );
  ND2 U96 ( .A(n186), .B(n523), .Z(n189) );
  NR2 U97 ( .A(n534), .B(n450), .Z(n188) );
  ND2 U98 ( .A(n268), .B(n267), .Z(n158) );
  ND2 U99 ( .A(n467), .B(n516), .Z(n267) );
  EN U100 ( .A(n495), .B(n467), .Z(n268) );
  IVP U101 ( .A(n441), .Z(n460) );
  IVP U102 ( .A(n442), .Z(n465) );
  IVP U103 ( .A(n477), .Z(n500) );
  IVP U104 ( .A(n510), .Z(n531) );
  IVP U105 ( .A(n476), .Z(n497) );
  IVP U106 ( .A(n510), .Z(n533) );
  IVP U107 ( .A(n477), .Z(n502) );
  IVP U108 ( .A(n510), .Z(n532) );
  IVP U109 ( .A(n442), .Z(n464) );
  IVP U110 ( .A(n477), .Z(n503) );
  IVP U111 ( .A(n476), .Z(n496) );
  IVP U112 ( .A(n509), .Z(n527) );
  IVP U113 ( .A(n510), .Z(n530) );
  IVP U114 ( .A(n476), .Z(n495) );
  IVP U115 ( .A(n510), .Z(n534) );
  IVP U116 ( .A(n442), .Z(n468) );
  AO7 U117 ( .A(n499), .B(n524), .C(n465), .Z(n165) );
  ND3 U118 ( .A(n248), .B(n247), .C(n246), .Z(n171) );
  ND2 U119 ( .A(n452), .B(n488), .Z(n247) );
  ND2 U120 ( .A(n532), .B(n488), .Z(n248) );
  ND2 U121 ( .A(n532), .B(n452), .Z(n246) );
  ND2 U122 ( .A(n233), .B(n232), .Z(n170) );
  MUX21L U123 ( .A(n230), .B(n231), .S(n464), .Z(n233) );
  ND2 U124 ( .A(n229), .B(n533), .Z(n232) );
  NR2 U125 ( .A(n533), .B(n489), .Z(n230) );
  ND2 U126 ( .A(n201), .B(n200), .Z(n167) );
  ND2 U127 ( .A(n502), .B(n522), .Z(n200) );
  MUX21L U128 ( .A(n522), .B(n199), .S(n463), .Z(n201) );
  NR2 U129 ( .A(n502), .B(n522), .Z(n199) );
  ND2 U130 ( .A(n212), .B(n211), .Z(n168) );
  ND2 U131 ( .A(n502), .B(n520), .Z(n211) );
  MUX21L U132 ( .A(n521), .B(n210), .S(n463), .Z(n212) );
  NR2 U133 ( .A(n502), .B(n520), .Z(n210) );
  ND2 U149 ( .A(n314), .B(n313), .Z(n177) );
  ND2 U150 ( .A(n310), .B(n512), .Z(n313) );
  MUX21L U151 ( .A(n311), .B(n312), .S(n496), .Z(n314) );
  NR2 U152 ( .A(n470), .B(n497), .Z(n310) );
  ND2 U153 ( .A(n250), .B(n249), .Z(n154) );
  ND2 U154 ( .A(n453), .B(n488), .Z(n249) );
  EN U155 ( .A(n527), .B(n500), .Z(n250) );
  ND2 U156 ( .A(n444), .B(n511), .Z(n338) );
  MUX21L U157 ( .A(n478), .B(n337), .S(n461), .Z(n339) );
  MUX21L U158 ( .A(n194), .B(n450), .S(n534), .Z(n166) );
  ND2 U159 ( .A(n450), .B(n492), .Z(n194) );
  MUX21L U160 ( .A(n282), .B(n281), .S(n498), .Z(n175) );
  ND2 U161 ( .A(n531), .B(n457), .Z(n282) );
  ND2 U162 ( .A(n530), .B(n467), .Z(n281) );
  MUX21L U178 ( .A(n214), .B(n213), .S(n502), .Z(n151) );
  ND2 U179 ( .A(n448), .B(n520), .Z(n213) );
  ND2 U180 ( .A(n533), .B(n448), .Z(n214) );
  MUX21L U181 ( .A(n486), .B(n517), .S(n466), .Z(n157) );
  MUX21L U182 ( .A(n514), .B(n484), .S(n468), .Z(n159) );
  IVP U183 ( .A(n509), .Z(n529) );
  IVP U184 ( .A(n509), .Z(n528) );
  IVP U185 ( .A(n443), .Z(n470) );
  IVP U186 ( .A(n441), .Z(n462) );
  IVP U187 ( .A(n476), .Z(n498) );
  IVP U188 ( .A(n476), .Z(n499) );
  AO7 U189 ( .A(n533), .B(n490), .C(n445), .Z(n169) );
  AO7 U190 ( .A(n499), .B(n517), .C(n455), .Z(n155) );
  NR2 U191 ( .A(n529), .B(n459), .Z(n312) );
  NR2 U192 ( .A(n532), .B(n489), .Z(n236) );
  ND2 U193 ( .A(n531), .B(n456), .Z(n174) );
  ND2 U194 ( .A(n238), .B(n237), .Z(n140) );
  ND2 U195 ( .A(n234), .B(n519), .Z(n237) );
  MUX21L U196 ( .A(n235), .B(n236), .S(n465), .Z(n238) );
  NR2 U197 ( .A(n465), .B(n500), .Z(n234) );
  ND2 U198 ( .A(n197), .B(n196), .Z(n136) );
  ND2 U199 ( .A(n463), .B(n492), .Z(n196) );
  MUX21L U200 ( .A(n195), .B(n534), .S(n463), .Z(n197) );
  NR2 U201 ( .A(n534), .B(n492), .Z(n195) );
  ND2 U202 ( .A(n183), .B(n182), .Z(n135) );
  ND2 U203 ( .A(n464), .B(n494), .Z(n182) );
  MUX21L U204 ( .A(n494), .B(n181), .S(n534), .Z(n183) );
  NR2 U205 ( .A(n464), .B(n494), .Z(n181) );
  ND2 U206 ( .A(n218), .B(n447), .Z(n138) );
  ND2 U207 ( .A(n533), .B(n501), .Z(n218) );
  MUX21L U208 ( .A(n490), .B(n519), .S(n462), .Z(n152) );
  MUX21L U209 ( .A(n205), .B(n204), .S(n534), .Z(n137) );
  ND2 U210 ( .A(n462), .B(n491), .Z(n205) );
  ND2 U211 ( .A(n502), .B(n462), .Z(n204) );
  IVP U212 ( .A(n441), .Z(n461) );
  IVP U213 ( .A(n443), .Z(n469) );
  IVP U214 ( .A(n477), .Z(n501) );
  ND2 U215 ( .A(n469), .B(n484), .Z(n300) );
  ND2 U216 ( .A(n469), .B(n513), .Z(n299) );
  ND2 U217 ( .A(n463), .B(n493), .Z(n192) );
  MUX21L U218 ( .A(n493), .B(n191), .S(n534), .Z(n193) );
  NR2 U219 ( .A(n463), .B(n493), .Z(n191) );
  ND2 U220 ( .A(n185), .B(n184), .Z(n122) );
  ND2 U221 ( .A(n534), .B(n451), .Z(n184) );
  EN U222 ( .A(n495), .B(n464), .Z(n185) );
  MUX21L U223 ( .A(n463), .B(n202), .S(n534), .Z(n124) );
  ND2 U224 ( .A(n463), .B(n491), .Z(n202) );
  ND2 U225 ( .A(n501), .B(n446), .Z(n222) );
  ND2 U226 ( .A(n341), .B(n340), .Z(n133) );
  ND2 U227 ( .A(n496), .B(n444), .Z(n340) );
  EO U228 ( .A(n526), .B(n460), .Z(n341) );
  MUX21L U229 ( .A(n283), .B(n498), .S(n467), .Z(n130) );
  ND2 U230 ( .A(n497), .B(n515), .Z(n283) );
  AO7 U231 ( .A(n531), .B(n498), .C(n456), .Z(n128) );
  ND2 U232 ( .A(n455), .B(n487), .Z(n142) );
  ND2 U233 ( .A(n452), .B(n518), .Z(n244) );
  ND2 U234 ( .A(n287), .B(n286), .Z(n117) );
  MUX21L U235 ( .A(n284), .B(n515), .S(n497), .Z(n286) );
  AO6 U236 ( .A(n499), .B(n457), .C(n285), .Z(n287) );
  ND2 U237 ( .A(n305), .B(n304), .Z(n118) );
  ND2 U238 ( .A(n483), .B(n513), .Z(n304) );
  MUX21L U239 ( .A(n483), .B(n303), .S(n469), .Z(n305) );
  ND2 U240 ( .A(n271), .B(n270), .Z(n116) );
  ND2 U241 ( .A(n531), .B(n456), .Z(n270) );
  MUX21L U242 ( .A(n486), .B(n269), .S(n467), .Z(n271) );
  NR2 U243 ( .A(n531), .B(n486), .Z(n269) );
  ND2 U244 ( .A(n241), .B(n240), .Z(n113) );
  ND2 U245 ( .A(n532), .B(n489), .Z(n240) );
  MUX21L U246 ( .A(n239), .B(n451), .S(n532), .Z(n241) );
  ND2 U247 ( .A(n208), .B(n207), .Z(n110) );
  MUX21L U248 ( .A(n206), .B(n521), .S(n502), .Z(n208) );
  ND2 U249 ( .A(n463), .B(n502), .Z(n207) );
  NR2 U250 ( .A(n462), .B(n521), .Z(n206) );
  MUX21L U251 ( .A(n325), .B(n527), .S(n461), .Z(n132) );
  ND2 U252 ( .A(n529), .B(n480), .Z(n325) );
  AO7 U253 ( .A(n499), .B(n466), .C(n517), .Z(n115) );
  ND2 U254 ( .A(n344), .B(n343), .Z(n120) );
  ND2 U255 ( .A(n528), .B(n495), .Z(n343) );
  MUX21L U256 ( .A(n342), .B(n444), .S(n495), .Z(n344) );
  NR2 U257 ( .A(n528), .B(n443), .Z(n342) );
  MUX21L U258 ( .A(n198), .B(n449), .S(n502), .Z(n109) );
  ND2 U259 ( .A(n449), .B(n523), .Z(n198) );
  ND2 U260 ( .A(n275), .B(n274), .Z(n100) );
  MUX21L U261 ( .A(n272), .B(n516), .S(n498), .Z(n274) );
  AO6 U262 ( .A(n498), .B(n457), .C(n273), .Z(n275) );
  ND2 U263 ( .A(n327), .B(n326), .Z(n119) );
  ND2 U264 ( .A(n480), .B(n512), .Z(n327) );
  ND2 U265 ( .A(n461), .B(n480), .Z(n326) );
  AO7 U266 ( .A(n532), .B(n451), .C(n500), .Z(n95) );
  NR2 U267 ( .A(n468), .B(n485), .Z(n291) );
  NR2 U268 ( .A(n497), .B(n514), .Z(n292) );
  NR2 U269 ( .A(n528), .B(n477), .Z(n346) );
  ND2 U270 ( .A(n295), .B(n294), .Z(n101) );
  NR2 U271 ( .A(n293), .B(n292), .Z(n295) );
  MUX21L U272 ( .A(n291), .B(n468), .S(n530), .Z(n294) );
  NR2 U273 ( .A(n498), .B(n458), .Z(n293) );
  ND2 U274 ( .A(n263), .B(n262), .Z(n99) );
  ND2 U275 ( .A(n531), .B(n487), .Z(n263) );
  ND2 U276 ( .A(n466), .B(n487), .Z(n262) );
  ND2 U277 ( .A(n349), .B(n348), .Z(n106) );
  NR2 U278 ( .A(n347), .B(n346), .Z(n349) );
  MUX21L U279 ( .A(n345), .B(n460), .S(n496), .Z(n348) );
  NR2 U280 ( .A(n527), .B(n443), .Z(n347) );
  ND2 U281 ( .A(n217), .B(n216), .Z(n93) );
  ND2 U282 ( .A(n447), .B(n519), .Z(n216) );
  MUX21L U283 ( .A(n490), .B(n215), .S(n462), .Z(n217) );
  ND2 U284 ( .A(n221), .B(n220), .Z(n94) );
  ND2 U285 ( .A(n501), .B(n446), .Z(n220) );
  ND2 U286 ( .A(n533), .B(n446), .Z(n221) );
  NR2 U287 ( .A(n460), .B(n511), .Z(n345) );
  NR2 U288 ( .A(n499), .B(n454), .Z(n256) );
  ND2 U289 ( .A(n465), .B(n518), .Z(n242) );
  EN U290 ( .A(n495), .B(n465), .Z(n243) );
  ND2 U291 ( .A(n499), .B(n454), .Z(n257) );
  MUX21L U292 ( .A(n256), .B(n455), .S(n531), .Z(n258) );
  ND2 U293 ( .A(n253), .B(n252), .Z(n79) );
  ND2 U294 ( .A(n500), .B(n453), .Z(n252) );
  MUX21L U295 ( .A(n251), .B(n454), .S(n532), .Z(n253) );
  NR2 U296 ( .A(n500), .B(n453), .Z(n251) );
  ND3 U297 ( .A(n278), .B(n277), .C(n276), .Z(n82) );
  ND2 U298 ( .A(n485), .B(n515), .Z(n277) );
  ND2 U299 ( .A(n467), .B(n516), .Z(n278) );
  ND2 U300 ( .A(n467), .B(n485), .Z(n276) );
  ND2 U301 ( .A(n297), .B(n296), .Z(n83) );
  ND2 U302 ( .A(n458), .B(n514), .Z(n296) );
  EO U303 ( .A(n495), .B(n469), .Z(n297) );
  ND2 U304 ( .A(n322), .B(n321), .Z(n86) );
  ND2 U305 ( .A(n530), .B(n496), .Z(n321) );
  MUX21L U306 ( .A(n320), .B(n459), .S(n496), .Z(n322) );
  NR2 U307 ( .A(n528), .B(n459), .Z(n320) );
  ND3 U308 ( .A(n491), .B(n523), .C(n449), .Z(n91) );
  ND2 U309 ( .A(n317), .B(n316), .Z(n85) );
  ND2 U310 ( .A(n528), .B(n482), .Z(n316) );
  MUX21L U311 ( .A(n482), .B(n315), .S(n470), .Z(n317) );
  NR2 U312 ( .A(n529), .B(n481), .Z(n315) );
  ND2 U313 ( .A(n330), .B(n329), .Z(n87) );
  ND2 U314 ( .A(n528), .B(n479), .Z(n329) );
  MUX21L U315 ( .A(n479), .B(n328), .S(n462), .Z(n330) );
  NR2 U316 ( .A(n528), .B(n479), .Z(n328) );
  MUX21L U317 ( .A(n336), .B(n335), .S(n461), .Z(n88) );
  ND2 U318 ( .A(n478), .B(n511), .Z(n335) );
  ND2 U319 ( .A(n528), .B(n496), .Z(n336) );
  MUX21L U320 ( .A(n483), .B(n301), .S(n469), .Z(n84) );
  ND2 U321 ( .A(n484), .B(n513), .Z(n301) );
  ND2 U322 ( .A(n219), .B(n447), .Z(n64) );
  ND2 U323 ( .A(n533), .B(n501), .Z(n219) );
  ND2 U324 ( .A(n319), .B(n318), .Z(n71) );
  ND2 U325 ( .A(n470), .B(n512), .Z(n318) );
  EN U326 ( .A(n495), .B(n470), .Z(n319) );
  MUX21L U327 ( .A(n49), .B(n48), .S(n432), .Z(n409) );
  ND2 U328 ( .A(n503), .B(n464), .Z(n48) );
  ND2 U329 ( .A(n261), .B(n260), .Z(n49) );
  ND2 U330 ( .A(n531), .B(n466), .Z(n261) );
  ND2 U331 ( .A(n431), .B(n43), .Z(n353) );
  MUX21L U332 ( .A(n417), .B(n416), .S(n435), .Z(n419) );
  AN3 U333 ( .A(n431), .B(n145), .C(n438), .Z(n417) );
  ND2 U334 ( .A(n290), .B(n289), .Z(n145) );
  MUX21L U335 ( .A(n413), .B(n412), .S(n432), .Z(n421) );
  NR3 U336 ( .A(n438), .B(n2), .C(n434), .Z(n412) );
  NR2 U337 ( .A(n438), .B(n1), .Z(n413) );
  MUX21L U338 ( .A(n415), .B(n414), .S(n438), .Z(n420) );
  NR2 U339 ( .A(n432), .B(n423), .Z(n414) );
  IVP U340 ( .A(n146), .Z(n423) );
  IVP U341 ( .A(n428), .Z(n431) );
  IVP U342 ( .A(n427), .Z(n430) );
  MUX21L U343 ( .A(n367), .B(n366), .S(n431), .Z(n370) );
  AN3 U344 ( .A(n125), .B(n434), .C(n438), .Z(n367) );
  AN3 U345 ( .A(n122), .B(n434), .C(n438), .Z(n366) );
  MUX21L U346 ( .A(n222), .B(n445), .S(n533), .Z(n125) );
  IVP U347 ( .A(n429), .Z(n432) );
  ND2 U348 ( .A(n434), .B(n426), .Z(n418) );
  AO2 U349 ( .A(n398), .B(n435), .C(n397), .D(n435), .Z(n406) );
  NR2 U350 ( .A(n439), .B(n427), .Z(n397) );
  NR2 U351 ( .A(n439), .B(n3), .Z(n398) );
  MUX21L U352 ( .A(n399), .B(n400), .S(n432), .Z(n408) );
  NR2 U353 ( .A(n439), .B(n422), .Z(n400) );
  NR3 U354 ( .A(n439), .B(n34), .C(n435), .Z(n399) );
  IVP U355 ( .A(n78), .Z(n422) );
  MUX21L U356 ( .A(n404), .B(n403), .S(n432), .Z(n405) );
  AN3 U357 ( .A(n438), .B(n460), .C(n434), .Z(n404) );
  ND2 U358 ( .A(n503), .B(n464), .Z(n76) );
  MUX21L U359 ( .A(n358), .B(n359), .S(n435), .Z(n361) );
  NR2 U360 ( .A(n439), .B(n429), .Z(n359) );
  ND2 U361 ( .A(n255), .B(n254), .Z(n65) );
  MUX21L U362 ( .A(n354), .B(n355), .S(n435), .Z(n363) );
  NR2 U363 ( .A(n439), .B(n59), .Z(n355) );
  MUX21L U364 ( .A(n356), .B(n357), .S(n435), .Z(n362) );
  ND2 U365 ( .A(n503), .B(n464), .Z(n63) );
  MUX21L U366 ( .A(n389), .B(n390), .S(n435), .Z(n395) );
  AN3 U367 ( .A(n61), .B(n426), .C(n438), .Z(n389) );
  ND2 U368 ( .A(n445), .B(n478), .Z(n61) );
  MUX21L U369 ( .A(n387), .B(n388), .S(n435), .Z(n396) );
  NR2 U370 ( .A(n439), .B(n427), .Z(n387) );
  AN3 U371 ( .A(n495), .B(n460), .C(n527), .Z(n57) );
  MUX21L U372 ( .A(n391), .B(n392), .S(n435), .Z(n394) );
  AO4 U373 ( .A(n498), .B(n468), .C(n530), .D(n468), .Z(n58) );
  MUX21L U374 ( .A(n373), .B(n53), .S(n431), .Z(n378) );
  ND2 U375 ( .A(n503), .B(n464), .Z(n53) );
  MUX21L U376 ( .A(n381), .B(n382), .S(n435), .Z(n383) );
  NR2 U377 ( .A(n432), .B(n36), .Z(n382) );
  EN U378 ( .A(n438), .B(n432), .Z(n410) );
  EN U379 ( .A(n434), .B(n432), .Z(n411) );
  ND2 U380 ( .A(n46), .B(n439), .Z(n386) );
  ND2 U381 ( .A(n298), .B(n458), .Z(n46) );
  ND2 U382 ( .A(n529), .B(n497), .Z(n298) );
  MUX21L U383 ( .A(n379), .B(n380), .S(n432), .Z(n384) );
  NR2 U384 ( .A(n439), .B(n435), .Z(n380) );
  ND2 U385 ( .A(n435), .B(n431), .Z(n385) );
  ND2 U386 ( .A(n440), .B(n435), .Z(n352) );
  NR2 U387 ( .A(n470), .B(n481), .Z(n178) );
  IVP U388 ( .A(n471), .Z(n472) );
  ND4 U389 ( .A(n421), .B(n420), .C(n419), .D(n418), .Z(n147) );
  IVP U390 ( .A(n504), .Z(n505) );
  ND3 U391 ( .A(n372), .B(n371), .C(n370), .Z(n127) );
  IVP U392 ( .A(n444), .Z(n474) );
  IVP U393 ( .A(n448), .Z(n475) );
  IVP U394 ( .A(n478), .Z(n507) );
  IVP U395 ( .A(n471), .Z(n473) );
  MUX21L U396 ( .A(n368), .B(n369), .S(n431), .Z(n371) );
  NR3 U397 ( .A(n439), .B(n534), .C(n435), .Z(n369) );
  AN3 U398 ( .A(n126), .B(n437), .C(n434), .Z(n368) );
  ND2 U399 ( .A(n245), .B(n244), .Z(n126) );
  MUX21L U400 ( .A(n364), .B(n365), .S(n435), .Z(n372) );
  AN3 U401 ( .A(n123), .B(n437), .C(n430), .Z(n365) );
  AN3 U402 ( .A(n124), .B(n430), .C(n438), .Z(n364) );
  ND2 U403 ( .A(n193), .B(n192), .Z(n123) );
  IVP U404 ( .A(n433), .Z(n436) );
  IVP U405 ( .A(n433), .Z(n434) );
  IVP U406 ( .A(n504), .Z(n506) );
  IVP U407 ( .A(n479), .Z(n508) );
  IVP U408 ( .A(n433), .Z(n435) );
  IVP U409 ( .A(n437), .Z(n440) );
  IVP U410 ( .A(n437), .Z(n438) );
  IVP U411 ( .A(n437), .Z(n439) );
  ND4 U412 ( .A(n408), .B(n407), .C(n406), .D(n405), .Z(n80) );
  MUX21L U413 ( .A(n402), .B(n401), .S(n432), .Z(n407) );
  AN3 U414 ( .A(n77), .B(n433), .C(n438), .Z(n401) );
  AN3 U415 ( .A(n79), .B(n433), .C(n438), .Z(n402) );
  ND2 U416 ( .A(n209), .B(n448), .Z(n77) );
  ND4 U417 ( .A(n363), .B(n362), .C(n361), .D(n360), .Z(n67) );
  ND4 U418 ( .A(n66), .B(n428), .C(n433), .D(n437), .Z(n360) );
  AO7 U419 ( .A(n531), .B(n499), .C(n466), .Z(n66) );
  ND4 U420 ( .A(n396), .B(n395), .C(n394), .D(n393), .Z(n62) );
  ND4 U421 ( .A(n378), .B(n377), .C(n376), .D(n375), .Z(n56) );
  ND3 U422 ( .A(n55), .B(n437), .C(n433), .Z(n375) );
  AO7 U423 ( .A(n531), .B(n499), .C(n466), .Z(n55) );
  MUX21L U424 ( .A(n374), .B(n437), .S(n432), .Z(n377) );
  AN3 U425 ( .A(n495), .B(n460), .C(n526), .Z(n54) );
  ND4 U426 ( .A(n60), .B(n435), .C(n428), .D(n437), .Z(n393) );
  AO7 U427 ( .A(n528), .B(n496), .C(n470), .Z(n60) );
  ND3 U428 ( .A(n411), .B(n410), .C(n409), .Z(n50) );
  ND2 U429 ( .A(n384), .B(n383), .Z(n52) );
  ND2 U430 ( .A(n431), .B(n433), .Z(n376) );
  AO7 U431 ( .A(n429), .B(n386), .C(n385), .Z(n47) );
  ND4 U432 ( .A(n439), .B(n435), .C(n432), .D(n43), .Z(n45) );
  NR2 U433 ( .A(n353), .B(n352), .Z(n44) );
  IVP U434 ( .A(n424), .Z(n425) );
  EN U435 ( .A(n35), .B(x[15]), .Z(N57) );
  ND2 U436 ( .A(x[14]), .B(func), .Z(n35) );
  IVP U437 ( .A(reset), .Z(n544) );
  MUX21H U438 ( .A(n47), .B(n45), .S(n425), .Z(N9) );
  MUX21H U439 ( .A(n52), .B(n50), .S(n425), .Z(N10) );
  MUX21H U440 ( .A(n62), .B(n56), .S(n425), .Z(N11) );
  MUX81P U441 ( .D0(n74), .D1(n70), .D2(n72), .D3(n68), .D4(n73), .D5(n69), 
        .D6(n71), .D7(n42), .A(n431), .B(n436), .C(n439), .Z(n75) );
  MUX21H U442 ( .A(n75), .B(n67), .S(n425), .Z(N12) );
  MUX81P U443 ( .D0(n88), .D1(n84), .D2(n86), .D3(n82), .D4(n87), .D5(n83), 
        .D6(n85), .D7(n81), .A(n431), .B(n436), .C(n440), .Z(n89) );
  MUX21H U444 ( .A(n89), .B(n80), .S(n425), .Z(N13) );
  MUX81P U445 ( .D0(n97), .D1(n93), .D2(n95), .D3(n91), .D4(n96), .D5(n92), 
        .D6(n94), .D7(n90), .A(n431), .B(n436), .C(n440), .Z(n98) );
  MUX81P U446 ( .D0(n106), .D1(n102), .D2(n104), .D3(n100), .D4(n105), .D5(
        n101), .D6(n103), .D7(n99), .A(n431), .B(n436), .C(n440), .Z(n107) );
  MUX21H U447 ( .A(n107), .B(n98), .S(n425), .Z(N14) );
  MUX81P U448 ( .D0(n524), .D1(n111), .D2(n113), .D3(n109), .D4(n524), .D5(
        n110), .D6(n112), .D7(n108), .A(n431), .B(n436), .C(n440), .Z(n114) );
  MUX81P U449 ( .D0(n120), .D1(n118), .D2(n481), .D3(n116), .D4(n119), .D5(
        n117), .D6(n482), .D7(n115), .A(n431), .B(n436), .C(n440), .Z(n121) );
  MUX21H U450 ( .A(n121), .B(n114), .S(n425), .Z(N15) );
  MUX81P U451 ( .D0(n133), .D1(n131), .D2(n525), .D3(n129), .D4(n132), .D5(
        n130), .D6(n525), .D7(n128), .A(n431), .B(n436), .C(n440), .Z(n134) );
  MUX21H U452 ( .A(n134), .B(n127), .S(n425), .Z(N16) );
  MUX81P U453 ( .D0(n142), .D1(n138), .D2(n140), .D3(n136), .D4(n141), .D5(
        n137), .D6(n139), .D7(n135), .A(n431), .B(n436), .C(n440), .Z(n143) );
  MUX21H U454 ( .A(n147), .B(n143), .S(n425), .Z(N17) );
  MUX81P U455 ( .D0(n155), .D1(n151), .D2(n153), .D3(n149), .D4(n154), .D5(
        n150), .D6(n152), .D7(n148), .A(n431), .B(n436), .C(n440), .Z(n156) );
  MUX81P U456 ( .D0(n163), .D1(n160), .D2(n465), .D3(n158), .D4(n162), .D5(
        n159), .D6(n161), .D7(n157), .A(n431), .B(n436), .C(n440), .Z(n164) );
  MUX21H U457 ( .A(n164), .B(n156), .S(n425), .Z(N18) );
  MUX81P U458 ( .D0(n172), .D1(n168), .D2(n170), .D3(n166), .D4(n171), .D5(
        n167), .D6(n169), .D7(n165), .A(n431), .B(n436), .C(n440), .Z(n173) );
  MUX81P U459 ( .D0(n525), .D1(n176), .D2(n178), .D3(n175), .D4(n179), .D5(n41), .D6(n177), .D7(n174), .A(n430), .B(n436), .C(n440), .Z(n180) );
  MUX21H U460 ( .A(n180), .B(n173), .S(n425), .Z(N19) );
  AN2P U461 ( .A(n526), .B(n460), .Z(n187) );
  AN2P U462 ( .A(n527), .B(n495), .Z(n215) );
  AN2P U463 ( .A(n527), .B(n495), .Z(n235) );
  AN2P U464 ( .A(n495), .B(n460), .Z(n239) );
  AN2P U465 ( .A(n527), .B(n460), .Z(n272) );
  AN2P U466 ( .A(n527), .B(n460), .Z(n284) );
  AN2P U467 ( .A(n527), .B(n495), .Z(n303) );
  AN2P U468 ( .A(n526), .B(n460), .Z(n311) );
  AN2P U469 ( .A(n526), .B(n495), .Z(n337) );
  AN2P U470 ( .A(n438), .B(n430), .Z(n354) );
  AN2P U471 ( .A(n64), .B(n430), .Z(n356) );
  AN2P U472 ( .A(n63), .B(n430), .Z(n357) );
  AN2P U473 ( .A(n438), .B(n65), .Z(n358) );
  AN2P U474 ( .A(n438), .B(n434), .Z(n373) );
  AN2P U475 ( .A(n434), .B(n54), .Z(n374) );
  AN2P U476 ( .A(n438), .B(n434), .Z(n379) );
  AN2P U477 ( .A(n430), .B(n51), .Z(n381) );
  AN2P U478 ( .A(n57), .B(n430), .Z(n388) );
  AN2P U479 ( .A(n59), .B(n438), .Z(n390) );
  AN2P U480 ( .A(n58), .B(n430), .Z(n391) );
  AN2P U481 ( .A(n438), .B(n430), .Z(n392) );
  AN2P U482 ( .A(n76), .B(n434), .Z(n403) );
  AN2P U483 ( .A(n510), .B(n434), .Z(n415) );
  AN2P U484 ( .A(n144), .B(n438), .Z(n416) );
  IV U485 ( .A(x[14]), .Z(n424) );
  IVA U486 ( .A(n542), .Z(n426) );
  IVA U487 ( .A(n542), .Z(n427) );
  IVA U488 ( .A(n542), .Z(n428) );
  IVA U489 ( .A(n542), .Z(n429) );
  IVP U490 ( .A(x[12]), .Z(n433) );
  IVA U491 ( .A(x[11]), .Z(n437) );
  IVA U492 ( .A(n472), .Z(n441) );
  IVA U493 ( .A(n472), .Z(n442) );
  IVA U494 ( .A(n472), .Z(n443) );
  IVA U495 ( .A(n472), .Z(n444) );
  IVA U496 ( .A(n473), .Z(n445) );
  IVA U497 ( .A(n473), .Z(n446) );
  IVA U498 ( .A(n473), .Z(n447) );
  IVA U499 ( .A(n473), .Z(n448) );
  IVA U500 ( .A(n473), .Z(n449) );
  IVA U501 ( .A(n474), .Z(n450) );
  IVA U502 ( .A(n474), .Z(n451) );
  IVA U503 ( .A(n474), .Z(n452) );
  IVA U504 ( .A(n474), .Z(n453) );
  IVA U505 ( .A(n474), .Z(n454) );
  IVA U506 ( .A(n475), .Z(n455) );
  IVA U507 ( .A(n475), .Z(n456) );
  IVA U508 ( .A(n475), .Z(n457) );
  IVA U509 ( .A(n475), .Z(n458) );
  IVA U510 ( .A(n475), .Z(n459) );
  IVP U511 ( .A(x[10]), .Z(n471) );
  IVA U512 ( .A(n505), .Z(n476) );
  IVA U513 ( .A(n505), .Z(n477) );
  IVA U514 ( .A(n505), .Z(n478) );
  IVA U515 ( .A(n505), .Z(n479) );
  IVA U516 ( .A(n506), .Z(n480) );
  IVA U517 ( .A(n506), .Z(n481) );
  IVA U518 ( .A(n506), .Z(n482) );
  IVA U519 ( .A(n506), .Z(n483) );
  IVA U520 ( .A(n506), .Z(n484) );
  IVA U521 ( .A(n507), .Z(n485) );
  IVA U522 ( .A(n507), .Z(n486) );
  IVA U523 ( .A(n507), .Z(n487) );
  IVA U524 ( .A(n507), .Z(n488) );
  IVA U525 ( .A(n507), .Z(n489) );
  IVA U526 ( .A(n508), .Z(n490) );
  IVA U527 ( .A(n508), .Z(n491) );
  IVA U528 ( .A(n508), .Z(n492) );
  IVA U529 ( .A(n508), .Z(n493) );
  IVA U530 ( .A(n508), .Z(n494) );
  IVP U531 ( .A(x[9]), .Z(n504) );
  IVA U532 ( .A(n536), .Z(n509) );
  IVA U533 ( .A(n536), .Z(n510) );
  IVA U534 ( .A(n537), .Z(n511) );
  IVA U535 ( .A(n537), .Z(n512) );
  IVA U536 ( .A(n537), .Z(n513) );
  IVA U537 ( .A(n538), .Z(n514) );
  IVA U538 ( .A(n538), .Z(n515) );
  IVA U539 ( .A(n538), .Z(n516) );
  IVA U540 ( .A(n539), .Z(n517) );
  IVA U541 ( .A(n539), .Z(n518) );
  IVA U542 ( .A(n539), .Z(n519) );
  IVA U543 ( .A(n540), .Z(n520) );
  IVA U544 ( .A(n540), .Z(n521) );
  IVA U545 ( .A(n540), .Z(n522) );
  IVA U546 ( .A(n541), .Z(n523) );
  IVA U547 ( .A(n541), .Z(n524) );
  IVA U548 ( .A(n541), .Z(n525) );
  IV U549 ( .A(n509), .Z(n526) );
  IVA U550 ( .A(x[8]), .Z(n535) );
  IVA U551 ( .A(n535), .Z(n536) );
  IVA U552 ( .A(n535), .Z(n537) );
  IVA U553 ( .A(n535), .Z(n538) );
  IVA U554 ( .A(n511), .Z(n539) );
  IVA U555 ( .A(n513), .Z(n540) );
  IVA U556 ( .A(n512), .Z(n541) );
  IVA U557 ( .A(n543), .Z(n542) );
  IV U558 ( .A(x[13]), .Z(n543) );
  EO U559 ( .A(Term1[25]), .B(\add_1242/carry[14] ), .Z(N50) );
  AN2 U560 ( .A(\add_1242/carry[13] ), .B(Term1[24]), .Z(\add_1242/carry[14] )
         );
  EO U561 ( .A(Term1[24]), .B(\add_1242/carry[13] ), .Z(N49) );
  AN2 U562 ( .A(\add_1242/carry[12] ), .B(Term1[23]), .Z(\add_1242/carry[13] )
         );
  EO U563 ( .A(Term1[23]), .B(\add_1242/carry[12] ), .Z(N48) );
  AN2 U564 ( .A(\add_1242/carry[11] ), .B(Term1[22]), .Z(\add_1242/carry[12] )
         );
  EO U565 ( .A(Term1[22]), .B(\add_1242/carry[11] ), .Z(N47) );
  AN2 U566 ( .A(\add_1242/carry[10] ), .B(Term1[21]), .Z(\add_1242/carry[11] )
         );
  EO U567 ( .A(Term1[21]), .B(\add_1242/carry[10] ), .Z(N46) );
  AN2 U568 ( .A(\add_1242/carry[9] ), .B(Term1[20]), .Z(\add_1242/carry[10] )
         );
  EO U569 ( .A(Term1[20]), .B(\add_1242/carry[9] ), .Z(N45) );
  AN2 U570 ( .A(\add_1242/carry[8] ), .B(Term1[19]), .Z(\add_1242/carry[9] )
         );
  EO U571 ( .A(Term1[19]), .B(\add_1242/carry[8] ), .Z(N44) );
  AN2 U572 ( .A(\add_1242/carry[7] ), .B(Term1[18]), .Z(\add_1242/carry[8] )
         );
  EO U573 ( .A(Term1[18]), .B(\add_1242/carry[7] ), .Z(N43) );
  AN2 U574 ( .A(\add_1242/carry[6] ), .B(Term1[17]), .Z(\add_1242/carry[7] )
         );
  EO U575 ( .A(Term1[17]), .B(\add_1242/carry[6] ), .Z(N42) );
  AN2 U576 ( .A(\add_1242/carry[5] ), .B(Term1[16]), .Z(\add_1242/carry[6] )
         );
  EO U577 ( .A(Term1[16]), .B(\add_1242/carry[5] ), .Z(N41) );
  AN2 U578 ( .A(\add_1242/carry[4] ), .B(Term1[15]), .Z(\add_1242/carry[5] )
         );
  EO U579 ( .A(Term1[15]), .B(\add_1242/carry[4] ), .Z(N40) );
  AN2 U580 ( .A(\add_1242/carry[3] ), .B(Term1[14]), .Z(\add_1242/carry[4] )
         );
  EO U581 ( .A(Term1[14]), .B(\add_1242/carry[3] ), .Z(N39) );
  AN2 U582 ( .A(\add_1242/carry[2] ), .B(Term1[13]), .Z(\add_1242/carry[3] )
         );
  EO U583 ( .A(Term1[13]), .B(\add_1242/carry[2] ), .Z(N38) );
  AN2 U584 ( .A(\add_1242/carry[1] ), .B(Term1[12]), .Z(\add_1242/carry[2] )
         );
  EO U585 ( .A(Term1[12]), .B(\add_1242/carry[1] ), .Z(N37) );
  AN2 U586 ( .A(\Term2[18] ), .B(Term1[11]), .Z(\add_1242/carry[1] ) );
  EO U587 ( .A(Term1[11]), .B(\Term2[18] ), .Z(N36) );
endmodule


module SinBlock_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   \A[9] , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59;
  assign SUM[10] = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];

  OR2P U2 ( .A(B[11]), .B(A[11]), .Z(n1) );
  AN2P U3 ( .A(n1), .B(n59), .Z(SUM[11]) );
  IVP U4 ( .A(n57), .Z(n13) );
  IVP U5 ( .A(n50), .Z(n11) );
  IVP U6 ( .A(n42), .Z(n9) );
  IVP U7 ( .A(n34), .Z(n7) );
  IVP U8 ( .A(n26), .Z(n5) );
  IVP U9 ( .A(n59), .Z(n14) );
  IVP U10 ( .A(n22), .Z(n4) );
  IVP U11 ( .A(n30), .Z(n6) );
  IVP U12 ( .A(n38), .Z(n8) );
  IVP U13 ( .A(n46), .Z(n10) );
  IVP U14 ( .A(n54), .Z(n12) );
  IVP U15 ( .A(n18), .Z(n3) );
  EN U16 ( .A(B[23]), .B(n15), .Z(SUM[23]) );
  AO6 U17 ( .A(n16), .B(n3), .C(n17), .Z(n15) );
  EO U18 ( .A(n16), .B(n19), .Z(SUM[22]) );
  NR2 U19 ( .A(n17), .B(n18), .Z(n19) );
  NR2 U20 ( .A(B[22]), .B(A[22]), .Z(n18) );
  AN2 U21 ( .A(B[22]), .B(A[22]), .Z(n17) );
  AO7 U22 ( .A(n20), .B(n21), .C(n22), .Z(n16) );
  EN U23 ( .A(n21), .B(n23), .Z(SUM[21]) );
  NR2 U24 ( .A(n4), .B(n20), .Z(n23) );
  NR2 U25 ( .A(B[21]), .B(A[21]), .Z(n20) );
  ND2 U26 ( .A(B[21]), .B(A[21]), .Z(n22) );
  AO6 U27 ( .A(n5), .B(n24), .C(n25), .Z(n21) );
  EO U28 ( .A(n24), .B(n27), .Z(SUM[20]) );
  NR2 U29 ( .A(n25), .B(n26), .Z(n27) );
  NR2 U30 ( .A(B[20]), .B(A[20]), .Z(n26) );
  AN2 U31 ( .A(B[20]), .B(A[20]), .Z(n25) );
  AO7 U32 ( .A(n28), .B(n29), .C(n30), .Z(n24) );
  EN U33 ( .A(n29), .B(n31), .Z(SUM[19]) );
  NR2 U34 ( .A(n6), .B(n28), .Z(n31) );
  NR2 U35 ( .A(B[19]), .B(A[19]), .Z(n28) );
  ND2 U36 ( .A(B[19]), .B(A[19]), .Z(n30) );
  AO6 U37 ( .A(n7), .B(n32), .C(n33), .Z(n29) );
  EO U38 ( .A(n32), .B(n35), .Z(SUM[18]) );
  NR2 U39 ( .A(n33), .B(n34), .Z(n35) );
  NR2 U40 ( .A(B[18]), .B(A[18]), .Z(n34) );
  AN2 U41 ( .A(B[18]), .B(A[18]), .Z(n33) );
  AO7 U42 ( .A(n36), .B(n37), .C(n38), .Z(n32) );
  EN U43 ( .A(n37), .B(n39), .Z(SUM[17]) );
  NR2 U44 ( .A(n8), .B(n36), .Z(n39) );
  NR2 U45 ( .A(B[17]), .B(A[17]), .Z(n36) );
  ND2 U46 ( .A(B[17]), .B(A[17]), .Z(n38) );
  AO6 U47 ( .A(n9), .B(n40), .C(n41), .Z(n37) );
  EO U48 ( .A(n40), .B(n43), .Z(SUM[16]) );
  NR2 U49 ( .A(n41), .B(n42), .Z(n43) );
  NR2 U50 ( .A(B[16]), .B(A[16]), .Z(n42) );
  AN2 U51 ( .A(B[16]), .B(A[16]), .Z(n41) );
  AO7 U52 ( .A(n44), .B(n45), .C(n46), .Z(n40) );
  EN U53 ( .A(n45), .B(n47), .Z(SUM[15]) );
  NR2 U54 ( .A(n10), .B(n44), .Z(n47) );
  NR2 U55 ( .A(B[15]), .B(A[15]), .Z(n44) );
  ND2 U56 ( .A(B[15]), .B(A[15]), .Z(n46) );
  AO6 U57 ( .A(n11), .B(n48), .C(n49), .Z(n45) );
  EO U58 ( .A(n48), .B(n51), .Z(SUM[14]) );
  NR2 U59 ( .A(n49), .B(n50), .Z(n51) );
  NR2 U60 ( .A(B[14]), .B(A[14]), .Z(n50) );
  AN2 U61 ( .A(B[14]), .B(A[14]), .Z(n49) );
  AO7 U62 ( .A(n52), .B(n53), .C(n54), .Z(n48) );
  EN U63 ( .A(n53), .B(n55), .Z(SUM[13]) );
  NR2 U64 ( .A(n12), .B(n52), .Z(n55) );
  NR2 U65 ( .A(B[13]), .B(A[13]), .Z(n52) );
  ND2 U66 ( .A(B[13]), .B(A[13]), .Z(n54) );
  AO6 U67 ( .A(n13), .B(n14), .C(n56), .Z(n53) );
  EO U68 ( .A(n14), .B(n58), .Z(SUM[12]) );
  NR2 U69 ( .A(n56), .B(n57), .Z(n58) );
  NR2 U70 ( .A(B[12]), .B(A[12]), .Z(n57) );
  AN2 U71 ( .A(B[12]), .B(A[12]), .Z(n56) );
  ND2 U72 ( .A(B[11]), .B(A[11]), .Z(n59) );
endmodule


module SinBlock_1_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [11:0] A;
  input [13:0] B;
  output [25:0] PRODUCT;
  input TC;
  wire   \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][13] ,
         \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] ,
         \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] ,
         \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][13] , \ab[8][12] , \ab[8][11] ,
         \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] , \ab[8][6] ,
         \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] ,
         \ab[8][0] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][13] ,
         \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] ,
         \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] ,
         \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][13] , \ab[3][12] , \ab[3][11] ,
         \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[0][13] , \ab[0][12] ,
         \ab[0][11] , \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] ,
         \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] ,
         \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] ,
         \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] ,
         \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] ,
         \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] ,
         \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][12] , \CARRYB[1][11] ,
         \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] ,
         \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[11][0] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][12] ,
         \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] ,
         \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] ,
         \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][12] ,
         \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] ,
         \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] ,
         \A2[17] , \A2[16] , \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] ,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8;

  SinBlock_1_DW01_add_1 FS_1 ( .A({1'b0, \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \SUMB[11][0] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[23] , 
        \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , 
        \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        PRODUCT[25:11], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8}) );
  FA1A S5_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\ab[10][13] ), .CO(
        \CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S3_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\ab[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S3_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\ab[8][13] ), .CO(
        \CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S3_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\ab[7][13] ), .CO(
        \CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S3_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\ab[6][13] ), .CO(
        \CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S3_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\ab[5][13] ), .CO(
        \CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S3_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\ab[4][13] ), .CO(
        \CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S3_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\ab[3][13] ), .CO(
        \CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S3_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\ab[2][13] ), .CO(
        \CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S3_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\ab[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S4_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(
        \CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S4_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), .CO(
        \CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S4_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(
        \CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S4_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(
        \CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S4_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(
        \CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S4_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(
        \CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S4_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(
        \CARRYB[11][0] ), .S(\SUMB[11][0] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S4_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(
        \CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S4_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(
        \CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(
        \CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  IVP U2 ( .A(A[0]), .Z(n10) );
  EO U3 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A1[12] ) );
  EO U4 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  EO U5 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A1[11] ) );
  EO U6 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A1[13] ) );
  EO U7 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A1[14] ) );
  EO U8 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A1[15] ) );
  EO U9 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A1[16] ) );
  EO U10 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A1[17] ) );
  EO U11 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A1[18] ) );
  EO U12 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A1[19] ) );
  EO U13 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A1[20] ) );
  EO U14 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A1[21] ) );
  EO U15 ( .A(\CARRYB[11][12] ), .B(\ab[11][13] ), .Z(\A1[22] ) );
  EO U16 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A1[10] ) );
  IVP U17 ( .A(A[1]), .Z(n11) );
  EO U18 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U19 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  IVP U20 ( .A(A[2]), .Z(n12) );
  EO U21 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U22 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U23 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  IVP U24 ( .A(A[3]), .Z(n13) );
  EO U25 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U26 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U27 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  IVP U28 ( .A(A[4]), .Z(n14) );
  EO U29 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U30 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  IVP U31 ( .A(A[5]), .Z(n15) );
  EO U32 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  IVP U33 ( .A(A[6]), .Z(n16) );
  IVP U34 ( .A(A[7]), .Z(n17) );
  IVP U35 ( .A(A[8]), .Z(n18) );
  IVP U36 ( .A(B[13]), .Z(n8) );
  IVP U37 ( .A(A[9]), .Z(n19) );
  IVP U38 ( .A(A[10]), .Z(n20) );
  IVP U39 ( .A(A[11]), .Z(n9) );
  IVP U40 ( .A(B[2]), .Z(n26) );
  IVP U41 ( .A(B[3]), .Z(n25) );
  IVP U42 ( .A(B[4]), .Z(n24) );
  IVP U43 ( .A(B[1]), .Z(n27) );
  IVP U44 ( .A(B[5]), .Z(n23) );
  IVP U45 ( .A(B[6]), .Z(n22) );
  IVP U46 ( .A(B[7]), .Z(n21) );
  IVP U47 ( .A(B[0]), .Z(n28) );
  IVP U48 ( .A(B[8]), .Z(n3) );
  IVP U49 ( .A(B[9]), .Z(n4) );
  IVP U50 ( .A(B[10]), .Z(n5) );
  IVP U51 ( .A(B[11]), .Z(n6) );
  IVP U52 ( .A(B[12]), .Z(n7) );
  AN2P U53 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A2[11] ) );
  AN2P U54 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A2[13] ) );
  AN2P U55 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A2[14] ) );
  AN2P U56 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A2[15] ) );
  AN2P U57 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A2[16] ) );
  AN2P U58 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A2[17] ) );
  AN2P U59 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A2[18] ) );
  AN2P U60 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A2[19] ) );
  AN2P U61 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A2[20] ) );
  AN2P U62 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A2[21] ) );
  AN2P U63 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A2[22] ) );
  AN2P U64 ( .A(\CARRYB[11][12] ), .B(\ab[11][13] ), .Z(\A2[23] ) );
  AN2P U65 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U66 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U67 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U68 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U69 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U70 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U71 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U72 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U73 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U74 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U75 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U76 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U77 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A2[12] ) );
  NR2 U79 ( .A(n19), .B(n4), .Z(\ab[9][9] ) );
  NR2 U80 ( .A(n19), .B(n3), .Z(\ab[9][8] ) );
  NR2 U81 ( .A(n19), .B(n21), .Z(\ab[9][7] ) );
  NR2 U82 ( .A(n19), .B(n22), .Z(\ab[9][6] ) );
  NR2 U83 ( .A(n19), .B(n23), .Z(\ab[9][5] ) );
  NR2 U84 ( .A(n19), .B(n24), .Z(\ab[9][4] ) );
  NR2 U85 ( .A(n19), .B(n25), .Z(\ab[9][3] ) );
  NR2 U86 ( .A(n19), .B(n26), .Z(\ab[9][2] ) );
  NR2 U87 ( .A(n19), .B(n27), .Z(\ab[9][1] ) );
  NR2 U88 ( .A(n19), .B(n8), .Z(\ab[9][13] ) );
  NR2 U89 ( .A(n19), .B(n7), .Z(\ab[9][12] ) );
  NR2 U90 ( .A(n19), .B(n6), .Z(\ab[9][11] ) );
  NR2 U91 ( .A(n19), .B(n5), .Z(\ab[9][10] ) );
  NR2 U92 ( .A(n19), .B(n28), .Z(\ab[9][0] ) );
  NR2 U93 ( .A(n4), .B(n18), .Z(\ab[8][9] ) );
  NR2 U94 ( .A(n3), .B(n18), .Z(\ab[8][8] ) );
  NR2 U95 ( .A(n21), .B(n18), .Z(\ab[8][7] ) );
  NR2 U96 ( .A(n22), .B(n18), .Z(\ab[8][6] ) );
  NR2 U97 ( .A(n23), .B(n18), .Z(\ab[8][5] ) );
  NR2 U98 ( .A(n24), .B(n18), .Z(\ab[8][4] ) );
  NR2 U99 ( .A(n25), .B(n18), .Z(\ab[8][3] ) );
  NR2 U100 ( .A(n26), .B(n18), .Z(\ab[8][2] ) );
  NR2 U101 ( .A(n27), .B(n18), .Z(\ab[8][1] ) );
  NR2 U102 ( .A(n8), .B(n18), .Z(\ab[8][13] ) );
  NR2 U103 ( .A(n7), .B(n18), .Z(\ab[8][12] ) );
  NR2 U104 ( .A(n6), .B(n18), .Z(\ab[8][11] ) );
  NR2 U105 ( .A(n5), .B(n18), .Z(\ab[8][10] ) );
  NR2 U106 ( .A(n28), .B(n18), .Z(\ab[8][0] ) );
  NR2 U107 ( .A(n4), .B(n17), .Z(\ab[7][9] ) );
  NR2 U108 ( .A(n3), .B(n17), .Z(\ab[7][8] ) );
  NR2 U109 ( .A(n21), .B(n17), .Z(\ab[7][7] ) );
  NR2 U110 ( .A(n22), .B(n17), .Z(\ab[7][6] ) );
  NR2 U111 ( .A(n23), .B(n17), .Z(\ab[7][5] ) );
  NR2 U112 ( .A(n24), .B(n17), .Z(\ab[7][4] ) );
  NR2 U113 ( .A(n25), .B(n17), .Z(\ab[7][3] ) );
  NR2 U114 ( .A(n26), .B(n17), .Z(\ab[7][2] ) );
  NR2 U115 ( .A(n27), .B(n17), .Z(\ab[7][1] ) );
  NR2 U116 ( .A(n8), .B(n17), .Z(\ab[7][13] ) );
  NR2 U117 ( .A(n7), .B(n17), .Z(\ab[7][12] ) );
  NR2 U118 ( .A(n6), .B(n17), .Z(\ab[7][11] ) );
  NR2 U119 ( .A(n5), .B(n17), .Z(\ab[7][10] ) );
  NR2 U120 ( .A(n28), .B(n17), .Z(\ab[7][0] ) );
  NR2 U121 ( .A(n4), .B(n16), .Z(\ab[6][9] ) );
  NR2 U122 ( .A(n3), .B(n16), .Z(\ab[6][8] ) );
  NR2 U123 ( .A(n21), .B(n16), .Z(\ab[6][7] ) );
  NR2 U124 ( .A(n22), .B(n16), .Z(\ab[6][6] ) );
  NR2 U125 ( .A(n23), .B(n16), .Z(\ab[6][5] ) );
  NR2 U126 ( .A(n24), .B(n16), .Z(\ab[6][4] ) );
  NR2 U127 ( .A(n25), .B(n16), .Z(\ab[6][3] ) );
  NR2 U128 ( .A(n26), .B(n16), .Z(\ab[6][2] ) );
  NR2 U129 ( .A(n27), .B(n16), .Z(\ab[6][1] ) );
  NR2 U130 ( .A(n8), .B(n16), .Z(\ab[6][13] ) );
  NR2 U131 ( .A(n7), .B(n16), .Z(\ab[6][12] ) );
  NR2 U132 ( .A(n6), .B(n16), .Z(\ab[6][11] ) );
  NR2 U133 ( .A(n5), .B(n16), .Z(\ab[6][10] ) );
  NR2 U134 ( .A(n28), .B(n16), .Z(\ab[6][0] ) );
  NR2 U135 ( .A(n4), .B(n15), .Z(\ab[5][9] ) );
  NR2 U136 ( .A(n3), .B(n15), .Z(\ab[5][8] ) );
  NR2 U137 ( .A(n21), .B(n15), .Z(\ab[5][7] ) );
  NR2 U138 ( .A(n22), .B(n15), .Z(\ab[5][6] ) );
  NR2 U139 ( .A(n23), .B(n15), .Z(\ab[5][5] ) );
  NR2 U140 ( .A(n24), .B(n15), .Z(\ab[5][4] ) );
  NR2 U141 ( .A(n25), .B(n15), .Z(\ab[5][3] ) );
  NR2 U142 ( .A(n26), .B(n15), .Z(\ab[5][2] ) );
  NR2 U143 ( .A(n27), .B(n15), .Z(\ab[5][1] ) );
  NR2 U144 ( .A(n8), .B(n15), .Z(\ab[5][13] ) );
  NR2 U145 ( .A(n7), .B(n15), .Z(\ab[5][12] ) );
  NR2 U146 ( .A(n6), .B(n15), .Z(\ab[5][11] ) );
  NR2 U147 ( .A(n5), .B(n15), .Z(\ab[5][10] ) );
  NR2 U148 ( .A(n28), .B(n15), .Z(\ab[5][0] ) );
  NR2 U149 ( .A(n4), .B(n14), .Z(\ab[4][9] ) );
  NR2 U150 ( .A(n3), .B(n14), .Z(\ab[4][8] ) );
  NR2 U151 ( .A(n21), .B(n14), .Z(\ab[4][7] ) );
  NR2 U152 ( .A(n22), .B(n14), .Z(\ab[4][6] ) );
  NR2 U153 ( .A(n23), .B(n14), .Z(\ab[4][5] ) );
  NR2 U154 ( .A(n24), .B(n14), .Z(\ab[4][4] ) );
  NR2 U155 ( .A(n25), .B(n14), .Z(\ab[4][3] ) );
  NR2 U156 ( .A(n26), .B(n14), .Z(\ab[4][2] ) );
  NR2 U157 ( .A(n27), .B(n14), .Z(\ab[4][1] ) );
  NR2 U158 ( .A(n8), .B(n14), .Z(\ab[4][13] ) );
  NR2 U159 ( .A(n7), .B(n14), .Z(\ab[4][12] ) );
  NR2 U160 ( .A(n6), .B(n14), .Z(\ab[4][11] ) );
  NR2 U161 ( .A(n5), .B(n14), .Z(\ab[4][10] ) );
  NR2 U162 ( .A(n28), .B(n14), .Z(\ab[4][0] ) );
  NR2 U163 ( .A(n4), .B(n13), .Z(\ab[3][9] ) );
  NR2 U164 ( .A(n3), .B(n13), .Z(\ab[3][8] ) );
  NR2 U165 ( .A(n21), .B(n13), .Z(\ab[3][7] ) );
  NR2 U166 ( .A(n22), .B(n13), .Z(\ab[3][6] ) );
  NR2 U167 ( .A(n23), .B(n13), .Z(\ab[3][5] ) );
  NR2 U168 ( .A(n24), .B(n13), .Z(\ab[3][4] ) );
  NR2 U169 ( .A(n25), .B(n13), .Z(\ab[3][3] ) );
  NR2 U170 ( .A(n26), .B(n13), .Z(\ab[3][2] ) );
  NR2 U171 ( .A(n27), .B(n13), .Z(\ab[3][1] ) );
  NR2 U172 ( .A(n8), .B(n13), .Z(\ab[3][13] ) );
  NR2 U173 ( .A(n7), .B(n13), .Z(\ab[3][12] ) );
  NR2 U174 ( .A(n6), .B(n13), .Z(\ab[3][11] ) );
  NR2 U175 ( .A(n5), .B(n13), .Z(\ab[3][10] ) );
  NR2 U176 ( .A(n28), .B(n13), .Z(\ab[3][0] ) );
  NR2 U177 ( .A(n4), .B(n12), .Z(\ab[2][9] ) );
  NR2 U178 ( .A(n3), .B(n12), .Z(\ab[2][8] ) );
  NR2 U179 ( .A(n21), .B(n12), .Z(\ab[2][7] ) );
  NR2 U180 ( .A(n22), .B(n12), .Z(\ab[2][6] ) );
  NR2 U181 ( .A(n23), .B(n12), .Z(\ab[2][5] ) );
  NR2 U182 ( .A(n24), .B(n12), .Z(\ab[2][4] ) );
  NR2 U183 ( .A(n25), .B(n12), .Z(\ab[2][3] ) );
  NR2 U184 ( .A(n26), .B(n12), .Z(\ab[2][2] ) );
  NR2 U185 ( .A(n27), .B(n12), .Z(\ab[2][1] ) );
  NR2 U186 ( .A(n8), .B(n12), .Z(\ab[2][13] ) );
  NR2 U187 ( .A(n7), .B(n12), .Z(\ab[2][12] ) );
  NR2 U188 ( .A(n6), .B(n12), .Z(\ab[2][11] ) );
  NR2 U189 ( .A(n5), .B(n12), .Z(\ab[2][10] ) );
  NR2 U190 ( .A(n28), .B(n12), .Z(\ab[2][0] ) );
  NR2 U191 ( .A(n4), .B(n11), .Z(\ab[1][9] ) );
  NR2 U192 ( .A(n3), .B(n11), .Z(\ab[1][8] ) );
  NR2 U193 ( .A(n21), .B(n11), .Z(\ab[1][7] ) );
  NR2 U194 ( .A(n22), .B(n11), .Z(\ab[1][6] ) );
  NR2 U195 ( .A(n23), .B(n11), .Z(\ab[1][5] ) );
  NR2 U196 ( .A(n24), .B(n11), .Z(\ab[1][4] ) );
  NR2 U197 ( .A(n25), .B(n11), .Z(\ab[1][3] ) );
  NR2 U198 ( .A(n26), .B(n11), .Z(\ab[1][2] ) );
  NR2 U199 ( .A(n8), .B(n11), .Z(\ab[1][13] ) );
  NR2 U200 ( .A(n7), .B(n11), .Z(\ab[1][12] ) );
  NR2 U201 ( .A(n6), .B(n11), .Z(\ab[1][11] ) );
  NR2 U202 ( .A(n5), .B(n11), .Z(\ab[1][10] ) );
  NR2 U203 ( .A(n4), .B(n9), .Z(\ab[11][9] ) );
  NR2 U204 ( .A(n3), .B(n9), .Z(\ab[11][8] ) );
  NR2 U205 ( .A(n21), .B(n9), .Z(\ab[11][7] ) );
  NR2 U206 ( .A(n22), .B(n9), .Z(\ab[11][6] ) );
  NR2 U207 ( .A(n23), .B(n9), .Z(\ab[11][5] ) );
  NR2 U208 ( .A(n24), .B(n9), .Z(\ab[11][4] ) );
  NR2 U209 ( .A(n25), .B(n9), .Z(\ab[11][3] ) );
  NR2 U210 ( .A(n26), .B(n9), .Z(\ab[11][2] ) );
  NR2 U211 ( .A(n27), .B(n9), .Z(\ab[11][1] ) );
  NR2 U212 ( .A(n8), .B(n9), .Z(\ab[11][13] ) );
  NR2 U213 ( .A(n7), .B(n9), .Z(\ab[11][12] ) );
  NR2 U214 ( .A(n6), .B(n9), .Z(\ab[11][11] ) );
  NR2 U215 ( .A(n5), .B(n9), .Z(\ab[11][10] ) );
  NR2 U216 ( .A(n28), .B(n9), .Z(\ab[11][0] ) );
  NR2 U217 ( .A(n4), .B(n20), .Z(\ab[10][9] ) );
  NR2 U218 ( .A(n3), .B(n20), .Z(\ab[10][8] ) );
  NR2 U219 ( .A(n21), .B(n20), .Z(\ab[10][7] ) );
  NR2 U220 ( .A(n22), .B(n20), .Z(\ab[10][6] ) );
  NR2 U221 ( .A(n23), .B(n20), .Z(\ab[10][5] ) );
  NR2 U222 ( .A(n24), .B(n20), .Z(\ab[10][4] ) );
  NR2 U223 ( .A(n25), .B(n20), .Z(\ab[10][3] ) );
  NR2 U224 ( .A(n26), .B(n20), .Z(\ab[10][2] ) );
  NR2 U225 ( .A(n27), .B(n20), .Z(\ab[10][1] ) );
  NR2 U226 ( .A(n8), .B(n20), .Z(\ab[10][13] ) );
  NR2 U227 ( .A(n7), .B(n20), .Z(\ab[10][12] ) );
  NR2 U228 ( .A(n6), .B(n20), .Z(\ab[10][11] ) );
  NR2 U229 ( .A(n5), .B(n20), .Z(\ab[10][10] ) );
  NR2 U230 ( .A(n28), .B(n20), .Z(\ab[10][0] ) );
  NR2 U231 ( .A(n4), .B(n10), .Z(\ab[0][9] ) );
  NR2 U232 ( .A(n3), .B(n10), .Z(\ab[0][8] ) );
  NR2 U233 ( .A(n21), .B(n10), .Z(\ab[0][7] ) );
  NR2 U234 ( .A(n22), .B(n10), .Z(\ab[0][6] ) );
  NR2 U235 ( .A(n23), .B(n10), .Z(\ab[0][5] ) );
  NR2 U236 ( .A(n24), .B(n10), .Z(\ab[0][4] ) );
  NR2 U237 ( .A(n25), .B(n10), .Z(\ab[0][3] ) );
  NR2 U238 ( .A(n26), .B(n10), .Z(\ab[0][2] ) );
  NR2 U239 ( .A(n8), .B(n10), .Z(\ab[0][13] ) );
  NR2 U240 ( .A(n7), .B(n10), .Z(\ab[0][12] ) );
  NR2 U241 ( .A(n6), .B(n10), .Z(\ab[0][11] ) );
  NR2 U242 ( .A(n5), .B(n10), .Z(\ab[0][10] ) );
  AN3 U243 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U244 ( .A(n11), .B(n27), .Z(\ab[1][1] ) );
endmodule


module SinBlock_1 ( clk, reset, func, x, sinValue );
  input [15:0] x;
  output [15:0] sinValue;
  input clk, reset, func;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         \Term2[18] , N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, sValue, N57, \add_1242/carry[14] ,
         \add_1242/carry[13] , \add_1242/carry[12] , \add_1242/carry[11] ,
         \add_1242/carry[10] , \add_1242/carry[9] , \add_1242/carry[8] ,
         \add_1242/carry[7] , \add_1242/carry[6] , \add_1242/carry[5] ,
         \add_1242/carry[4] , \add_1242/carry[3] , \add_1242/carry[2] ,
         \add_1242/carry[1] , n34, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n547;
  wire   [25:11] Term1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10;

  SinBlock_1_DW02_mult_0 mult_1238 ( .A({n40, N9, N10, N11, N12, N13, N14, N15, 
        N16, N17, N18, N19}), .B({n542, x[12:0]}), .TC(1'b0), .PRODUCT({N34, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  FDS2L \Term1_reg[25]  ( .CR(1'b1), .D(N34), .LD(n544), .CP(clk), .Q(
        Term1[25]) );
  FDS2L \Term1_reg[24]  ( .CR(1'b1), .D(N33), .LD(n544), .CP(clk), .Q(
        Term1[24]) );
  FDS2L \Term1_reg[23]  ( .CR(1'b1), .D(N32), .LD(n544), .CP(clk), .Q(
        Term1[23]) );
  FDS2L \Term1_reg[22]  ( .CR(1'b1), .D(N31), .LD(n544), .CP(clk), .Q(
        Term1[22]) );
  FDS2L \Term1_reg[21]  ( .CR(1'b1), .D(N30), .LD(n544), .CP(clk), .Q(
        Term1[21]) );
  FDS2L \Term1_reg[20]  ( .CR(1'b1), .D(N29), .LD(n544), .CP(clk), .Q(
        Term1[20]) );
  FDS2L \Term1_reg[19]  ( .CR(1'b1), .D(N28), .LD(n544), .CP(clk), .Q(
        Term1[19]) );
  FDS2L \Term1_reg[18]  ( .CR(1'b1), .D(N27), .LD(n544), .CP(clk), .Q(
        Term1[18]) );
  FDS2L \Term1_reg[17]  ( .CR(1'b1), .D(N26), .LD(n544), .CP(clk), .Q(
        Term1[17]) );
  FDS2L \Term1_reg[16]  ( .CR(1'b1), .D(N25), .LD(n544), .CP(clk), .Q(
        Term1[16]) );
  FDS2L \Term1_reg[15]  ( .CR(1'b1), .D(N24), .LD(n544), .CP(clk), .Q(
        Term1[15]) );
  FDS2L \Term1_reg[14]  ( .CR(1'b1), .D(N23), .LD(n544), .CP(clk), .Q(
        Term1[14]) );
  FDS2L \Term1_reg[13]  ( .CR(1'b1), .D(N22), .LD(n544), .CP(clk), .Q(
        Term1[13]) );
  FDS2L \Term1_reg[12]  ( .CR(1'b1), .D(N21), .LD(n544), .CP(clk), .Q(
        Term1[12]) );
  FDS2L \Term1_reg[11]  ( .CR(1'b1), .D(N20), .LD(n544), .CP(clk), .Q(
        Term1[11]) );
  FDS2L \Term2_reg[18]  ( .CR(1'b1), .D(1'b1), .LD(n544), .CP(clk), .Q(
        \Term2[18] ) );
  FDS2L \sinValue_reg[14]  ( .CR(1'b1), .D(N50), .LD(n544), .CP(clk), .Q(
        sinValue[14]) );
  FDS2L \sinValue_reg[13]  ( .CR(1'b1), .D(N49), .LD(n544), .CP(clk), .Q(
        sinValue[13]) );
  FDS2L \sinValue_reg[12]  ( .CR(1'b1), .D(N48), .LD(n544), .CP(clk), .Q(
        sinValue[12]) );
  FDS2L \sinValue_reg[11]  ( .CR(1'b1), .D(N47), .LD(n544), .CP(clk), .Q(
        sinValue[11]) );
  FDS2L \sinValue_reg[10]  ( .CR(1'b1), .D(N46), .LD(n544), .CP(clk), .Q(
        sinValue[10]) );
  FDS2L \sinValue_reg[9]  ( .CR(1'b1), .D(N45), .LD(n544), .CP(clk), .Q(
        sinValue[9]) );
  FDS2L \sinValue_reg[8]  ( .CR(1'b1), .D(N44), .LD(n544), .CP(clk), .Q(
        sinValue[8]) );
  FDS2L \sinValue_reg[7]  ( .CR(1'b1), .D(N43), .LD(n544), .CP(clk), .Q(
        sinValue[7]) );
  FDS2L \sinValue_reg[6]  ( .CR(1'b1), .D(N42), .LD(n544), .CP(clk), .Q(
        sinValue[6]) );
  FDS2L \sinValue_reg[5]  ( .CR(1'b1), .D(N41), .LD(n544), .CP(clk), .Q(
        sinValue[5]) );
  FDS2L \sinValue_reg[4]  ( .CR(1'b1), .D(N40), .LD(n544), .CP(clk), .Q(
        sinValue[4]) );
  FDS2L \sinValue_reg[3]  ( .CR(1'b1), .D(N39), .LD(n544), .CP(clk), .Q(
        sinValue[3]) );
  FDS2L \sinValue_reg[2]  ( .CR(1'b1), .D(N38), .LD(n544), .CP(clk), .Q(
        sinValue[2]) );
  FDS2L \sinValue_reg[1]  ( .CR(1'b1), .D(N37), .LD(n544), .CP(clk), .Q(
        sinValue[1]) );
  FDS2L \sinValue_reg[0]  ( .CR(1'b1), .D(N36), .LD(n544), .CP(clk), .Q(
        sinValue[0]) );
  FDS2L sValue_reg ( .CR(1'b1), .D(N57), .LD(n544), .CP(clk), .Q(sValue) );
  FDS2L \sinValue_reg[15]  ( .CR(1'b1), .D(sValue), .LD(n544), .CP(clk), .Q(
        sinValue[15]) );
  AN2P U3 ( .A(n339), .B(n338), .Z(n34) );
  AN2P U4 ( .A(n300), .B(n299), .Z(n36) );
  AN2P U5 ( .A(n243), .B(n242), .Z(n37) );
  AN2P U6 ( .A(n258), .B(n257), .Z(n38) );
  AN2P U7 ( .A(n324), .B(n323), .Z(n39) );
  AN2P U8 ( .A(n425), .B(n44), .Z(n40) );
  NR2 U9 ( .A(n463), .B(n503), .Z(n186) );
  NR2 U10 ( .A(n500), .B(n465), .Z(n229) );
  NR2 U11 ( .A(n532), .B(n500), .Z(n231) );
  EO U12 ( .A(n527), .B(n495), .Z(n163) );
  ND2 U13 ( .A(n529), .B(n332), .Z(n179) );
  ND2 U14 ( .A(n496), .B(n461), .Z(n332) );
  ND2 U15 ( .A(n502), .B(n203), .Z(n150) );
  ND2 U16 ( .A(n534), .B(n462), .Z(n203) );
  ND2 U17 ( .A(n334), .B(n333), .Z(n162) );
  ND2 U18 ( .A(n528), .B(n460), .Z(n333) );
  EN U19 ( .A(n527), .B(n496), .Z(n334) );
  ND2 U20 ( .A(n468), .B(n530), .Z(n289) );
  AN2P U21 ( .A(n530), .B(n468), .Z(n41) );
  MUX21L U22 ( .A(n530), .B(n503), .S(n464), .Z(n148) );
  MUX21L U23 ( .A(n500), .B(n465), .S(n532), .Z(n153) );
  MUX21L U24 ( .A(n530), .B(n288), .S(n497), .Z(n290) );
  NR2 U25 ( .A(n529), .B(n468), .Z(n288) );
  ND2 U26 ( .A(n266), .B(n265), .Z(n144) );
  ND2 U27 ( .A(n466), .B(n498), .Z(n265) );
  MUX21L U28 ( .A(n264), .B(n499), .S(n531), .Z(n266) );
  NR2 U29 ( .A(n499), .B(n466), .Z(n264) );
  AO4 U30 ( .A(n496), .B(n462), .C(n528), .D(n461), .Z(n146) );
  AO4 U31 ( .A(n529), .B(n469), .C(n529), .D(n497), .Z(n176) );
  AO7 U32 ( .A(n528), .B(n496), .C(n470), .Z(n161) );
  AO7 U33 ( .A(n532), .B(n500), .C(n465), .Z(n141) );
  ND2 U34 ( .A(n497), .B(n302), .Z(n160) );
  ND2 U35 ( .A(n529), .B(n469), .Z(n302) );
  ND2 U36 ( .A(n225), .B(n224), .Z(n139) );
  ND2 U37 ( .A(n461), .B(n501), .Z(n224) );
  MUX21L U38 ( .A(n223), .B(n501), .S(n533), .Z(n225) );
  NR2 U39 ( .A(n501), .B(n462), .Z(n223) );
  EO U40 ( .A(n495), .B(n465), .Z(n245) );
  EN U41 ( .A(n527), .B(n498), .Z(n129) );
  EN U42 ( .A(n527), .B(n469), .Z(n131) );
  NR2 U43 ( .A(n530), .B(n467), .Z(n285) );
  ND2 U44 ( .A(n228), .B(n227), .Z(n112) );
  ND2 U45 ( .A(n461), .B(n501), .Z(n227) );
  MUX21L U46 ( .A(n226), .B(n501), .S(n533), .Z(n228) );
  NR2 U47 ( .A(n501), .B(n461), .Z(n226) );
  EO U48 ( .A(n526), .B(n501), .Z(n111) );
  ND2 U49 ( .A(n503), .B(n464), .Z(n108) );
  NR2 U50 ( .A(n531), .B(n467), .Z(n273) );
  AO4 U51 ( .A(n502), .B(n463), .C(n534), .D(n462), .Z(n92) );
  EN U52 ( .A(n527), .B(n499), .Z(n97) );
  EN U53 ( .A(n527), .B(n500), .Z(n96) );
  ND2 U54 ( .A(n307), .B(n306), .Z(n102) );
  EN U55 ( .A(n527), .B(n469), .Z(n307) );
  ND2 U56 ( .A(n496), .B(n469), .Z(n306) );
  ND2 U57 ( .A(n503), .B(n464), .Z(n90) );
  EO U58 ( .A(n527), .B(n470), .Z(n103) );
  EO U59 ( .A(n527), .B(n470), .Z(n104) );
  EO U60 ( .A(n527), .B(n461), .Z(n105) );
  AO4 U61 ( .A(n501), .B(n462), .C(n533), .D(n462), .Z(n78) );
  EO U62 ( .A(n495), .B(n466), .Z(n81) );
  ND2 U63 ( .A(n533), .B(n502), .Z(n209) );
  ND2 U64 ( .A(n280), .B(n279), .Z(n68) );
  EN U65 ( .A(n495), .B(n467), .Z(n280) );
  EN U66 ( .A(n527), .B(n467), .Z(n279) );
  ND2 U67 ( .A(n500), .B(n466), .Z(n254) );
  ND2 U68 ( .A(n532), .B(n465), .Z(n255) );
  AO4 U69 ( .A(n498), .B(n468), .C(n530), .D(n468), .Z(n69) );
  AO7 U70 ( .A(n529), .B(n497), .C(n470), .Z(n72) );
  ND2 U71 ( .A(n351), .B(n350), .Z(n74) );
  ND2 U72 ( .A(n503), .B(n460), .Z(n350) );
  ND2 U73 ( .A(n530), .B(n460), .Z(n351) );
  ND2 U74 ( .A(n309), .B(n308), .Z(n70) );
  ND2 U75 ( .A(n529), .B(n469), .Z(n309) );
  ND2 U76 ( .A(n497), .B(n469), .Z(n308) );
  AN2P U77 ( .A(n498), .B(n467), .Z(n42) );
  MUX21L U78 ( .A(n461), .B(n331), .S(n497), .Z(n73) );
  ND2 U79 ( .A(n527), .B(n461), .Z(n331) );
  AN3 U80 ( .A(n495), .B(n460), .C(n526), .Z(n59) );
  ND2 U81 ( .A(n529), .B(n470), .Z(n324) );
  ND2 U82 ( .A(n498), .B(n470), .Z(n323) );
  AO4 U83 ( .A(n497), .B(n468), .C(n530), .D(n468), .Z(n51) );
  ND2 U84 ( .A(n499), .B(n466), .Z(n260) );
  AN2P U85 ( .A(n503), .B(n464), .Z(n43) );
  IVP U86 ( .A(n442), .Z(n466) );
  IVP U87 ( .A(n442), .Z(n463) );
  IVP U88 ( .A(n442), .Z(n467) );
  ND2 U89 ( .A(n259), .B(n518), .Z(n172) );
  EO U90 ( .A(n495), .B(n466), .Z(n259) );
  ND2 U91 ( .A(n190), .B(n189), .Z(n149) );
  MUX21L U92 ( .A(n187), .B(n188), .S(n503), .Z(n190) );
  ND2 U93 ( .A(n186), .B(n523), .Z(n189) );
  NR2 U94 ( .A(n534), .B(n450), .Z(n188) );
  ND2 U95 ( .A(n268), .B(n267), .Z(n158) );
  ND2 U96 ( .A(n467), .B(n516), .Z(n267) );
  EN U97 ( .A(n495), .B(n467), .Z(n268) );
  IVP U98 ( .A(n441), .Z(n460) );
  IVP U99 ( .A(n442), .Z(n465) );
  IVP U100 ( .A(n477), .Z(n500) );
  IVP U101 ( .A(n510), .Z(n531) );
  IVP U102 ( .A(n476), .Z(n497) );
  IVP U103 ( .A(n510), .Z(n533) );
  IVP U104 ( .A(n477), .Z(n502) );
  IVP U105 ( .A(n510), .Z(n532) );
  IVP U106 ( .A(n442), .Z(n464) );
  IVP U107 ( .A(n477), .Z(n503) );
  IVP U108 ( .A(n476), .Z(n496) );
  IVP U109 ( .A(n509), .Z(n527) );
  IVP U110 ( .A(n510), .Z(n530) );
  IVP U111 ( .A(n476), .Z(n495) );
  IVP U112 ( .A(n510), .Z(n534) );
  IVP U113 ( .A(n442), .Z(n468) );
  AO7 U114 ( .A(n499), .B(n524), .C(n465), .Z(n165) );
  ND3 U115 ( .A(n248), .B(n247), .C(n246), .Z(n171) );
  ND2 U116 ( .A(n452), .B(n488), .Z(n247) );
  ND2 U117 ( .A(n532), .B(n488), .Z(n248) );
  ND2 U118 ( .A(n532), .B(n452), .Z(n246) );
  ND2 U119 ( .A(n233), .B(n232), .Z(n170) );
  MUX21L U120 ( .A(n230), .B(n231), .S(n464), .Z(n233) );
  ND2 U121 ( .A(n229), .B(n533), .Z(n232) );
  NR2 U122 ( .A(n533), .B(n489), .Z(n230) );
  ND2 U123 ( .A(n201), .B(n200), .Z(n167) );
  ND2 U124 ( .A(n502), .B(n522), .Z(n200) );
  MUX21L U125 ( .A(n522), .B(n199), .S(n463), .Z(n201) );
  NR2 U126 ( .A(n502), .B(n522), .Z(n199) );
  ND2 U127 ( .A(n212), .B(n211), .Z(n168) );
  ND2 U128 ( .A(n502), .B(n520), .Z(n211) );
  MUX21L U129 ( .A(n521), .B(n210), .S(n463), .Z(n212) );
  NR2 U130 ( .A(n502), .B(n520), .Z(n210) );
  ND2 U149 ( .A(n314), .B(n313), .Z(n177) );
  ND2 U150 ( .A(n310), .B(n512), .Z(n313) );
  MUX21L U151 ( .A(n311), .B(n312), .S(n496), .Z(n314) );
  NR2 U152 ( .A(n470), .B(n497), .Z(n310) );
  ND2 U153 ( .A(n250), .B(n249), .Z(n154) );
  ND2 U154 ( .A(n453), .B(n488), .Z(n249) );
  EN U155 ( .A(n527), .B(n500), .Z(n250) );
  ND2 U156 ( .A(n444), .B(n511), .Z(n338) );
  MUX21L U157 ( .A(n478), .B(n337), .S(n461), .Z(n339) );
  MUX21L U158 ( .A(n194), .B(n450), .S(n534), .Z(n166) );
  ND2 U159 ( .A(n450), .B(n492), .Z(n194) );
  MUX21L U160 ( .A(n282), .B(n281), .S(n498), .Z(n175) );
  ND2 U161 ( .A(n531), .B(n457), .Z(n282) );
  ND2 U162 ( .A(n530), .B(n467), .Z(n281) );
  MUX21L U178 ( .A(n214), .B(n213), .S(n502), .Z(n151) );
  ND2 U179 ( .A(n448), .B(n520), .Z(n213) );
  ND2 U180 ( .A(n533), .B(n448), .Z(n214) );
  MUX21L U181 ( .A(n486), .B(n517), .S(n466), .Z(n157) );
  MUX21L U182 ( .A(n514), .B(n484), .S(n468), .Z(n159) );
  IVP U183 ( .A(n509), .Z(n529) );
  IVP U184 ( .A(n509), .Z(n528) );
  IVP U185 ( .A(n443), .Z(n470) );
  IVP U186 ( .A(n441), .Z(n462) );
  IVP U187 ( .A(n476), .Z(n498) );
  IVP U188 ( .A(n476), .Z(n499) );
  AO7 U189 ( .A(n533), .B(n490), .C(n445), .Z(n169) );
  AO7 U190 ( .A(n499), .B(n517), .C(n455), .Z(n155) );
  NR2 U191 ( .A(n529), .B(n459), .Z(n312) );
  NR2 U192 ( .A(n532), .B(n489), .Z(n236) );
  ND2 U193 ( .A(n531), .B(n456), .Z(n174) );
  ND2 U194 ( .A(n238), .B(n237), .Z(n140) );
  ND2 U195 ( .A(n234), .B(n519), .Z(n237) );
  MUX21L U196 ( .A(n235), .B(n236), .S(n465), .Z(n238) );
  NR2 U197 ( .A(n465), .B(n500), .Z(n234) );
  ND2 U198 ( .A(n197), .B(n196), .Z(n136) );
  ND2 U199 ( .A(n463), .B(n492), .Z(n196) );
  MUX21L U200 ( .A(n195), .B(n534), .S(n463), .Z(n197) );
  NR2 U201 ( .A(n534), .B(n492), .Z(n195) );
  ND2 U202 ( .A(n183), .B(n182), .Z(n135) );
  ND2 U203 ( .A(n464), .B(n494), .Z(n182) );
  MUX21L U204 ( .A(n494), .B(n181), .S(n534), .Z(n183) );
  NR2 U205 ( .A(n464), .B(n494), .Z(n181) );
  ND2 U206 ( .A(n218), .B(n447), .Z(n138) );
  ND2 U207 ( .A(n533), .B(n501), .Z(n218) );
  MUX21L U208 ( .A(n490), .B(n519), .S(n462), .Z(n152) );
  MUX21L U209 ( .A(n205), .B(n204), .S(n534), .Z(n137) );
  ND2 U210 ( .A(n462), .B(n491), .Z(n205) );
  ND2 U211 ( .A(n502), .B(n462), .Z(n204) );
  IVP U212 ( .A(n441), .Z(n461) );
  IVP U213 ( .A(n443), .Z(n469) );
  IVP U214 ( .A(n477), .Z(n501) );
  ND2 U215 ( .A(n469), .B(n484), .Z(n300) );
  ND2 U216 ( .A(n469), .B(n513), .Z(n299) );
  ND2 U217 ( .A(n463), .B(n493), .Z(n192) );
  MUX21L U218 ( .A(n493), .B(n191), .S(n534), .Z(n193) );
  NR2 U219 ( .A(n463), .B(n493), .Z(n191) );
  ND2 U220 ( .A(n185), .B(n184), .Z(n122) );
  ND2 U221 ( .A(n534), .B(n451), .Z(n184) );
  EN U222 ( .A(n495), .B(n464), .Z(n185) );
  MUX21L U223 ( .A(n463), .B(n202), .S(n534), .Z(n124) );
  ND2 U224 ( .A(n463), .B(n491), .Z(n202) );
  ND2 U225 ( .A(n501), .B(n446), .Z(n222) );
  ND2 U226 ( .A(n341), .B(n340), .Z(n133) );
  ND2 U227 ( .A(n496), .B(n444), .Z(n340) );
  EO U228 ( .A(n526), .B(n460), .Z(n341) );
  MUX21L U229 ( .A(n283), .B(n498), .S(n467), .Z(n130) );
  ND2 U230 ( .A(n497), .B(n515), .Z(n283) );
  AO7 U231 ( .A(n531), .B(n498), .C(n456), .Z(n128) );
  ND2 U232 ( .A(n455), .B(n487), .Z(n142) );
  ND2 U233 ( .A(n452), .B(n518), .Z(n244) );
  ND2 U234 ( .A(n287), .B(n286), .Z(n117) );
  MUX21L U235 ( .A(n284), .B(n515), .S(n497), .Z(n286) );
  AO6 U236 ( .A(n499), .B(n457), .C(n285), .Z(n287) );
  ND2 U237 ( .A(n305), .B(n304), .Z(n118) );
  ND2 U238 ( .A(n483), .B(n513), .Z(n304) );
  MUX21L U239 ( .A(n483), .B(n303), .S(n469), .Z(n305) );
  ND2 U240 ( .A(n271), .B(n270), .Z(n116) );
  ND2 U241 ( .A(n531), .B(n456), .Z(n270) );
  MUX21L U242 ( .A(n486), .B(n269), .S(n467), .Z(n271) );
  NR2 U243 ( .A(n531), .B(n486), .Z(n269) );
  ND2 U244 ( .A(n241), .B(n240), .Z(n113) );
  ND2 U245 ( .A(n532), .B(n489), .Z(n240) );
  MUX21L U246 ( .A(n239), .B(n451), .S(n532), .Z(n241) );
  ND2 U247 ( .A(n208), .B(n207), .Z(n110) );
  MUX21L U248 ( .A(n206), .B(n521), .S(n502), .Z(n208) );
  ND2 U249 ( .A(n463), .B(n502), .Z(n207) );
  NR2 U250 ( .A(n462), .B(n521), .Z(n206) );
  MUX21L U251 ( .A(n325), .B(n527), .S(n461), .Z(n132) );
  ND2 U252 ( .A(n529), .B(n480), .Z(n325) );
  AO7 U253 ( .A(n499), .B(n466), .C(n517), .Z(n115) );
  ND2 U254 ( .A(n344), .B(n343), .Z(n120) );
  ND2 U255 ( .A(n528), .B(n495), .Z(n343) );
  MUX21L U256 ( .A(n342), .B(n444), .S(n495), .Z(n344) );
  NR2 U257 ( .A(n528), .B(n443), .Z(n342) );
  MUX21L U258 ( .A(n198), .B(n449), .S(n502), .Z(n109) );
  ND2 U259 ( .A(n449), .B(n523), .Z(n198) );
  ND2 U260 ( .A(n275), .B(n274), .Z(n100) );
  MUX21L U261 ( .A(n272), .B(n516), .S(n498), .Z(n274) );
  AO6 U262 ( .A(n498), .B(n457), .C(n273), .Z(n275) );
  ND2 U263 ( .A(n327), .B(n326), .Z(n119) );
  ND2 U264 ( .A(n480), .B(n512), .Z(n327) );
  ND2 U265 ( .A(n461), .B(n480), .Z(n326) );
  AO7 U266 ( .A(n532), .B(n451), .C(n500), .Z(n95) );
  NR2 U267 ( .A(n468), .B(n485), .Z(n291) );
  NR2 U268 ( .A(n497), .B(n514), .Z(n292) );
  NR2 U269 ( .A(n528), .B(n477), .Z(n346) );
  ND2 U270 ( .A(n295), .B(n294), .Z(n101) );
  NR2 U271 ( .A(n293), .B(n292), .Z(n295) );
  MUX21L U272 ( .A(n291), .B(n468), .S(n530), .Z(n294) );
  NR2 U273 ( .A(n498), .B(n458), .Z(n293) );
  ND2 U274 ( .A(n263), .B(n262), .Z(n99) );
  ND2 U275 ( .A(n531), .B(n487), .Z(n263) );
  ND2 U276 ( .A(n466), .B(n487), .Z(n262) );
  ND2 U277 ( .A(n349), .B(n348), .Z(n106) );
  NR2 U278 ( .A(n347), .B(n346), .Z(n349) );
  MUX21L U279 ( .A(n345), .B(n460), .S(n496), .Z(n348) );
  NR2 U280 ( .A(n527), .B(n443), .Z(n347) );
  ND2 U281 ( .A(n217), .B(n216), .Z(n93) );
  ND2 U282 ( .A(n447), .B(n519), .Z(n216) );
  MUX21L U283 ( .A(n490), .B(n215), .S(n462), .Z(n217) );
  ND2 U284 ( .A(n221), .B(n220), .Z(n94) );
  ND2 U285 ( .A(n501), .B(n446), .Z(n220) );
  ND2 U286 ( .A(n533), .B(n446), .Z(n221) );
  NR2 U287 ( .A(n460), .B(n511), .Z(n345) );
  NR2 U288 ( .A(n499), .B(n454), .Z(n256) );
  ND2 U289 ( .A(n465), .B(n518), .Z(n242) );
  EN U290 ( .A(n495), .B(n465), .Z(n243) );
  ND2 U291 ( .A(n499), .B(n454), .Z(n257) );
  MUX21L U292 ( .A(n256), .B(n455), .S(n531), .Z(n258) );
  ND2 U293 ( .A(n253), .B(n252), .Z(n79) );
  ND2 U294 ( .A(n500), .B(n453), .Z(n252) );
  MUX21L U295 ( .A(n251), .B(n454), .S(n532), .Z(n253) );
  NR2 U296 ( .A(n500), .B(n453), .Z(n251) );
  ND3 U297 ( .A(n278), .B(n277), .C(n276), .Z(n82) );
  ND2 U298 ( .A(n485), .B(n515), .Z(n277) );
  ND2 U299 ( .A(n467), .B(n516), .Z(n278) );
  ND2 U300 ( .A(n467), .B(n485), .Z(n276) );
  ND2 U301 ( .A(n297), .B(n296), .Z(n83) );
  ND2 U302 ( .A(n458), .B(n514), .Z(n296) );
  EO U303 ( .A(n495), .B(n469), .Z(n297) );
  ND2 U304 ( .A(n322), .B(n321), .Z(n86) );
  ND2 U305 ( .A(n530), .B(n496), .Z(n321) );
  MUX21L U306 ( .A(n320), .B(n459), .S(n496), .Z(n322) );
  NR2 U307 ( .A(n528), .B(n459), .Z(n320) );
  ND3 U308 ( .A(n491), .B(n523), .C(n449), .Z(n91) );
  ND2 U309 ( .A(n317), .B(n316), .Z(n85) );
  ND2 U310 ( .A(n528), .B(n482), .Z(n316) );
  MUX21L U311 ( .A(n482), .B(n315), .S(n470), .Z(n317) );
  NR2 U312 ( .A(n529), .B(n481), .Z(n315) );
  ND2 U313 ( .A(n330), .B(n329), .Z(n87) );
  ND2 U314 ( .A(n528), .B(n479), .Z(n329) );
  MUX21L U315 ( .A(n479), .B(n328), .S(n462), .Z(n330) );
  NR2 U316 ( .A(n528), .B(n479), .Z(n328) );
  MUX21L U317 ( .A(n336), .B(n335), .S(n461), .Z(n88) );
  ND2 U318 ( .A(n478), .B(n511), .Z(n335) );
  ND2 U319 ( .A(n528), .B(n496), .Z(n336) );
  MUX21L U320 ( .A(n483), .B(n301), .S(n469), .Z(n84) );
  ND2 U321 ( .A(n484), .B(n513), .Z(n301) );
  ND2 U322 ( .A(n219), .B(n447), .Z(n64) );
  ND2 U323 ( .A(n533), .B(n501), .Z(n219) );
  ND2 U324 ( .A(n319), .B(n318), .Z(n71) );
  ND2 U325 ( .A(n470), .B(n512), .Z(n318) );
  EN U326 ( .A(n495), .B(n470), .Z(n319) );
  MUX21L U327 ( .A(n49), .B(n48), .S(n432), .Z(n409) );
  ND2 U328 ( .A(n503), .B(n464), .Z(n48) );
  ND2 U329 ( .A(n261), .B(n260), .Z(n49) );
  ND2 U330 ( .A(n531), .B(n466), .Z(n261) );
  ND2 U331 ( .A(n431), .B(n43), .Z(n353) );
  MUX21L U332 ( .A(n417), .B(n416), .S(n435), .Z(n419) );
  AN3 U333 ( .A(n431), .B(n145), .C(n438), .Z(n417) );
  ND2 U334 ( .A(n290), .B(n289), .Z(n145) );
  MUX21L U335 ( .A(n413), .B(n412), .S(n432), .Z(n421) );
  NR3 U336 ( .A(n438), .B(n36), .C(n434), .Z(n412) );
  NR2 U337 ( .A(n438), .B(n34), .Z(n413) );
  MUX21L U338 ( .A(n415), .B(n414), .S(n438), .Z(n420) );
  NR2 U339 ( .A(n432), .B(n423), .Z(n414) );
  IVP U340 ( .A(n146), .Z(n423) );
  IVP U341 ( .A(n428), .Z(n431) );
  IVP U342 ( .A(n427), .Z(n430) );
  MUX21L U343 ( .A(n367), .B(n366), .S(n431), .Z(n370) );
  AN3 U344 ( .A(n125), .B(n434), .C(n438), .Z(n367) );
  AN3 U345 ( .A(n122), .B(n434), .C(n438), .Z(n366) );
  MUX21L U346 ( .A(n222), .B(n445), .S(n533), .Z(n125) );
  IVP U347 ( .A(n429), .Z(n432) );
  ND2 U348 ( .A(n434), .B(n426), .Z(n418) );
  AO2 U349 ( .A(n398), .B(n435), .C(n397), .D(n435), .Z(n406) );
  NR2 U350 ( .A(n439), .B(n427), .Z(n397) );
  NR2 U351 ( .A(n439), .B(n37), .Z(n398) );
  MUX21L U352 ( .A(n399), .B(n400), .S(n432), .Z(n408) );
  NR2 U353 ( .A(n439), .B(n422), .Z(n400) );
  NR3 U354 ( .A(n439), .B(n38), .C(n435), .Z(n399) );
  IVP U355 ( .A(n78), .Z(n422) );
  MUX21L U356 ( .A(n404), .B(n403), .S(n432), .Z(n405) );
  AN3 U357 ( .A(n438), .B(n460), .C(n434), .Z(n404) );
  ND2 U358 ( .A(n503), .B(n464), .Z(n76) );
  MUX21L U359 ( .A(n358), .B(n359), .S(n435), .Z(n361) );
  NR2 U360 ( .A(n439), .B(n429), .Z(n359) );
  ND2 U361 ( .A(n255), .B(n254), .Z(n65) );
  MUX21L U362 ( .A(n354), .B(n355), .S(n435), .Z(n363) );
  NR2 U363 ( .A(n439), .B(n59), .Z(n355) );
  MUX21L U364 ( .A(n356), .B(n357), .S(n435), .Z(n362) );
  ND2 U365 ( .A(n503), .B(n464), .Z(n63) );
  MUX21L U366 ( .A(n389), .B(n390), .S(n435), .Z(n395) );
  AN3 U367 ( .A(n61), .B(n426), .C(n438), .Z(n389) );
  ND2 U368 ( .A(n445), .B(n478), .Z(n61) );
  MUX21L U369 ( .A(n387), .B(n388), .S(n435), .Z(n396) );
  NR2 U370 ( .A(n439), .B(n427), .Z(n387) );
  AN3 U371 ( .A(n495), .B(n460), .C(n527), .Z(n57) );
  MUX21L U372 ( .A(n391), .B(n392), .S(n435), .Z(n394) );
  AO4 U373 ( .A(n498), .B(n468), .C(n530), .D(n468), .Z(n58) );
  MUX21L U374 ( .A(n373), .B(n53), .S(n431), .Z(n378) );
  ND2 U375 ( .A(n503), .B(n464), .Z(n53) );
  MUX21L U376 ( .A(n381), .B(n382), .S(n435), .Z(n383) );
  NR2 U377 ( .A(n432), .B(n39), .Z(n382) );
  EN U378 ( .A(n438), .B(n432), .Z(n410) );
  EN U379 ( .A(n434), .B(n432), .Z(n411) );
  ND2 U380 ( .A(n46), .B(n439), .Z(n386) );
  ND2 U381 ( .A(n298), .B(n458), .Z(n46) );
  ND2 U382 ( .A(n529), .B(n497), .Z(n298) );
  MUX21L U383 ( .A(n379), .B(n380), .S(n432), .Z(n384) );
  NR2 U384 ( .A(n439), .B(n435), .Z(n380) );
  ND2 U385 ( .A(n435), .B(n431), .Z(n385) );
  ND2 U386 ( .A(n440), .B(n435), .Z(n352) );
  NR2 U387 ( .A(n470), .B(n481), .Z(n178) );
  IVP U388 ( .A(n471), .Z(n472) );
  ND4 U389 ( .A(n421), .B(n420), .C(n419), .D(n418), .Z(n147) );
  IVP U390 ( .A(n504), .Z(n505) );
  ND3 U391 ( .A(n372), .B(n371), .C(n370), .Z(n127) );
  IVP U392 ( .A(n444), .Z(n474) );
  IVP U393 ( .A(n448), .Z(n475) );
  IVP U394 ( .A(n478), .Z(n507) );
  IVP U395 ( .A(n471), .Z(n473) );
  MUX21L U396 ( .A(n368), .B(n369), .S(n431), .Z(n371) );
  NR3 U397 ( .A(n439), .B(n534), .C(n435), .Z(n369) );
  AN3 U398 ( .A(n126), .B(n437), .C(n434), .Z(n368) );
  ND2 U399 ( .A(n245), .B(n244), .Z(n126) );
  MUX21L U400 ( .A(n364), .B(n365), .S(n435), .Z(n372) );
  AN3 U401 ( .A(n123), .B(n437), .C(n430), .Z(n365) );
  AN3 U402 ( .A(n124), .B(n430), .C(n438), .Z(n364) );
  ND2 U403 ( .A(n193), .B(n192), .Z(n123) );
  IVP U404 ( .A(n433), .Z(n436) );
  IVP U405 ( .A(n433), .Z(n434) );
  IVP U406 ( .A(n504), .Z(n506) );
  IVP U407 ( .A(n479), .Z(n508) );
  IVP U408 ( .A(n433), .Z(n435) );
  IVP U409 ( .A(n437), .Z(n440) );
  IVP U410 ( .A(n437), .Z(n438) );
  IVP U411 ( .A(n437), .Z(n439) );
  ND4 U412 ( .A(n408), .B(n407), .C(n406), .D(n405), .Z(n80) );
  MUX21L U413 ( .A(n402), .B(n401), .S(n432), .Z(n407) );
  AN3 U414 ( .A(n77), .B(n433), .C(n438), .Z(n401) );
  AN3 U415 ( .A(n79), .B(n433), .C(n438), .Z(n402) );
  ND2 U416 ( .A(n209), .B(n448), .Z(n77) );
  ND4 U417 ( .A(n363), .B(n362), .C(n361), .D(n360), .Z(n67) );
  ND4 U418 ( .A(n66), .B(n428), .C(n433), .D(n437), .Z(n360) );
  AO7 U419 ( .A(n531), .B(n499), .C(n466), .Z(n66) );
  ND4 U420 ( .A(n396), .B(n395), .C(n394), .D(n393), .Z(n62) );
  ND4 U421 ( .A(n378), .B(n377), .C(n376), .D(n375), .Z(n56) );
  ND3 U422 ( .A(n55), .B(n437), .C(n433), .Z(n375) );
  AO7 U423 ( .A(n531), .B(n499), .C(n466), .Z(n55) );
  MUX21L U424 ( .A(n374), .B(n437), .S(n432), .Z(n377) );
  AN3 U425 ( .A(n495), .B(n460), .C(n526), .Z(n54) );
  ND4 U426 ( .A(n60), .B(n435), .C(n428), .D(n437), .Z(n393) );
  AO7 U427 ( .A(n528), .B(n496), .C(n470), .Z(n60) );
  ND3 U428 ( .A(n411), .B(n410), .C(n409), .Z(n50) );
  ND2 U429 ( .A(n384), .B(n383), .Z(n52) );
  ND2 U430 ( .A(n431), .B(n433), .Z(n376) );
  AO7 U431 ( .A(n429), .B(n386), .C(n385), .Z(n47) );
  ND4 U432 ( .A(n439), .B(n435), .C(n432), .D(n43), .Z(n45) );
  NR2 U433 ( .A(n353), .B(n352), .Z(n44) );
  IVP U434 ( .A(n424), .Z(n425) );
  EN U435 ( .A(n547), .B(x[15]), .Z(N57) );
  ND2 U436 ( .A(x[14]), .B(func), .Z(n547) );
  IVP U437 ( .A(reset), .Z(n544) );
  MUX21H U438 ( .A(n47), .B(n45), .S(n425), .Z(N9) );
  MUX21H U439 ( .A(n52), .B(n50), .S(n425), .Z(N10) );
  MUX21H U440 ( .A(n62), .B(n56), .S(n425), .Z(N11) );
  MUX81P U441 ( .D0(n74), .D1(n70), .D2(n72), .D3(n68), .D4(n73), .D5(n69), 
        .D6(n71), .D7(n42), .A(n431), .B(n436), .C(n439), .Z(n75) );
  MUX21H U442 ( .A(n75), .B(n67), .S(n425), .Z(N12) );
  MUX81P U443 ( .D0(n88), .D1(n84), .D2(n86), .D3(n82), .D4(n87), .D5(n83), 
        .D6(n85), .D7(n81), .A(n431), .B(n436), .C(n440), .Z(n89) );
  MUX21H U444 ( .A(n89), .B(n80), .S(n425), .Z(N13) );
  MUX81P U445 ( .D0(n97), .D1(n93), .D2(n95), .D3(n91), .D4(n96), .D5(n92), 
        .D6(n94), .D7(n90), .A(n431), .B(n436), .C(n440), .Z(n98) );
  MUX81P U446 ( .D0(n106), .D1(n102), .D2(n104), .D3(n100), .D4(n105), .D5(
        n101), .D6(n103), .D7(n99), .A(n431), .B(n436), .C(n440), .Z(n107) );
  MUX21H U447 ( .A(n107), .B(n98), .S(n425), .Z(N14) );
  MUX81P U448 ( .D0(n524), .D1(n111), .D2(n113), .D3(n109), .D4(n524), .D5(
        n110), .D6(n112), .D7(n108), .A(n431), .B(n436), .C(n440), .Z(n114) );
  MUX81P U449 ( .D0(n120), .D1(n118), .D2(n481), .D3(n116), .D4(n119), .D5(
        n117), .D6(n482), .D7(n115), .A(n431), .B(n436), .C(n440), .Z(n121) );
  MUX21H U450 ( .A(n121), .B(n114), .S(n425), .Z(N15) );
  MUX81P U451 ( .D0(n133), .D1(n131), .D2(n525), .D3(n129), .D4(n132), .D5(
        n130), .D6(n525), .D7(n128), .A(n431), .B(n436), .C(n440), .Z(n134) );
  MUX21H U452 ( .A(n134), .B(n127), .S(n425), .Z(N16) );
  MUX81P U453 ( .D0(n142), .D1(n138), .D2(n140), .D3(n136), .D4(n141), .D5(
        n137), .D6(n139), .D7(n135), .A(n431), .B(n436), .C(n440), .Z(n143) );
  MUX21H U454 ( .A(n147), .B(n143), .S(n425), .Z(N17) );
  MUX81P U455 ( .D0(n155), .D1(n151), .D2(n153), .D3(n149), .D4(n154), .D5(
        n150), .D6(n152), .D7(n148), .A(n431), .B(n436), .C(n440), .Z(n156) );
  MUX81P U456 ( .D0(n163), .D1(n160), .D2(n465), .D3(n158), .D4(n162), .D5(
        n159), .D6(n161), .D7(n157), .A(n431), .B(n436), .C(n440), .Z(n164) );
  MUX21H U457 ( .A(n164), .B(n156), .S(n425), .Z(N18) );
  MUX81P U458 ( .D0(n172), .D1(n168), .D2(n170), .D3(n166), .D4(n171), .D5(
        n167), .D6(n169), .D7(n165), .A(n431), .B(n436), .C(n440), .Z(n173) );
  MUX81P U459 ( .D0(n525), .D1(n176), .D2(n178), .D3(n175), .D4(n179), .D5(n41), .D6(n177), .D7(n174), .A(n430), .B(n436), .C(n440), .Z(n180) );
  MUX21H U460 ( .A(n180), .B(n173), .S(n425), .Z(N19) );
  AN2P U461 ( .A(n526), .B(n460), .Z(n187) );
  AN2P U462 ( .A(n527), .B(n495), .Z(n215) );
  AN2P U463 ( .A(n527), .B(n495), .Z(n235) );
  AN2P U464 ( .A(n495), .B(n460), .Z(n239) );
  AN2P U465 ( .A(n527), .B(n460), .Z(n272) );
  AN2P U466 ( .A(n527), .B(n460), .Z(n284) );
  AN2P U467 ( .A(n527), .B(n495), .Z(n303) );
  AN2P U468 ( .A(n526), .B(n460), .Z(n311) );
  AN2P U469 ( .A(n526), .B(n495), .Z(n337) );
  AN2P U470 ( .A(n438), .B(n430), .Z(n354) );
  AN2P U471 ( .A(n64), .B(n430), .Z(n356) );
  AN2P U472 ( .A(n63), .B(n430), .Z(n357) );
  AN2P U473 ( .A(n438), .B(n65), .Z(n358) );
  AN2P U474 ( .A(n438), .B(n434), .Z(n373) );
  AN2P U475 ( .A(n434), .B(n54), .Z(n374) );
  AN2P U476 ( .A(n438), .B(n434), .Z(n379) );
  AN2P U477 ( .A(n430), .B(n51), .Z(n381) );
  AN2P U478 ( .A(n57), .B(n430), .Z(n388) );
  AN2P U479 ( .A(n59), .B(n438), .Z(n390) );
  AN2P U480 ( .A(n58), .B(n430), .Z(n391) );
  AN2P U481 ( .A(n438), .B(n430), .Z(n392) );
  AN2P U482 ( .A(n76), .B(n434), .Z(n403) );
  AN2P U483 ( .A(n510), .B(n434), .Z(n415) );
  AN2P U484 ( .A(n144), .B(n438), .Z(n416) );
  IV U485 ( .A(x[14]), .Z(n424) );
  IVA U486 ( .A(n542), .Z(n426) );
  IVA U487 ( .A(n542), .Z(n427) );
  IVA U488 ( .A(n542), .Z(n428) );
  IVA U489 ( .A(n542), .Z(n429) );
  IVP U490 ( .A(x[12]), .Z(n433) );
  IVA U491 ( .A(x[11]), .Z(n437) );
  IVA U492 ( .A(n472), .Z(n441) );
  IVA U493 ( .A(n472), .Z(n442) );
  IVA U494 ( .A(n472), .Z(n443) );
  IVA U495 ( .A(n472), .Z(n444) );
  IVA U496 ( .A(n473), .Z(n445) );
  IVA U497 ( .A(n473), .Z(n446) );
  IVA U498 ( .A(n473), .Z(n447) );
  IVA U499 ( .A(n473), .Z(n448) );
  IVA U500 ( .A(n473), .Z(n449) );
  IVA U501 ( .A(n474), .Z(n450) );
  IVA U502 ( .A(n474), .Z(n451) );
  IVA U503 ( .A(n474), .Z(n452) );
  IVA U504 ( .A(n474), .Z(n453) );
  IVA U505 ( .A(n474), .Z(n454) );
  IVA U506 ( .A(n475), .Z(n455) );
  IVA U507 ( .A(n475), .Z(n456) );
  IVA U508 ( .A(n475), .Z(n457) );
  IVA U509 ( .A(n475), .Z(n458) );
  IVA U510 ( .A(n475), .Z(n459) );
  IVP U511 ( .A(x[10]), .Z(n471) );
  IVA U512 ( .A(n505), .Z(n476) );
  IVA U513 ( .A(n505), .Z(n477) );
  IVA U514 ( .A(n505), .Z(n478) );
  IVA U515 ( .A(n505), .Z(n479) );
  IVA U516 ( .A(n506), .Z(n480) );
  IVA U517 ( .A(n506), .Z(n481) );
  IVA U518 ( .A(n506), .Z(n482) );
  IVA U519 ( .A(n506), .Z(n483) );
  IVA U520 ( .A(n506), .Z(n484) );
  IVA U521 ( .A(n507), .Z(n485) );
  IVA U522 ( .A(n507), .Z(n486) );
  IVA U523 ( .A(n507), .Z(n487) );
  IVA U524 ( .A(n507), .Z(n488) );
  IVA U525 ( .A(n507), .Z(n489) );
  IVA U526 ( .A(n508), .Z(n490) );
  IVA U527 ( .A(n508), .Z(n491) );
  IVA U528 ( .A(n508), .Z(n492) );
  IVA U529 ( .A(n508), .Z(n493) );
  IVA U530 ( .A(n508), .Z(n494) );
  IVP U531 ( .A(x[9]), .Z(n504) );
  IVA U532 ( .A(n536), .Z(n509) );
  IVA U533 ( .A(n536), .Z(n510) );
  IVA U534 ( .A(n537), .Z(n511) );
  IVA U535 ( .A(n537), .Z(n512) );
  IVA U536 ( .A(n537), .Z(n513) );
  IVA U537 ( .A(n538), .Z(n514) );
  IVA U538 ( .A(n538), .Z(n515) );
  IVA U539 ( .A(n538), .Z(n516) );
  IVA U540 ( .A(n539), .Z(n517) );
  IVA U541 ( .A(n539), .Z(n518) );
  IVA U542 ( .A(n539), .Z(n519) );
  IVA U543 ( .A(n540), .Z(n520) );
  IVA U544 ( .A(n540), .Z(n521) );
  IVA U545 ( .A(n540), .Z(n522) );
  IVA U546 ( .A(n541), .Z(n523) );
  IVA U547 ( .A(n541), .Z(n524) );
  IVA U548 ( .A(n541), .Z(n525) );
  IV U549 ( .A(n509), .Z(n526) );
  IVA U550 ( .A(x[8]), .Z(n535) );
  IVA U551 ( .A(n535), .Z(n536) );
  IVA U552 ( .A(n535), .Z(n537) );
  IVA U553 ( .A(n535), .Z(n538) );
  IVA U554 ( .A(n511), .Z(n539) );
  IVA U555 ( .A(n513), .Z(n540) );
  IVA U556 ( .A(n512), .Z(n541) );
  IVA U557 ( .A(n543), .Z(n542) );
  IV U558 ( .A(x[13]), .Z(n543) );
  EO U559 ( .A(Term1[25]), .B(\add_1242/carry[14] ), .Z(N50) );
  AN2 U560 ( .A(\add_1242/carry[13] ), .B(Term1[24]), .Z(\add_1242/carry[14] )
         );
  EO U561 ( .A(Term1[24]), .B(\add_1242/carry[13] ), .Z(N49) );
  AN2 U562 ( .A(\add_1242/carry[12] ), .B(Term1[23]), .Z(\add_1242/carry[13] )
         );
  EO U563 ( .A(Term1[23]), .B(\add_1242/carry[12] ), .Z(N48) );
  AN2 U564 ( .A(\add_1242/carry[11] ), .B(Term1[22]), .Z(\add_1242/carry[12] )
         );
  EO U565 ( .A(Term1[22]), .B(\add_1242/carry[11] ), .Z(N47) );
  AN2 U566 ( .A(\add_1242/carry[10] ), .B(Term1[21]), .Z(\add_1242/carry[11] )
         );
  EO U567 ( .A(Term1[21]), .B(\add_1242/carry[10] ), .Z(N46) );
  AN2 U568 ( .A(\add_1242/carry[9] ), .B(Term1[20]), .Z(\add_1242/carry[10] )
         );
  EO U569 ( .A(Term1[20]), .B(\add_1242/carry[9] ), .Z(N45) );
  AN2 U570 ( .A(\add_1242/carry[8] ), .B(Term1[19]), .Z(\add_1242/carry[9] )
         );
  EO U571 ( .A(Term1[19]), .B(\add_1242/carry[8] ), .Z(N44) );
  AN2 U572 ( .A(\add_1242/carry[7] ), .B(Term1[18]), .Z(\add_1242/carry[8] )
         );
  EO U573 ( .A(Term1[18]), .B(\add_1242/carry[7] ), .Z(N43) );
  AN2 U574 ( .A(\add_1242/carry[6] ), .B(Term1[17]), .Z(\add_1242/carry[7] )
         );
  EO U575 ( .A(Term1[17]), .B(\add_1242/carry[6] ), .Z(N42) );
  AN2 U576 ( .A(\add_1242/carry[5] ), .B(Term1[16]), .Z(\add_1242/carry[6] )
         );
  EO U577 ( .A(Term1[16]), .B(\add_1242/carry[5] ), .Z(N41) );
  AN2 U578 ( .A(\add_1242/carry[4] ), .B(Term1[15]), .Z(\add_1242/carry[5] )
         );
  EO U579 ( .A(Term1[15]), .B(\add_1242/carry[4] ), .Z(N40) );
  AN2 U580 ( .A(\add_1242/carry[3] ), .B(Term1[14]), .Z(\add_1242/carry[4] )
         );
  EO U581 ( .A(Term1[14]), .B(\add_1242/carry[3] ), .Z(N39) );
  AN2 U582 ( .A(\add_1242/carry[2] ), .B(Term1[13]), .Z(\add_1242/carry[3] )
         );
  EO U583 ( .A(Term1[13]), .B(\add_1242/carry[2] ), .Z(N38) );
  AN2 U584 ( .A(\add_1242/carry[1] ), .B(Term1[12]), .Z(\add_1242/carry[2] )
         );
  EO U585 ( .A(Term1[12]), .B(\add_1242/carry[1] ), .Z(N37) );
  AN2 U586 ( .A(\Term2[18] ), .B(Term1[11]), .Z(\add_1242/carry[1] ) );
  EO U587 ( .A(Term1[11]), .B(\Term2[18] ), .Z(N36) );
endmodule


module AWGN_DW01_add_1 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;

  IVP U2 ( .A(n67), .Z(n14) );
  IVP U3 ( .A(n59), .Z(n12) );
  IVP U4 ( .A(n51), .Z(n10) );
  IVP U5 ( .A(n43), .Z(n8) );
  IVP U6 ( .A(n35), .Z(n6) );
  IVP U7 ( .A(n27), .Z(n4) );
  IVP U8 ( .A(n18), .Z(n1) );
  IVP U9 ( .A(n23), .Z(n3) );
  IVP U10 ( .A(n31), .Z(n5) );
  IVP U11 ( .A(n39), .Z(n7) );
  IVP U12 ( .A(n47), .Z(n9) );
  IVP U13 ( .A(n55), .Z(n11) );
  IVP U14 ( .A(n63), .Z(n13) );
  IVP U15 ( .A(n69), .Z(n15) );
  IVP U16 ( .A(n19), .Z(n2) );
  ND2 U17 ( .A(A[14]), .B(B[14]), .Z(n70) );
  EO U18 ( .A(n16), .B(B[29]), .Z(SUM[29]) );
  AO7 U19 ( .A(n17), .B(n2), .C(n18), .Z(n16) );
  EO U20 ( .A(n19), .B(n20), .Z(SUM[28]) );
  NR2 U21 ( .A(n1), .B(n17), .Z(n20) );
  NR2 U22 ( .A(B[28]), .B(A[28]), .Z(n17) );
  ND2 U23 ( .A(B[28]), .B(A[28]), .Z(n18) );
  AO7 U24 ( .A(n21), .B(n22), .C(n23), .Z(n19) );
  EN U25 ( .A(n22), .B(n24), .Z(SUM[27]) );
  NR2 U26 ( .A(n3), .B(n21), .Z(n24) );
  NR2 U27 ( .A(B[27]), .B(A[27]), .Z(n21) );
  ND2 U28 ( .A(B[27]), .B(A[27]), .Z(n23) );
  AO6 U29 ( .A(n4), .B(n25), .C(n26), .Z(n22) );
  EO U30 ( .A(n25), .B(n28), .Z(SUM[26]) );
  NR2 U31 ( .A(n26), .B(n27), .Z(n28) );
  NR2 U32 ( .A(B[26]), .B(A[26]), .Z(n27) );
  AN2 U33 ( .A(B[26]), .B(A[26]), .Z(n26) );
  AO7 U34 ( .A(n29), .B(n30), .C(n31), .Z(n25) );
  EN U35 ( .A(n30), .B(n32), .Z(SUM[25]) );
  NR2 U36 ( .A(n5), .B(n29), .Z(n32) );
  NR2 U37 ( .A(B[25]), .B(A[25]), .Z(n29) );
  ND2 U38 ( .A(B[25]), .B(A[25]), .Z(n31) );
  AO6 U39 ( .A(n6), .B(n33), .C(n34), .Z(n30) );
  EO U40 ( .A(n33), .B(n36), .Z(SUM[24]) );
  NR2 U41 ( .A(n34), .B(n35), .Z(n36) );
  NR2 U42 ( .A(B[24]), .B(A[24]), .Z(n35) );
  AN2 U43 ( .A(B[24]), .B(A[24]), .Z(n34) );
  AO7 U44 ( .A(n37), .B(n38), .C(n39), .Z(n33) );
  EN U45 ( .A(n38), .B(n40), .Z(SUM[23]) );
  NR2 U46 ( .A(n7), .B(n37), .Z(n40) );
  NR2 U47 ( .A(B[23]), .B(A[23]), .Z(n37) );
  ND2 U48 ( .A(B[23]), .B(A[23]), .Z(n39) );
  AO6 U49 ( .A(n8), .B(n41), .C(n42), .Z(n38) );
  EO U50 ( .A(n41), .B(n44), .Z(SUM[22]) );
  NR2 U51 ( .A(n42), .B(n43), .Z(n44) );
  NR2 U52 ( .A(B[22]), .B(A[22]), .Z(n43) );
  AN2 U53 ( .A(B[22]), .B(A[22]), .Z(n42) );
  AO7 U54 ( .A(n45), .B(n46), .C(n47), .Z(n41) );
  EN U55 ( .A(n46), .B(n48), .Z(SUM[21]) );
  NR2 U56 ( .A(n9), .B(n45), .Z(n48) );
  NR2 U57 ( .A(B[21]), .B(A[21]), .Z(n45) );
  ND2 U58 ( .A(B[21]), .B(A[21]), .Z(n47) );
  AO6 U59 ( .A(n10), .B(n49), .C(n50), .Z(n46) );
  EO U60 ( .A(n49), .B(n52), .Z(SUM[20]) );
  NR2 U61 ( .A(n50), .B(n51), .Z(n52) );
  NR2 U62 ( .A(B[20]), .B(A[20]), .Z(n51) );
  AN2 U63 ( .A(B[20]), .B(A[20]), .Z(n50) );
  AO7 U64 ( .A(n53), .B(n54), .C(n55), .Z(n49) );
  EN U65 ( .A(n54), .B(n56), .Z(SUM[19]) );
  NR2 U66 ( .A(n11), .B(n53), .Z(n56) );
  NR2 U67 ( .A(B[19]), .B(A[19]), .Z(n53) );
  ND2 U68 ( .A(B[19]), .B(A[19]), .Z(n55) );
  AO6 U69 ( .A(n12), .B(n57), .C(n58), .Z(n54) );
  EO U70 ( .A(n57), .B(n60), .Z(SUM[18]) );
  NR2 U71 ( .A(n58), .B(n59), .Z(n60) );
  NR2 U72 ( .A(B[18]), .B(A[18]), .Z(n59) );
  AN2 U73 ( .A(B[18]), .B(A[18]), .Z(n58) );
  AO7 U74 ( .A(n61), .B(n62), .C(n63), .Z(n57) );
  EN U75 ( .A(n62), .B(n64), .Z(SUM[17]) );
  NR2 U76 ( .A(n13), .B(n61), .Z(n64) );
  NR2 U77 ( .A(B[17]), .B(A[17]), .Z(n61) );
  ND2 U78 ( .A(B[17]), .B(A[17]), .Z(n63) );
  AO6 U79 ( .A(n14), .B(n65), .C(n66), .Z(n62) );
  EO U80 ( .A(n65), .B(n68), .Z(SUM[16]) );
  NR2 U81 ( .A(n66), .B(n67), .Z(n68) );
  NR2 U82 ( .A(B[16]), .B(A[16]), .Z(n67) );
  AN2 U83 ( .A(B[16]), .B(A[16]), .Z(n66) );
  AO7 U84 ( .A(n69), .B(n70), .C(n71), .Z(n65) );
  EO U85 ( .A(n72), .B(n70), .Z(SUM[15]) );
  ND2 U86 ( .A(n15), .B(n71), .Z(n72) );
  ND2 U87 ( .A(B[15]), .B(A[15]), .Z(n71) );
  NR2 U88 ( .A(B[15]), .B(A[15]), .Z(n69) );
endmodule


module AWGN_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [14:0] A;
  input [16:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[14][16] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][16] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][16] ,
         \ab[12][15] , \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] ,
         \ab[12][10] , \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] ,
         \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] ,
         \ab[12][0] , \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] ,
         \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] ,
         \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] ,
         \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][16] ,
         \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] ,
         \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] ,
         \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] ,
         \ab[7][0] , \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] ,
         \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] ,
         \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] ,
         \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][16] ,
         \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] ,
         \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] ,
         \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] ,
         \ab[2][0] , \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][13] , \CARRYB[14][12] , \CARRYB[14][11] ,
         \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][15] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[14][0] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] ,
         \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] ,
         \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] ,
         \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] ,
         \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] ,
         \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] ,
         \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][15] , \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] ,
         \SUMB[1][11] , \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] ,
         \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , \A1[28] , \A1[27] , \A1[26] , \A1[25] ,
         \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] ,
         \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[29] , \A2[28] , \A2[27] , \A2[26] ,
         \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] ,
         \A2[18] , \A2[17] , \A2[16] , \A2[15] , \A2[14] , n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  AWGN_DW01_add_1 FS_1 ( .A({1'b0, \A1[28] , \A1[27] , \A1[26] , \A1[25] , 
        \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , 
        \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \SUMB[14][0] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[29] , \A2[28] , 
        \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , 
        \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , \A2[14] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[31:17], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14}) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S5_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\ab[13][16] ), .CO(
        \CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S3_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\ab[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S3_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\ab[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S3_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\ab[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S3_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\ab[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S3_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\ab[8][16] ), .CO(
        \CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S3_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\ab[7][16] ), .CO(
        \CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S3_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\ab[6][16] ), .CO(
        \CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S3_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\ab[5][16] ), .CO(
        \CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S3_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\ab[4][16] ), .CO(
        \CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S3_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\ab[3][16] ), .CO(
        \CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S3_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\ab[2][16] ), .CO(
        \CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S3_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\ab[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S4_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S4_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S4_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S4_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), .CO(
        \CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S4_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), .CO(
        \CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S4_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), .CO(
        \CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S4_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), .CO(
        \CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S4_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(
        \CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S4_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(
        \CARRYB[14][0] ), .S(\SUMB[14][0] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S4_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(
        \CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S4_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(
        \CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S4_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), .CO(
        \CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), .CO(
        \CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  EO U2 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A1[15] ) );
  EO U3 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A1[14] ) );
  EO U4 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A1[16] ) );
  EO U5 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A1[18] ) );
  EO U6 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A1[17] ) );
  EO U7 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A1[20] ) );
  EO U8 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A1[19] ) );
  EO U9 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A1[21] ) );
  EO U10 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A1[22] ) );
  EO U11 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A1[23] ) );
  EO U12 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A1[24] ) );
  EO U13 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A1[25] ) );
  EO U14 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A1[26] ) );
  EO U15 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A1[27] ) );
  EO U16 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A1[28] ) );
  EO U17 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A1[13] ) );
  EO U18 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U19 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U20 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U21 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U22 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U23 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U24 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U25 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U26 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U27 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U28 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U29 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U30 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U31 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  IVP U32 ( .A(A[1]), .Z(n33) );
  IVP U33 ( .A(B[2]), .Z(n17) );
  IVP U34 ( .A(B[3]), .Z(n16) );
  IVP U35 ( .A(B[4]), .Z(n15) );
  IVP U36 ( .A(B[1]), .Z(n18) );
  IVP U37 ( .A(A[2]), .Z(n32) );
  IVP U38 ( .A(A[0]), .Z(n34) );
  IVP U39 ( .A(B[5]), .Z(n14) );
  IVP U40 ( .A(B[6]), .Z(n13) );
  EO U41 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  IVP U42 ( .A(B[7]), .Z(n12) );
  IVP U43 ( .A(B[0]), .Z(n19) );
  IVP U44 ( .A(B[8]), .Z(n11) );
  IVP U45 ( .A(A[3]), .Z(n31) );
  IVP U46 ( .A(B[9]), .Z(n10) );
  IVP U47 ( .A(B[10]), .Z(n9) );
  IVP U48 ( .A(A[4]), .Z(n30) );
  IVP U49 ( .A(B[11]), .Z(n8) );
  IVP U50 ( .A(B[12]), .Z(n7) );
  IVP U51 ( .A(A[5]), .Z(n29) );
  IVP U52 ( .A(B[13]), .Z(n6) );
  IVP U53 ( .A(B[14]), .Z(n5) );
  IVP U54 ( .A(B[15]), .Z(n4) );
  IVP U55 ( .A(B[16]), .Z(n3) );
  IVP U56 ( .A(A[6]), .Z(n28) );
  IVP U57 ( .A(A[7]), .Z(n27) );
  IVP U58 ( .A(A[8]), .Z(n26) );
  IVP U59 ( .A(A[9]), .Z(n25) );
  IVP U60 ( .A(A[10]), .Z(n24) );
  IVP U61 ( .A(A[11]), .Z(n23) );
  IVP U62 ( .A(A[12]), .Z(n22) );
  IVP U63 ( .A(A[13]), .Z(n21) );
  IVP U64 ( .A(A[14]), .Z(n20) );
  AN2P U65 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A2[14] ) );
  AN2P U66 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A2[16] ) );
  AN2P U67 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A2[17] ) );
  AN2P U68 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A2[18] ) );
  AN2P U69 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A2[19] ) );
  AN2P U70 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A2[20] ) );
  AN2P U71 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A2[21] ) );
  AN2P U72 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A2[22] ) );
  AN2P U73 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A2[23] ) );
  AN2P U74 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A2[24] ) );
  AN2P U75 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A2[25] ) );
  AN2P U76 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A2[26] ) );
  AN2P U77 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A2[27] ) );
  AN2P U78 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A2[28] ) );
  AN2P U79 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A2[29] ) );
  AN2P U80 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U81 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U82 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U83 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U84 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U85 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U86 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U87 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U88 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U89 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U90 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U91 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U92 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U93 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U94 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U95 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A2[15] ) );
  NR2 U97 ( .A(n25), .B(n10), .Z(\ab[9][9] ) );
  NR2 U98 ( .A(n25), .B(n11), .Z(\ab[9][8] ) );
  NR2 U99 ( .A(n25), .B(n12), .Z(\ab[9][7] ) );
  NR2 U100 ( .A(n25), .B(n13), .Z(\ab[9][6] ) );
  NR2 U101 ( .A(n25), .B(n14), .Z(\ab[9][5] ) );
  NR2 U102 ( .A(n25), .B(n15), .Z(\ab[9][4] ) );
  NR2 U103 ( .A(n25), .B(n16), .Z(\ab[9][3] ) );
  NR2 U104 ( .A(n25), .B(n17), .Z(\ab[9][2] ) );
  NR2 U105 ( .A(n25), .B(n18), .Z(\ab[9][1] ) );
  NR2 U106 ( .A(n25), .B(n3), .Z(\ab[9][16] ) );
  NR2 U107 ( .A(n25), .B(n4), .Z(\ab[9][15] ) );
  NR2 U108 ( .A(n25), .B(n5), .Z(\ab[9][14] ) );
  NR2 U109 ( .A(n25), .B(n6), .Z(\ab[9][13] ) );
  NR2 U110 ( .A(n25), .B(n7), .Z(\ab[9][12] ) );
  NR2 U111 ( .A(n25), .B(n8), .Z(\ab[9][11] ) );
  NR2 U112 ( .A(n25), .B(n9), .Z(\ab[9][10] ) );
  NR2 U113 ( .A(n25), .B(n19), .Z(\ab[9][0] ) );
  NR2 U114 ( .A(n10), .B(n26), .Z(\ab[8][9] ) );
  NR2 U115 ( .A(n11), .B(n26), .Z(\ab[8][8] ) );
  NR2 U116 ( .A(n12), .B(n26), .Z(\ab[8][7] ) );
  NR2 U117 ( .A(n13), .B(n26), .Z(\ab[8][6] ) );
  NR2 U118 ( .A(n14), .B(n26), .Z(\ab[8][5] ) );
  NR2 U119 ( .A(n15), .B(n26), .Z(\ab[8][4] ) );
  NR2 U120 ( .A(n16), .B(n26), .Z(\ab[8][3] ) );
  NR2 U121 ( .A(n17), .B(n26), .Z(\ab[8][2] ) );
  NR2 U122 ( .A(n18), .B(n26), .Z(\ab[8][1] ) );
  NR2 U123 ( .A(n3), .B(n26), .Z(\ab[8][16] ) );
  NR2 U124 ( .A(n4), .B(n26), .Z(\ab[8][15] ) );
  NR2 U125 ( .A(n5), .B(n26), .Z(\ab[8][14] ) );
  NR2 U126 ( .A(n6), .B(n26), .Z(\ab[8][13] ) );
  NR2 U127 ( .A(n7), .B(n26), .Z(\ab[8][12] ) );
  NR2 U128 ( .A(n8), .B(n26), .Z(\ab[8][11] ) );
  NR2 U129 ( .A(n9), .B(n26), .Z(\ab[8][10] ) );
  NR2 U130 ( .A(n19), .B(n26), .Z(\ab[8][0] ) );
  NR2 U131 ( .A(n10), .B(n27), .Z(\ab[7][9] ) );
  NR2 U132 ( .A(n11), .B(n27), .Z(\ab[7][8] ) );
  NR2 U133 ( .A(n12), .B(n27), .Z(\ab[7][7] ) );
  NR2 U134 ( .A(n13), .B(n27), .Z(\ab[7][6] ) );
  NR2 U135 ( .A(n14), .B(n27), .Z(\ab[7][5] ) );
  NR2 U136 ( .A(n15), .B(n27), .Z(\ab[7][4] ) );
  NR2 U137 ( .A(n16), .B(n27), .Z(\ab[7][3] ) );
  NR2 U138 ( .A(n17), .B(n27), .Z(\ab[7][2] ) );
  NR2 U139 ( .A(n18), .B(n27), .Z(\ab[7][1] ) );
  NR2 U140 ( .A(n3), .B(n27), .Z(\ab[7][16] ) );
  NR2 U141 ( .A(n4), .B(n27), .Z(\ab[7][15] ) );
  NR2 U142 ( .A(n5), .B(n27), .Z(\ab[7][14] ) );
  NR2 U143 ( .A(n6), .B(n27), .Z(\ab[7][13] ) );
  NR2 U144 ( .A(n7), .B(n27), .Z(\ab[7][12] ) );
  NR2 U145 ( .A(n8), .B(n27), .Z(\ab[7][11] ) );
  NR2 U146 ( .A(n9), .B(n27), .Z(\ab[7][10] ) );
  NR2 U147 ( .A(n19), .B(n27), .Z(\ab[7][0] ) );
  NR2 U148 ( .A(n10), .B(n28), .Z(\ab[6][9] ) );
  NR2 U149 ( .A(n11), .B(n28), .Z(\ab[6][8] ) );
  NR2 U150 ( .A(n12), .B(n28), .Z(\ab[6][7] ) );
  NR2 U151 ( .A(n13), .B(n28), .Z(\ab[6][6] ) );
  NR2 U152 ( .A(n14), .B(n28), .Z(\ab[6][5] ) );
  NR2 U153 ( .A(n15), .B(n28), .Z(\ab[6][4] ) );
  NR2 U154 ( .A(n16), .B(n28), .Z(\ab[6][3] ) );
  NR2 U155 ( .A(n17), .B(n28), .Z(\ab[6][2] ) );
  NR2 U156 ( .A(n18), .B(n28), .Z(\ab[6][1] ) );
  NR2 U157 ( .A(n3), .B(n28), .Z(\ab[6][16] ) );
  NR2 U158 ( .A(n4), .B(n28), .Z(\ab[6][15] ) );
  NR2 U159 ( .A(n5), .B(n28), .Z(\ab[6][14] ) );
  NR2 U160 ( .A(n6), .B(n28), .Z(\ab[6][13] ) );
  NR2 U161 ( .A(n7), .B(n28), .Z(\ab[6][12] ) );
  NR2 U162 ( .A(n8), .B(n28), .Z(\ab[6][11] ) );
  NR2 U163 ( .A(n9), .B(n28), .Z(\ab[6][10] ) );
  NR2 U164 ( .A(n19), .B(n28), .Z(\ab[6][0] ) );
  NR2 U165 ( .A(n10), .B(n29), .Z(\ab[5][9] ) );
  NR2 U166 ( .A(n11), .B(n29), .Z(\ab[5][8] ) );
  NR2 U167 ( .A(n12), .B(n29), .Z(\ab[5][7] ) );
  NR2 U168 ( .A(n13), .B(n29), .Z(\ab[5][6] ) );
  NR2 U169 ( .A(n14), .B(n29), .Z(\ab[5][5] ) );
  NR2 U170 ( .A(n15), .B(n29), .Z(\ab[5][4] ) );
  NR2 U171 ( .A(n16), .B(n29), .Z(\ab[5][3] ) );
  NR2 U172 ( .A(n17), .B(n29), .Z(\ab[5][2] ) );
  NR2 U173 ( .A(n18), .B(n29), .Z(\ab[5][1] ) );
  NR2 U174 ( .A(n3), .B(n29), .Z(\ab[5][16] ) );
  NR2 U175 ( .A(n4), .B(n29), .Z(\ab[5][15] ) );
  NR2 U176 ( .A(n5), .B(n29), .Z(\ab[5][14] ) );
  NR2 U177 ( .A(n6), .B(n29), .Z(\ab[5][13] ) );
  NR2 U178 ( .A(n7), .B(n29), .Z(\ab[5][12] ) );
  NR2 U179 ( .A(n8), .B(n29), .Z(\ab[5][11] ) );
  NR2 U180 ( .A(n9), .B(n29), .Z(\ab[5][10] ) );
  NR2 U181 ( .A(n19), .B(n29), .Z(\ab[5][0] ) );
  NR2 U182 ( .A(n10), .B(n30), .Z(\ab[4][9] ) );
  NR2 U183 ( .A(n11), .B(n30), .Z(\ab[4][8] ) );
  NR2 U184 ( .A(n12), .B(n30), .Z(\ab[4][7] ) );
  NR2 U185 ( .A(n13), .B(n30), .Z(\ab[4][6] ) );
  NR2 U186 ( .A(n14), .B(n30), .Z(\ab[4][5] ) );
  NR2 U187 ( .A(n15), .B(n30), .Z(\ab[4][4] ) );
  NR2 U188 ( .A(n16), .B(n30), .Z(\ab[4][3] ) );
  NR2 U189 ( .A(n17), .B(n30), .Z(\ab[4][2] ) );
  NR2 U190 ( .A(n18), .B(n30), .Z(\ab[4][1] ) );
  NR2 U191 ( .A(n3), .B(n30), .Z(\ab[4][16] ) );
  NR2 U192 ( .A(n4), .B(n30), .Z(\ab[4][15] ) );
  NR2 U193 ( .A(n5), .B(n30), .Z(\ab[4][14] ) );
  NR2 U194 ( .A(n6), .B(n30), .Z(\ab[4][13] ) );
  NR2 U195 ( .A(n7), .B(n30), .Z(\ab[4][12] ) );
  NR2 U196 ( .A(n8), .B(n30), .Z(\ab[4][11] ) );
  NR2 U197 ( .A(n9), .B(n30), .Z(\ab[4][10] ) );
  NR2 U198 ( .A(n19), .B(n30), .Z(\ab[4][0] ) );
  NR2 U199 ( .A(n10), .B(n31), .Z(\ab[3][9] ) );
  NR2 U200 ( .A(n11), .B(n31), .Z(\ab[3][8] ) );
  NR2 U201 ( .A(n12), .B(n31), .Z(\ab[3][7] ) );
  NR2 U202 ( .A(n13), .B(n31), .Z(\ab[3][6] ) );
  NR2 U203 ( .A(n14), .B(n31), .Z(\ab[3][5] ) );
  NR2 U204 ( .A(n15), .B(n31), .Z(\ab[3][4] ) );
  NR2 U205 ( .A(n16), .B(n31), .Z(\ab[3][3] ) );
  NR2 U206 ( .A(n17), .B(n31), .Z(\ab[3][2] ) );
  NR2 U207 ( .A(n18), .B(n31), .Z(\ab[3][1] ) );
  NR2 U208 ( .A(n3), .B(n31), .Z(\ab[3][16] ) );
  NR2 U209 ( .A(n4), .B(n31), .Z(\ab[3][15] ) );
  NR2 U210 ( .A(n5), .B(n31), .Z(\ab[3][14] ) );
  NR2 U211 ( .A(n6), .B(n31), .Z(\ab[3][13] ) );
  NR2 U212 ( .A(n7), .B(n31), .Z(\ab[3][12] ) );
  NR2 U213 ( .A(n8), .B(n31), .Z(\ab[3][11] ) );
  NR2 U214 ( .A(n9), .B(n31), .Z(\ab[3][10] ) );
  NR2 U215 ( .A(n19), .B(n31), .Z(\ab[3][0] ) );
  NR2 U216 ( .A(n10), .B(n32), .Z(\ab[2][9] ) );
  NR2 U217 ( .A(n11), .B(n32), .Z(\ab[2][8] ) );
  NR2 U218 ( .A(n12), .B(n32), .Z(\ab[2][7] ) );
  NR2 U219 ( .A(n13), .B(n32), .Z(\ab[2][6] ) );
  NR2 U220 ( .A(n14), .B(n32), .Z(\ab[2][5] ) );
  NR2 U221 ( .A(n15), .B(n32), .Z(\ab[2][4] ) );
  NR2 U222 ( .A(n16), .B(n32), .Z(\ab[2][3] ) );
  NR2 U223 ( .A(n17), .B(n32), .Z(\ab[2][2] ) );
  NR2 U224 ( .A(n18), .B(n32), .Z(\ab[2][1] ) );
  NR2 U225 ( .A(n3), .B(n32), .Z(\ab[2][16] ) );
  NR2 U226 ( .A(n4), .B(n32), .Z(\ab[2][15] ) );
  NR2 U227 ( .A(n5), .B(n32), .Z(\ab[2][14] ) );
  NR2 U228 ( .A(n6), .B(n32), .Z(\ab[2][13] ) );
  NR2 U229 ( .A(n7), .B(n32), .Z(\ab[2][12] ) );
  NR2 U230 ( .A(n8), .B(n32), .Z(\ab[2][11] ) );
  NR2 U231 ( .A(n9), .B(n32), .Z(\ab[2][10] ) );
  NR2 U232 ( .A(n19), .B(n32), .Z(\ab[2][0] ) );
  NR2 U233 ( .A(n10), .B(n33), .Z(\ab[1][9] ) );
  NR2 U234 ( .A(n11), .B(n33), .Z(\ab[1][8] ) );
  NR2 U235 ( .A(n12), .B(n33), .Z(\ab[1][7] ) );
  NR2 U236 ( .A(n13), .B(n33), .Z(\ab[1][6] ) );
  NR2 U237 ( .A(n14), .B(n33), .Z(\ab[1][5] ) );
  NR2 U238 ( .A(n15), .B(n33), .Z(\ab[1][4] ) );
  NR2 U239 ( .A(n16), .B(n33), .Z(\ab[1][3] ) );
  NR2 U240 ( .A(n17), .B(n33), .Z(\ab[1][2] ) );
  NR2 U241 ( .A(n3), .B(n33), .Z(\ab[1][16] ) );
  NR2 U242 ( .A(n4), .B(n33), .Z(\ab[1][15] ) );
  NR2 U243 ( .A(n5), .B(n33), .Z(\ab[1][14] ) );
  NR2 U244 ( .A(n6), .B(n33), .Z(\ab[1][13] ) );
  NR2 U245 ( .A(n7), .B(n33), .Z(\ab[1][12] ) );
  NR2 U246 ( .A(n8), .B(n33), .Z(\ab[1][11] ) );
  NR2 U247 ( .A(n9), .B(n33), .Z(\ab[1][10] ) );
  NR2 U248 ( .A(n10), .B(n20), .Z(\ab[14][9] ) );
  NR2 U249 ( .A(n11), .B(n20), .Z(\ab[14][8] ) );
  NR2 U250 ( .A(n12), .B(n20), .Z(\ab[14][7] ) );
  NR2 U251 ( .A(n13), .B(n20), .Z(\ab[14][6] ) );
  NR2 U252 ( .A(n14), .B(n20), .Z(\ab[14][5] ) );
  NR2 U253 ( .A(n15), .B(n20), .Z(\ab[14][4] ) );
  NR2 U254 ( .A(n16), .B(n20), .Z(\ab[14][3] ) );
  NR2 U255 ( .A(n17), .B(n20), .Z(\ab[14][2] ) );
  NR2 U256 ( .A(n18), .B(n20), .Z(\ab[14][1] ) );
  NR2 U257 ( .A(n3), .B(n20), .Z(\ab[14][16] ) );
  NR2 U258 ( .A(n4), .B(n20), .Z(\ab[14][15] ) );
  NR2 U259 ( .A(n5), .B(n20), .Z(\ab[14][14] ) );
  NR2 U260 ( .A(n6), .B(n20), .Z(\ab[14][13] ) );
  NR2 U261 ( .A(n7), .B(n20), .Z(\ab[14][12] ) );
  NR2 U262 ( .A(n8), .B(n20), .Z(\ab[14][11] ) );
  NR2 U263 ( .A(n9), .B(n20), .Z(\ab[14][10] ) );
  NR2 U264 ( .A(n19), .B(n20), .Z(\ab[14][0] ) );
  NR2 U265 ( .A(n10), .B(n21), .Z(\ab[13][9] ) );
  NR2 U266 ( .A(n11), .B(n21), .Z(\ab[13][8] ) );
  NR2 U267 ( .A(n12), .B(n21), .Z(\ab[13][7] ) );
  NR2 U268 ( .A(n13), .B(n21), .Z(\ab[13][6] ) );
  NR2 U269 ( .A(n14), .B(n21), .Z(\ab[13][5] ) );
  NR2 U270 ( .A(n15), .B(n21), .Z(\ab[13][4] ) );
  NR2 U271 ( .A(n16), .B(n21), .Z(\ab[13][3] ) );
  NR2 U272 ( .A(n17), .B(n21), .Z(\ab[13][2] ) );
  NR2 U273 ( .A(n18), .B(n21), .Z(\ab[13][1] ) );
  NR2 U274 ( .A(n3), .B(n21), .Z(\ab[13][16] ) );
  NR2 U275 ( .A(n4), .B(n21), .Z(\ab[13][15] ) );
  NR2 U276 ( .A(n5), .B(n21), .Z(\ab[13][14] ) );
  NR2 U277 ( .A(n6), .B(n21), .Z(\ab[13][13] ) );
  NR2 U278 ( .A(n7), .B(n21), .Z(\ab[13][12] ) );
  NR2 U279 ( .A(n8), .B(n21), .Z(\ab[13][11] ) );
  NR2 U280 ( .A(n9), .B(n21), .Z(\ab[13][10] ) );
  NR2 U281 ( .A(n19), .B(n21), .Z(\ab[13][0] ) );
  NR2 U282 ( .A(n10), .B(n22), .Z(\ab[12][9] ) );
  NR2 U283 ( .A(n11), .B(n22), .Z(\ab[12][8] ) );
  NR2 U284 ( .A(n12), .B(n22), .Z(\ab[12][7] ) );
  NR2 U285 ( .A(n13), .B(n22), .Z(\ab[12][6] ) );
  NR2 U286 ( .A(n14), .B(n22), .Z(\ab[12][5] ) );
  NR2 U287 ( .A(n15), .B(n22), .Z(\ab[12][4] ) );
  NR2 U288 ( .A(n16), .B(n22), .Z(\ab[12][3] ) );
  NR2 U289 ( .A(n17), .B(n22), .Z(\ab[12][2] ) );
  NR2 U290 ( .A(n18), .B(n22), .Z(\ab[12][1] ) );
  NR2 U291 ( .A(n3), .B(n22), .Z(\ab[12][16] ) );
  NR2 U292 ( .A(n4), .B(n22), .Z(\ab[12][15] ) );
  NR2 U293 ( .A(n5), .B(n22), .Z(\ab[12][14] ) );
  NR2 U294 ( .A(n6), .B(n22), .Z(\ab[12][13] ) );
  NR2 U295 ( .A(n7), .B(n22), .Z(\ab[12][12] ) );
  NR2 U296 ( .A(n8), .B(n22), .Z(\ab[12][11] ) );
  NR2 U297 ( .A(n9), .B(n22), .Z(\ab[12][10] ) );
  NR2 U298 ( .A(n19), .B(n22), .Z(\ab[12][0] ) );
  NR2 U299 ( .A(n10), .B(n23), .Z(\ab[11][9] ) );
  NR2 U300 ( .A(n11), .B(n23), .Z(\ab[11][8] ) );
  NR2 U301 ( .A(n12), .B(n23), .Z(\ab[11][7] ) );
  NR2 U302 ( .A(n13), .B(n23), .Z(\ab[11][6] ) );
  NR2 U303 ( .A(n14), .B(n23), .Z(\ab[11][5] ) );
  NR2 U304 ( .A(n15), .B(n23), .Z(\ab[11][4] ) );
  NR2 U305 ( .A(n16), .B(n23), .Z(\ab[11][3] ) );
  NR2 U306 ( .A(n17), .B(n23), .Z(\ab[11][2] ) );
  NR2 U307 ( .A(n18), .B(n23), .Z(\ab[11][1] ) );
  NR2 U308 ( .A(n3), .B(n23), .Z(\ab[11][16] ) );
  NR2 U309 ( .A(n4), .B(n23), .Z(\ab[11][15] ) );
  NR2 U310 ( .A(n5), .B(n23), .Z(\ab[11][14] ) );
  NR2 U311 ( .A(n6), .B(n23), .Z(\ab[11][13] ) );
  NR2 U312 ( .A(n7), .B(n23), .Z(\ab[11][12] ) );
  NR2 U313 ( .A(n8), .B(n23), .Z(\ab[11][11] ) );
  NR2 U314 ( .A(n9), .B(n23), .Z(\ab[11][10] ) );
  NR2 U315 ( .A(n19), .B(n23), .Z(\ab[11][0] ) );
  NR2 U316 ( .A(n10), .B(n24), .Z(\ab[10][9] ) );
  NR2 U317 ( .A(n11), .B(n24), .Z(\ab[10][8] ) );
  NR2 U318 ( .A(n12), .B(n24), .Z(\ab[10][7] ) );
  NR2 U319 ( .A(n13), .B(n24), .Z(\ab[10][6] ) );
  NR2 U320 ( .A(n14), .B(n24), .Z(\ab[10][5] ) );
  NR2 U321 ( .A(n15), .B(n24), .Z(\ab[10][4] ) );
  NR2 U322 ( .A(n16), .B(n24), .Z(\ab[10][3] ) );
  NR2 U323 ( .A(n17), .B(n24), .Z(\ab[10][2] ) );
  NR2 U324 ( .A(n18), .B(n24), .Z(\ab[10][1] ) );
  NR2 U325 ( .A(n3), .B(n24), .Z(\ab[10][16] ) );
  NR2 U326 ( .A(n4), .B(n24), .Z(\ab[10][15] ) );
  NR2 U327 ( .A(n5), .B(n24), .Z(\ab[10][14] ) );
  NR2 U328 ( .A(n6), .B(n24), .Z(\ab[10][13] ) );
  NR2 U329 ( .A(n7), .B(n24), .Z(\ab[10][12] ) );
  NR2 U330 ( .A(n8), .B(n24), .Z(\ab[10][11] ) );
  NR2 U331 ( .A(n9), .B(n24), .Z(\ab[10][10] ) );
  NR2 U332 ( .A(n19), .B(n24), .Z(\ab[10][0] ) );
  NR2 U333 ( .A(n10), .B(n34), .Z(\ab[0][9] ) );
  NR2 U334 ( .A(n11), .B(n34), .Z(\ab[0][8] ) );
  NR2 U335 ( .A(n12), .B(n34), .Z(\ab[0][7] ) );
  NR2 U336 ( .A(n13), .B(n34), .Z(\ab[0][6] ) );
  NR2 U337 ( .A(n14), .B(n34), .Z(\ab[0][5] ) );
  NR2 U338 ( .A(n15), .B(n34), .Z(\ab[0][4] ) );
  NR2 U339 ( .A(n16), .B(n34), .Z(\ab[0][3] ) );
  NR2 U340 ( .A(n17), .B(n34), .Z(\ab[0][2] ) );
  NR2 U341 ( .A(n3), .B(n34), .Z(\ab[0][16] ) );
  NR2 U342 ( .A(n4), .B(n34), .Z(\ab[0][15] ) );
  NR2 U343 ( .A(n5), .B(n34), .Z(\ab[0][14] ) );
  NR2 U344 ( .A(n6), .B(n34), .Z(\ab[0][13] ) );
  NR2 U345 ( .A(n7), .B(n34), .Z(\ab[0][12] ) );
  NR2 U346 ( .A(n8), .B(n34), .Z(\ab[0][11] ) );
  NR2 U347 ( .A(n9), .B(n34), .Z(\ab[0][10] ) );
  AN3 U348 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U349 ( .A(n33), .B(n18), .Z(\ab[1][1] ) );
endmodule


module AWGN_DW01_add_0 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;

  IVP U2 ( .A(n67), .Z(n14) );
  IVP U3 ( .A(n59), .Z(n12) );
  IVP U4 ( .A(n51), .Z(n10) );
  IVP U5 ( .A(n43), .Z(n8) );
  IVP U6 ( .A(n35), .Z(n6) );
  IVP U7 ( .A(n27), .Z(n4) );
  IVP U8 ( .A(n18), .Z(n1) );
  IVP U9 ( .A(n23), .Z(n3) );
  IVP U10 ( .A(n31), .Z(n5) );
  IVP U11 ( .A(n39), .Z(n7) );
  IVP U12 ( .A(n47), .Z(n9) );
  IVP U13 ( .A(n55), .Z(n11) );
  IVP U14 ( .A(n63), .Z(n13) );
  IVP U15 ( .A(n69), .Z(n15) );
  IVP U16 ( .A(n19), .Z(n2) );
  ND2 U17 ( .A(A[14]), .B(B[14]), .Z(n70) );
  EO U18 ( .A(n16), .B(B[29]), .Z(SUM[29]) );
  AO7 U19 ( .A(n17), .B(n2), .C(n18), .Z(n16) );
  EO U20 ( .A(n19), .B(n20), .Z(SUM[28]) );
  NR2 U21 ( .A(n1), .B(n17), .Z(n20) );
  NR2 U22 ( .A(B[28]), .B(A[28]), .Z(n17) );
  ND2 U23 ( .A(B[28]), .B(A[28]), .Z(n18) );
  AO7 U24 ( .A(n21), .B(n22), .C(n23), .Z(n19) );
  EN U25 ( .A(n22), .B(n24), .Z(SUM[27]) );
  NR2 U26 ( .A(n3), .B(n21), .Z(n24) );
  NR2 U27 ( .A(B[27]), .B(A[27]), .Z(n21) );
  ND2 U28 ( .A(B[27]), .B(A[27]), .Z(n23) );
  AO6 U29 ( .A(n4), .B(n25), .C(n26), .Z(n22) );
  EO U30 ( .A(n25), .B(n28), .Z(SUM[26]) );
  NR2 U31 ( .A(n26), .B(n27), .Z(n28) );
  NR2 U32 ( .A(B[26]), .B(A[26]), .Z(n27) );
  AN2 U33 ( .A(B[26]), .B(A[26]), .Z(n26) );
  AO7 U34 ( .A(n29), .B(n30), .C(n31), .Z(n25) );
  EN U35 ( .A(n30), .B(n32), .Z(SUM[25]) );
  NR2 U36 ( .A(n5), .B(n29), .Z(n32) );
  NR2 U37 ( .A(B[25]), .B(A[25]), .Z(n29) );
  ND2 U38 ( .A(B[25]), .B(A[25]), .Z(n31) );
  AO6 U39 ( .A(n6), .B(n33), .C(n34), .Z(n30) );
  EO U40 ( .A(n33), .B(n36), .Z(SUM[24]) );
  NR2 U41 ( .A(n34), .B(n35), .Z(n36) );
  NR2 U42 ( .A(B[24]), .B(A[24]), .Z(n35) );
  AN2 U43 ( .A(B[24]), .B(A[24]), .Z(n34) );
  AO7 U44 ( .A(n37), .B(n38), .C(n39), .Z(n33) );
  EN U45 ( .A(n38), .B(n40), .Z(SUM[23]) );
  NR2 U46 ( .A(n7), .B(n37), .Z(n40) );
  NR2 U47 ( .A(B[23]), .B(A[23]), .Z(n37) );
  ND2 U48 ( .A(B[23]), .B(A[23]), .Z(n39) );
  AO6 U49 ( .A(n8), .B(n41), .C(n42), .Z(n38) );
  EO U50 ( .A(n41), .B(n44), .Z(SUM[22]) );
  NR2 U51 ( .A(n42), .B(n43), .Z(n44) );
  NR2 U52 ( .A(B[22]), .B(A[22]), .Z(n43) );
  AN2 U53 ( .A(B[22]), .B(A[22]), .Z(n42) );
  AO7 U54 ( .A(n45), .B(n46), .C(n47), .Z(n41) );
  EN U55 ( .A(n46), .B(n48), .Z(SUM[21]) );
  NR2 U56 ( .A(n9), .B(n45), .Z(n48) );
  NR2 U57 ( .A(B[21]), .B(A[21]), .Z(n45) );
  ND2 U58 ( .A(B[21]), .B(A[21]), .Z(n47) );
  AO6 U59 ( .A(n10), .B(n49), .C(n50), .Z(n46) );
  EO U60 ( .A(n49), .B(n52), .Z(SUM[20]) );
  NR2 U61 ( .A(n50), .B(n51), .Z(n52) );
  NR2 U62 ( .A(B[20]), .B(A[20]), .Z(n51) );
  AN2 U63 ( .A(B[20]), .B(A[20]), .Z(n50) );
  AO7 U64 ( .A(n53), .B(n54), .C(n55), .Z(n49) );
  EN U65 ( .A(n54), .B(n56), .Z(SUM[19]) );
  NR2 U66 ( .A(n11), .B(n53), .Z(n56) );
  NR2 U67 ( .A(B[19]), .B(A[19]), .Z(n53) );
  ND2 U68 ( .A(B[19]), .B(A[19]), .Z(n55) );
  AO6 U69 ( .A(n12), .B(n57), .C(n58), .Z(n54) );
  EO U70 ( .A(n57), .B(n60), .Z(SUM[18]) );
  NR2 U71 ( .A(n58), .B(n59), .Z(n60) );
  NR2 U72 ( .A(B[18]), .B(A[18]), .Z(n59) );
  AN2 U73 ( .A(B[18]), .B(A[18]), .Z(n58) );
  AO7 U74 ( .A(n61), .B(n62), .C(n63), .Z(n57) );
  EN U75 ( .A(n62), .B(n64), .Z(SUM[17]) );
  NR2 U76 ( .A(n13), .B(n61), .Z(n64) );
  NR2 U77 ( .A(B[17]), .B(A[17]), .Z(n61) );
  ND2 U78 ( .A(B[17]), .B(A[17]), .Z(n63) );
  AO6 U79 ( .A(n14), .B(n65), .C(n66), .Z(n62) );
  EO U80 ( .A(n65), .B(n68), .Z(SUM[16]) );
  NR2 U81 ( .A(n66), .B(n67), .Z(n68) );
  NR2 U82 ( .A(B[16]), .B(A[16]), .Z(n67) );
  AN2 U83 ( .A(B[16]), .B(A[16]), .Z(n66) );
  AO7 U84 ( .A(n69), .B(n70), .C(n71), .Z(n65) );
  EO U85 ( .A(n72), .B(n70), .Z(SUM[15]) );
  ND2 U86 ( .A(n15), .B(n71), .Z(n72) );
  ND2 U87 ( .A(B[15]), .B(A[15]), .Z(n71) );
  NR2 U88 ( .A(B[15]), .B(A[15]), .Z(n69) );
endmodule


module AWGN_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [14:0] A;
  input [16:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[14][16] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][16] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][16] ,
         \ab[12][15] , \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] ,
         \ab[12][10] , \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] ,
         \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] ,
         \ab[12][0] , \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] ,
         \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] ,
         \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] ,
         \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][16] ,
         \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] ,
         \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] ,
         \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] ,
         \ab[7][0] , \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] ,
         \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] ,
         \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] ,
         \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][16] ,
         \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] ,
         \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] ,
         \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] ,
         \ab[2][0] , \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][13] , \CARRYB[14][12] , \CARRYB[14][11] ,
         \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][15] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[14][0] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] ,
         \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] ,
         \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] ,
         \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] ,
         \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] ,
         \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] ,
         \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][15] , \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] ,
         \SUMB[1][11] , \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] ,
         \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , \A1[28] , \A1[27] , \A1[26] , \A1[25] ,
         \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] ,
         \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[29] , \A2[28] , \A2[27] , \A2[26] ,
         \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] ,
         \A2[18] , \A2[17] , \A2[16] , \A2[15] , \A2[14] , n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  AWGN_DW01_add_0 FS_1 ( .A({1'b0, \A1[28] , \A1[27] , \A1[26] , \A1[25] , 
        \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , 
        \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \SUMB[14][0] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[29] , \A2[28] , 
        \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , 
        \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , \A2[14] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[31:17], SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14}) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S5_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\ab[13][16] ), .CO(
        \CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S3_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\ab[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S3_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\ab[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S3_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\ab[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S3_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\ab[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S3_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\ab[8][16] ), .CO(
        \CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S3_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\ab[7][16] ), .CO(
        \CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S3_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\ab[6][16] ), .CO(
        \CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S3_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\ab[5][16] ), .CO(
        \CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S3_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\ab[4][16] ), .CO(
        \CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S3_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\ab[3][16] ), .CO(
        \CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S3_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\ab[2][16] ), .CO(
        \CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S3_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\ab[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S4_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S4_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S4_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S4_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), .CO(
        \CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S4_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), .CO(
        \CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S4_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), .CO(
        \CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S4_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), .CO(
        \CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S4_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(
        \CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S4_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(
        \CARRYB[14][0] ), .S(\SUMB[14][0] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S4_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(
        \CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S4_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(
        \CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S4_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), .CO(
        \CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), .CO(
        \CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  EO U2 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A1[15] ) );
  EO U3 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A1[14] ) );
  EO U4 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A1[16] ) );
  EO U5 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A1[18] ) );
  EO U6 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A1[17] ) );
  EO U7 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A1[20] ) );
  EO U8 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A1[19] ) );
  EO U9 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A1[21] ) );
  EO U10 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A1[22] ) );
  EO U11 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A1[23] ) );
  EO U12 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A1[24] ) );
  EO U13 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A1[25] ) );
  EO U14 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A1[26] ) );
  EO U15 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A1[27] ) );
  EO U16 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A1[28] ) );
  EO U17 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A1[13] ) );
  EO U18 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U19 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U20 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U21 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U22 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U23 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U24 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U25 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U26 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U27 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U28 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U29 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U30 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U31 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  IVP U32 ( .A(A[1]), .Z(n33) );
  IVP U33 ( .A(B[2]), .Z(n17) );
  IVP U34 ( .A(B[3]), .Z(n16) );
  IVP U35 ( .A(B[4]), .Z(n15) );
  IVP U36 ( .A(B[1]), .Z(n18) );
  IVP U37 ( .A(A[2]), .Z(n32) );
  IVP U38 ( .A(A[0]), .Z(n34) );
  IVP U39 ( .A(B[5]), .Z(n14) );
  IVP U40 ( .A(B[6]), .Z(n13) );
  EO U41 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  IVP U42 ( .A(B[7]), .Z(n12) );
  IVP U43 ( .A(B[0]), .Z(n19) );
  IVP U44 ( .A(B[8]), .Z(n11) );
  IVP U45 ( .A(A[3]), .Z(n31) );
  IVP U46 ( .A(B[9]), .Z(n10) );
  IVP U47 ( .A(B[10]), .Z(n9) );
  IVP U48 ( .A(A[4]), .Z(n30) );
  IVP U49 ( .A(B[11]), .Z(n8) );
  IVP U50 ( .A(B[12]), .Z(n7) );
  IVP U51 ( .A(A[5]), .Z(n29) );
  IVP U52 ( .A(B[13]), .Z(n6) );
  IVP U53 ( .A(B[14]), .Z(n5) );
  IVP U54 ( .A(B[15]), .Z(n4) );
  IVP U55 ( .A(B[16]), .Z(n3) );
  IVP U56 ( .A(A[6]), .Z(n28) );
  IVP U57 ( .A(A[7]), .Z(n27) );
  IVP U58 ( .A(A[8]), .Z(n26) );
  IVP U59 ( .A(A[9]), .Z(n25) );
  IVP U60 ( .A(A[10]), .Z(n24) );
  IVP U61 ( .A(A[11]), .Z(n23) );
  IVP U62 ( .A(A[12]), .Z(n22) );
  IVP U63 ( .A(A[13]), .Z(n21) );
  IVP U64 ( .A(A[14]), .Z(n20) );
  AN2P U65 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A2[14] ) );
  AN2P U66 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A2[16] ) );
  AN2P U67 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A2[17] ) );
  AN2P U68 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A2[18] ) );
  AN2P U69 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A2[19] ) );
  AN2P U70 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A2[20] ) );
  AN2P U71 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A2[21] ) );
  AN2P U72 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A2[22] ) );
  AN2P U73 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A2[23] ) );
  AN2P U74 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A2[24] ) );
  AN2P U75 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A2[25] ) );
  AN2P U76 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A2[26] ) );
  AN2P U77 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A2[27] ) );
  AN2P U78 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A2[28] ) );
  AN2P U79 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A2[29] ) );
  AN2P U80 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U81 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U82 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U83 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U84 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U85 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U86 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U87 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U88 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U89 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U90 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U91 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U92 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U93 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U94 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U95 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A2[15] ) );
  NR2 U97 ( .A(n25), .B(n10), .Z(\ab[9][9] ) );
  NR2 U98 ( .A(n25), .B(n11), .Z(\ab[9][8] ) );
  NR2 U99 ( .A(n25), .B(n12), .Z(\ab[9][7] ) );
  NR2 U100 ( .A(n25), .B(n13), .Z(\ab[9][6] ) );
  NR2 U101 ( .A(n25), .B(n14), .Z(\ab[9][5] ) );
  NR2 U102 ( .A(n25), .B(n15), .Z(\ab[9][4] ) );
  NR2 U103 ( .A(n25), .B(n16), .Z(\ab[9][3] ) );
  NR2 U104 ( .A(n25), .B(n17), .Z(\ab[9][2] ) );
  NR2 U105 ( .A(n25), .B(n18), .Z(\ab[9][1] ) );
  NR2 U106 ( .A(n25), .B(n3), .Z(\ab[9][16] ) );
  NR2 U107 ( .A(n25), .B(n4), .Z(\ab[9][15] ) );
  NR2 U108 ( .A(n25), .B(n5), .Z(\ab[9][14] ) );
  NR2 U109 ( .A(n25), .B(n6), .Z(\ab[9][13] ) );
  NR2 U110 ( .A(n25), .B(n7), .Z(\ab[9][12] ) );
  NR2 U111 ( .A(n25), .B(n8), .Z(\ab[9][11] ) );
  NR2 U112 ( .A(n25), .B(n9), .Z(\ab[9][10] ) );
  NR2 U113 ( .A(n25), .B(n19), .Z(\ab[9][0] ) );
  NR2 U114 ( .A(n10), .B(n26), .Z(\ab[8][9] ) );
  NR2 U115 ( .A(n11), .B(n26), .Z(\ab[8][8] ) );
  NR2 U116 ( .A(n12), .B(n26), .Z(\ab[8][7] ) );
  NR2 U117 ( .A(n13), .B(n26), .Z(\ab[8][6] ) );
  NR2 U118 ( .A(n14), .B(n26), .Z(\ab[8][5] ) );
  NR2 U119 ( .A(n15), .B(n26), .Z(\ab[8][4] ) );
  NR2 U120 ( .A(n16), .B(n26), .Z(\ab[8][3] ) );
  NR2 U121 ( .A(n17), .B(n26), .Z(\ab[8][2] ) );
  NR2 U122 ( .A(n18), .B(n26), .Z(\ab[8][1] ) );
  NR2 U123 ( .A(n3), .B(n26), .Z(\ab[8][16] ) );
  NR2 U124 ( .A(n4), .B(n26), .Z(\ab[8][15] ) );
  NR2 U125 ( .A(n5), .B(n26), .Z(\ab[8][14] ) );
  NR2 U126 ( .A(n6), .B(n26), .Z(\ab[8][13] ) );
  NR2 U127 ( .A(n7), .B(n26), .Z(\ab[8][12] ) );
  NR2 U128 ( .A(n8), .B(n26), .Z(\ab[8][11] ) );
  NR2 U129 ( .A(n9), .B(n26), .Z(\ab[8][10] ) );
  NR2 U130 ( .A(n19), .B(n26), .Z(\ab[8][0] ) );
  NR2 U131 ( .A(n10), .B(n27), .Z(\ab[7][9] ) );
  NR2 U132 ( .A(n11), .B(n27), .Z(\ab[7][8] ) );
  NR2 U133 ( .A(n12), .B(n27), .Z(\ab[7][7] ) );
  NR2 U134 ( .A(n13), .B(n27), .Z(\ab[7][6] ) );
  NR2 U135 ( .A(n14), .B(n27), .Z(\ab[7][5] ) );
  NR2 U136 ( .A(n15), .B(n27), .Z(\ab[7][4] ) );
  NR2 U137 ( .A(n16), .B(n27), .Z(\ab[7][3] ) );
  NR2 U138 ( .A(n17), .B(n27), .Z(\ab[7][2] ) );
  NR2 U139 ( .A(n18), .B(n27), .Z(\ab[7][1] ) );
  NR2 U140 ( .A(n3), .B(n27), .Z(\ab[7][16] ) );
  NR2 U141 ( .A(n4), .B(n27), .Z(\ab[7][15] ) );
  NR2 U142 ( .A(n5), .B(n27), .Z(\ab[7][14] ) );
  NR2 U143 ( .A(n6), .B(n27), .Z(\ab[7][13] ) );
  NR2 U144 ( .A(n7), .B(n27), .Z(\ab[7][12] ) );
  NR2 U145 ( .A(n8), .B(n27), .Z(\ab[7][11] ) );
  NR2 U146 ( .A(n9), .B(n27), .Z(\ab[7][10] ) );
  NR2 U147 ( .A(n19), .B(n27), .Z(\ab[7][0] ) );
  NR2 U148 ( .A(n10), .B(n28), .Z(\ab[6][9] ) );
  NR2 U149 ( .A(n11), .B(n28), .Z(\ab[6][8] ) );
  NR2 U150 ( .A(n12), .B(n28), .Z(\ab[6][7] ) );
  NR2 U151 ( .A(n13), .B(n28), .Z(\ab[6][6] ) );
  NR2 U152 ( .A(n14), .B(n28), .Z(\ab[6][5] ) );
  NR2 U153 ( .A(n15), .B(n28), .Z(\ab[6][4] ) );
  NR2 U154 ( .A(n16), .B(n28), .Z(\ab[6][3] ) );
  NR2 U155 ( .A(n17), .B(n28), .Z(\ab[6][2] ) );
  NR2 U156 ( .A(n18), .B(n28), .Z(\ab[6][1] ) );
  NR2 U157 ( .A(n3), .B(n28), .Z(\ab[6][16] ) );
  NR2 U158 ( .A(n4), .B(n28), .Z(\ab[6][15] ) );
  NR2 U159 ( .A(n5), .B(n28), .Z(\ab[6][14] ) );
  NR2 U160 ( .A(n6), .B(n28), .Z(\ab[6][13] ) );
  NR2 U161 ( .A(n7), .B(n28), .Z(\ab[6][12] ) );
  NR2 U162 ( .A(n8), .B(n28), .Z(\ab[6][11] ) );
  NR2 U163 ( .A(n9), .B(n28), .Z(\ab[6][10] ) );
  NR2 U164 ( .A(n19), .B(n28), .Z(\ab[6][0] ) );
  NR2 U165 ( .A(n10), .B(n29), .Z(\ab[5][9] ) );
  NR2 U166 ( .A(n11), .B(n29), .Z(\ab[5][8] ) );
  NR2 U167 ( .A(n12), .B(n29), .Z(\ab[5][7] ) );
  NR2 U168 ( .A(n13), .B(n29), .Z(\ab[5][6] ) );
  NR2 U169 ( .A(n14), .B(n29), .Z(\ab[5][5] ) );
  NR2 U170 ( .A(n15), .B(n29), .Z(\ab[5][4] ) );
  NR2 U171 ( .A(n16), .B(n29), .Z(\ab[5][3] ) );
  NR2 U172 ( .A(n17), .B(n29), .Z(\ab[5][2] ) );
  NR2 U173 ( .A(n18), .B(n29), .Z(\ab[5][1] ) );
  NR2 U174 ( .A(n3), .B(n29), .Z(\ab[5][16] ) );
  NR2 U175 ( .A(n4), .B(n29), .Z(\ab[5][15] ) );
  NR2 U176 ( .A(n5), .B(n29), .Z(\ab[5][14] ) );
  NR2 U177 ( .A(n6), .B(n29), .Z(\ab[5][13] ) );
  NR2 U178 ( .A(n7), .B(n29), .Z(\ab[5][12] ) );
  NR2 U179 ( .A(n8), .B(n29), .Z(\ab[5][11] ) );
  NR2 U180 ( .A(n9), .B(n29), .Z(\ab[5][10] ) );
  NR2 U181 ( .A(n19), .B(n29), .Z(\ab[5][0] ) );
  NR2 U182 ( .A(n10), .B(n30), .Z(\ab[4][9] ) );
  NR2 U183 ( .A(n11), .B(n30), .Z(\ab[4][8] ) );
  NR2 U184 ( .A(n12), .B(n30), .Z(\ab[4][7] ) );
  NR2 U185 ( .A(n13), .B(n30), .Z(\ab[4][6] ) );
  NR2 U186 ( .A(n14), .B(n30), .Z(\ab[4][5] ) );
  NR2 U187 ( .A(n15), .B(n30), .Z(\ab[4][4] ) );
  NR2 U188 ( .A(n16), .B(n30), .Z(\ab[4][3] ) );
  NR2 U189 ( .A(n17), .B(n30), .Z(\ab[4][2] ) );
  NR2 U190 ( .A(n18), .B(n30), .Z(\ab[4][1] ) );
  NR2 U191 ( .A(n3), .B(n30), .Z(\ab[4][16] ) );
  NR2 U192 ( .A(n4), .B(n30), .Z(\ab[4][15] ) );
  NR2 U193 ( .A(n5), .B(n30), .Z(\ab[4][14] ) );
  NR2 U194 ( .A(n6), .B(n30), .Z(\ab[4][13] ) );
  NR2 U195 ( .A(n7), .B(n30), .Z(\ab[4][12] ) );
  NR2 U196 ( .A(n8), .B(n30), .Z(\ab[4][11] ) );
  NR2 U197 ( .A(n9), .B(n30), .Z(\ab[4][10] ) );
  NR2 U198 ( .A(n19), .B(n30), .Z(\ab[4][0] ) );
  NR2 U199 ( .A(n10), .B(n31), .Z(\ab[3][9] ) );
  NR2 U200 ( .A(n11), .B(n31), .Z(\ab[3][8] ) );
  NR2 U201 ( .A(n12), .B(n31), .Z(\ab[3][7] ) );
  NR2 U202 ( .A(n13), .B(n31), .Z(\ab[3][6] ) );
  NR2 U203 ( .A(n14), .B(n31), .Z(\ab[3][5] ) );
  NR2 U204 ( .A(n15), .B(n31), .Z(\ab[3][4] ) );
  NR2 U205 ( .A(n16), .B(n31), .Z(\ab[3][3] ) );
  NR2 U206 ( .A(n17), .B(n31), .Z(\ab[3][2] ) );
  NR2 U207 ( .A(n18), .B(n31), .Z(\ab[3][1] ) );
  NR2 U208 ( .A(n3), .B(n31), .Z(\ab[3][16] ) );
  NR2 U209 ( .A(n4), .B(n31), .Z(\ab[3][15] ) );
  NR2 U210 ( .A(n5), .B(n31), .Z(\ab[3][14] ) );
  NR2 U211 ( .A(n6), .B(n31), .Z(\ab[3][13] ) );
  NR2 U212 ( .A(n7), .B(n31), .Z(\ab[3][12] ) );
  NR2 U213 ( .A(n8), .B(n31), .Z(\ab[3][11] ) );
  NR2 U214 ( .A(n9), .B(n31), .Z(\ab[3][10] ) );
  NR2 U215 ( .A(n19), .B(n31), .Z(\ab[3][0] ) );
  NR2 U216 ( .A(n10), .B(n32), .Z(\ab[2][9] ) );
  NR2 U217 ( .A(n11), .B(n32), .Z(\ab[2][8] ) );
  NR2 U218 ( .A(n12), .B(n32), .Z(\ab[2][7] ) );
  NR2 U219 ( .A(n13), .B(n32), .Z(\ab[2][6] ) );
  NR2 U220 ( .A(n14), .B(n32), .Z(\ab[2][5] ) );
  NR2 U221 ( .A(n15), .B(n32), .Z(\ab[2][4] ) );
  NR2 U222 ( .A(n16), .B(n32), .Z(\ab[2][3] ) );
  NR2 U223 ( .A(n17), .B(n32), .Z(\ab[2][2] ) );
  NR2 U224 ( .A(n18), .B(n32), .Z(\ab[2][1] ) );
  NR2 U225 ( .A(n3), .B(n32), .Z(\ab[2][16] ) );
  NR2 U226 ( .A(n4), .B(n32), .Z(\ab[2][15] ) );
  NR2 U227 ( .A(n5), .B(n32), .Z(\ab[2][14] ) );
  NR2 U228 ( .A(n6), .B(n32), .Z(\ab[2][13] ) );
  NR2 U229 ( .A(n7), .B(n32), .Z(\ab[2][12] ) );
  NR2 U230 ( .A(n8), .B(n32), .Z(\ab[2][11] ) );
  NR2 U231 ( .A(n9), .B(n32), .Z(\ab[2][10] ) );
  NR2 U232 ( .A(n19), .B(n32), .Z(\ab[2][0] ) );
  NR2 U233 ( .A(n10), .B(n33), .Z(\ab[1][9] ) );
  NR2 U234 ( .A(n11), .B(n33), .Z(\ab[1][8] ) );
  NR2 U235 ( .A(n12), .B(n33), .Z(\ab[1][7] ) );
  NR2 U236 ( .A(n13), .B(n33), .Z(\ab[1][6] ) );
  NR2 U237 ( .A(n14), .B(n33), .Z(\ab[1][5] ) );
  NR2 U238 ( .A(n15), .B(n33), .Z(\ab[1][4] ) );
  NR2 U239 ( .A(n16), .B(n33), .Z(\ab[1][3] ) );
  NR2 U240 ( .A(n17), .B(n33), .Z(\ab[1][2] ) );
  NR2 U241 ( .A(n3), .B(n33), .Z(\ab[1][16] ) );
  NR2 U242 ( .A(n4), .B(n33), .Z(\ab[1][15] ) );
  NR2 U243 ( .A(n5), .B(n33), .Z(\ab[1][14] ) );
  NR2 U244 ( .A(n6), .B(n33), .Z(\ab[1][13] ) );
  NR2 U245 ( .A(n7), .B(n33), .Z(\ab[1][12] ) );
  NR2 U246 ( .A(n8), .B(n33), .Z(\ab[1][11] ) );
  NR2 U247 ( .A(n9), .B(n33), .Z(\ab[1][10] ) );
  NR2 U248 ( .A(n10), .B(n20), .Z(\ab[14][9] ) );
  NR2 U249 ( .A(n11), .B(n20), .Z(\ab[14][8] ) );
  NR2 U250 ( .A(n12), .B(n20), .Z(\ab[14][7] ) );
  NR2 U251 ( .A(n13), .B(n20), .Z(\ab[14][6] ) );
  NR2 U252 ( .A(n14), .B(n20), .Z(\ab[14][5] ) );
  NR2 U253 ( .A(n15), .B(n20), .Z(\ab[14][4] ) );
  NR2 U254 ( .A(n16), .B(n20), .Z(\ab[14][3] ) );
  NR2 U255 ( .A(n17), .B(n20), .Z(\ab[14][2] ) );
  NR2 U256 ( .A(n18), .B(n20), .Z(\ab[14][1] ) );
  NR2 U257 ( .A(n3), .B(n20), .Z(\ab[14][16] ) );
  NR2 U258 ( .A(n4), .B(n20), .Z(\ab[14][15] ) );
  NR2 U259 ( .A(n5), .B(n20), .Z(\ab[14][14] ) );
  NR2 U260 ( .A(n6), .B(n20), .Z(\ab[14][13] ) );
  NR2 U261 ( .A(n7), .B(n20), .Z(\ab[14][12] ) );
  NR2 U262 ( .A(n8), .B(n20), .Z(\ab[14][11] ) );
  NR2 U263 ( .A(n9), .B(n20), .Z(\ab[14][10] ) );
  NR2 U264 ( .A(n19), .B(n20), .Z(\ab[14][0] ) );
  NR2 U265 ( .A(n10), .B(n21), .Z(\ab[13][9] ) );
  NR2 U266 ( .A(n11), .B(n21), .Z(\ab[13][8] ) );
  NR2 U267 ( .A(n12), .B(n21), .Z(\ab[13][7] ) );
  NR2 U268 ( .A(n13), .B(n21), .Z(\ab[13][6] ) );
  NR2 U269 ( .A(n14), .B(n21), .Z(\ab[13][5] ) );
  NR2 U270 ( .A(n15), .B(n21), .Z(\ab[13][4] ) );
  NR2 U271 ( .A(n16), .B(n21), .Z(\ab[13][3] ) );
  NR2 U272 ( .A(n17), .B(n21), .Z(\ab[13][2] ) );
  NR2 U273 ( .A(n18), .B(n21), .Z(\ab[13][1] ) );
  NR2 U274 ( .A(n3), .B(n21), .Z(\ab[13][16] ) );
  NR2 U275 ( .A(n4), .B(n21), .Z(\ab[13][15] ) );
  NR2 U276 ( .A(n5), .B(n21), .Z(\ab[13][14] ) );
  NR2 U277 ( .A(n6), .B(n21), .Z(\ab[13][13] ) );
  NR2 U278 ( .A(n7), .B(n21), .Z(\ab[13][12] ) );
  NR2 U279 ( .A(n8), .B(n21), .Z(\ab[13][11] ) );
  NR2 U280 ( .A(n9), .B(n21), .Z(\ab[13][10] ) );
  NR2 U281 ( .A(n19), .B(n21), .Z(\ab[13][0] ) );
  NR2 U282 ( .A(n10), .B(n22), .Z(\ab[12][9] ) );
  NR2 U283 ( .A(n11), .B(n22), .Z(\ab[12][8] ) );
  NR2 U284 ( .A(n12), .B(n22), .Z(\ab[12][7] ) );
  NR2 U285 ( .A(n13), .B(n22), .Z(\ab[12][6] ) );
  NR2 U286 ( .A(n14), .B(n22), .Z(\ab[12][5] ) );
  NR2 U287 ( .A(n15), .B(n22), .Z(\ab[12][4] ) );
  NR2 U288 ( .A(n16), .B(n22), .Z(\ab[12][3] ) );
  NR2 U289 ( .A(n17), .B(n22), .Z(\ab[12][2] ) );
  NR2 U290 ( .A(n18), .B(n22), .Z(\ab[12][1] ) );
  NR2 U291 ( .A(n3), .B(n22), .Z(\ab[12][16] ) );
  NR2 U292 ( .A(n4), .B(n22), .Z(\ab[12][15] ) );
  NR2 U293 ( .A(n5), .B(n22), .Z(\ab[12][14] ) );
  NR2 U294 ( .A(n6), .B(n22), .Z(\ab[12][13] ) );
  NR2 U295 ( .A(n7), .B(n22), .Z(\ab[12][12] ) );
  NR2 U296 ( .A(n8), .B(n22), .Z(\ab[12][11] ) );
  NR2 U297 ( .A(n9), .B(n22), .Z(\ab[12][10] ) );
  NR2 U298 ( .A(n19), .B(n22), .Z(\ab[12][0] ) );
  NR2 U299 ( .A(n10), .B(n23), .Z(\ab[11][9] ) );
  NR2 U300 ( .A(n11), .B(n23), .Z(\ab[11][8] ) );
  NR2 U301 ( .A(n12), .B(n23), .Z(\ab[11][7] ) );
  NR2 U302 ( .A(n13), .B(n23), .Z(\ab[11][6] ) );
  NR2 U303 ( .A(n14), .B(n23), .Z(\ab[11][5] ) );
  NR2 U304 ( .A(n15), .B(n23), .Z(\ab[11][4] ) );
  NR2 U305 ( .A(n16), .B(n23), .Z(\ab[11][3] ) );
  NR2 U306 ( .A(n17), .B(n23), .Z(\ab[11][2] ) );
  NR2 U307 ( .A(n18), .B(n23), .Z(\ab[11][1] ) );
  NR2 U308 ( .A(n3), .B(n23), .Z(\ab[11][16] ) );
  NR2 U309 ( .A(n4), .B(n23), .Z(\ab[11][15] ) );
  NR2 U310 ( .A(n5), .B(n23), .Z(\ab[11][14] ) );
  NR2 U311 ( .A(n6), .B(n23), .Z(\ab[11][13] ) );
  NR2 U312 ( .A(n7), .B(n23), .Z(\ab[11][12] ) );
  NR2 U313 ( .A(n8), .B(n23), .Z(\ab[11][11] ) );
  NR2 U314 ( .A(n9), .B(n23), .Z(\ab[11][10] ) );
  NR2 U315 ( .A(n19), .B(n23), .Z(\ab[11][0] ) );
  NR2 U316 ( .A(n10), .B(n24), .Z(\ab[10][9] ) );
  NR2 U317 ( .A(n11), .B(n24), .Z(\ab[10][8] ) );
  NR2 U318 ( .A(n12), .B(n24), .Z(\ab[10][7] ) );
  NR2 U319 ( .A(n13), .B(n24), .Z(\ab[10][6] ) );
  NR2 U320 ( .A(n14), .B(n24), .Z(\ab[10][5] ) );
  NR2 U321 ( .A(n15), .B(n24), .Z(\ab[10][4] ) );
  NR2 U322 ( .A(n16), .B(n24), .Z(\ab[10][3] ) );
  NR2 U323 ( .A(n17), .B(n24), .Z(\ab[10][2] ) );
  NR2 U324 ( .A(n18), .B(n24), .Z(\ab[10][1] ) );
  NR2 U325 ( .A(n3), .B(n24), .Z(\ab[10][16] ) );
  NR2 U326 ( .A(n4), .B(n24), .Z(\ab[10][15] ) );
  NR2 U327 ( .A(n5), .B(n24), .Z(\ab[10][14] ) );
  NR2 U328 ( .A(n6), .B(n24), .Z(\ab[10][13] ) );
  NR2 U329 ( .A(n7), .B(n24), .Z(\ab[10][12] ) );
  NR2 U330 ( .A(n8), .B(n24), .Z(\ab[10][11] ) );
  NR2 U331 ( .A(n9), .B(n24), .Z(\ab[10][10] ) );
  NR2 U332 ( .A(n19), .B(n24), .Z(\ab[10][0] ) );
  NR2 U333 ( .A(n10), .B(n34), .Z(\ab[0][9] ) );
  NR2 U334 ( .A(n11), .B(n34), .Z(\ab[0][8] ) );
  NR2 U335 ( .A(n12), .B(n34), .Z(\ab[0][7] ) );
  NR2 U336 ( .A(n13), .B(n34), .Z(\ab[0][6] ) );
  NR2 U337 ( .A(n14), .B(n34), .Z(\ab[0][5] ) );
  NR2 U338 ( .A(n15), .B(n34), .Z(\ab[0][4] ) );
  NR2 U339 ( .A(n16), .B(n34), .Z(\ab[0][3] ) );
  NR2 U340 ( .A(n17), .B(n34), .Z(\ab[0][2] ) );
  NR2 U341 ( .A(n3), .B(n34), .Z(\ab[0][16] ) );
  NR2 U342 ( .A(n4), .B(n34), .Z(\ab[0][15] ) );
  NR2 U343 ( .A(n5), .B(n34), .Z(\ab[0][14] ) );
  NR2 U344 ( .A(n6), .B(n34), .Z(\ab[0][13] ) );
  NR2 U345 ( .A(n7), .B(n34), .Z(\ab[0][12] ) );
  NR2 U346 ( .A(n8), .B(n34), .Z(\ab[0][11] ) );
  NR2 U347 ( .A(n9), .B(n34), .Z(\ab[0][10] ) );
  AN3 U348 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U349 ( .A(n33), .B(n18), .Z(\ab[1][1] ) );
endmodule


module AWGN ( clk, reset, Valid, X0_Out, X1_Out );
  output [15:0] X0_Out;
  output [15:0] X1_Out;
  input clk, reset;
  output Valid;
  wire   Valid0, Valid1, Valid2, Valid3, Valid4, Valid5, Valid6, Valid7,
         Valid8, Valid9, Valid10, Valid11, Valid12, Valid13, Valid14, Valid15,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535;
  wire   [31:0] Taus1;
  wire   [31:0] Taus2;
  wire   [47:0] LogIn;
  wire   [15:0] Angle;
  wire   [15:0] Sin2;
  wire   [15:0] Sin11;
  wire   [15:0] Cos2;
  wire   [15:0] Cos11;
  wire   [15:0] Sin3;
  wire   [15:0] Cos3;
  wire   [15:0] Sin4;
  wire   [15:0] Cos4;
  wire   [15:0] Sin5;
  wire   [15:0] Cos5;
  wire   [15:0] Sin6;
  wire   [15:0] Cos6;
  wire   [15:0] Sin7;
  wire   [15:0] Cos7;
  wire   [15:0] Sin8;
  wire   [15:0] Cos8;
  wire   [15:0] Sin1;
  wire   [15:0] Cos1;
  wire   [15:0] Sin;
  wire   [15:0] Cos;
  wire   [30:0] LogOut2;
  wire   [30:0] LogOut;
  wire   [15:0] X0;
  wire   [15:0] X1;
  wire   [16:0] SqrtOut;
  wire   [31:17] RegX0;
  wire   [31:17] RegX1;
  wire   [15:0] X01;
  wire   [15:0] X11;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34;

  FDS2LP \LogIn_reg[47]  ( .CR(1'b1), .D(Taus1[31]), .LD(n490), .CP(clk), .Q(
        LogIn[47]) );
  FDS2LP \LogIn_reg[32]  ( .CR(1'b1), .D(Taus1[16]), .LD(n489), .CP(clk), .Q(
        LogIn[32]) );
  FDS2LP \LogIn_reg[26]  ( .CR(1'b1), .D(Taus1[10]), .LD(n489), .CP(clk), .Q(
        LogIn[26]) );
  FDS2LP \LogIn_reg[1]  ( .CR(1'b1), .D(Taus2[17]), .LD(n487), .CP(clk), .Q(
        LogIn[1]) );
  FDS2LP \LogIn_reg[0]  ( .CR(1'b1), .D(Taus2[16]), .LD(n487), .CP(clk), .Q(
        LogIn[0]) );
  Taus_0 T1 ( .clk(clk), .reset(reset), .Tout(Taus1) );
  Taus_1 T2 ( .clk(clk), .reset(reset), .Tout(Taus2) );
  LOG_POLY L1 ( .clk(clk), .reset(reset), .LogIn(LogIn), .LogOut({LogOut[30:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  SQRT_POLY S1 ( .clk(clk), .reset(reset), .RootIn(LogOut2), .RootOut(SqrtOut)
         );
  SinBlock_0 SinInst1 ( .clk(clk), .reset(reset), .func(1'b0), .x(Angle), 
        .sinValue(Sin11) );
  SinBlock_1 CosInst1 ( .clk(clk), .reset(reset), .func(1'b1), .x(Angle), 
        .sinValue(Cos11) );
  AWGN_DW02_mult_1 mult_68 ( .A(Sin[14:0]), .B(SqrtOut), .TC(1'b0), .PRODUCT({
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17}) );
  AWGN_DW02_mult_0 mult_69 ( .A(Cos[14:0]), .B(SqrtOut), .TC(1'b0), .PRODUCT({
        N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, 
        N20, SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34}) );
  FD1P \LogIn_reg[27]  ( .D(n486), .CP(clk), .Q(LogIn[27]) );
  FD1P \LogIn_reg[2]  ( .D(n484), .CP(clk), .Q(LogIn[2]) );
  FDS2L \Angle_reg[15]  ( .CR(1'b1), .D(Taus2[15]), .LD(n529), .CP(clk), .Q(
        Angle[15]) );
  FDS2L \Sin_reg[14]  ( .CR(1'b1), .D(Sin1[14]), .LD(n506), .CP(clk), .Q(
        Sin[14]) );
  FDS2L \Cos_reg[14]  ( .CR(1'b1), .D(Cos1[14]), .LD(n505), .CP(clk), .Q(
        Cos[14]) );
  FDS2L \Sin_reg[13]  ( .CR(1'b1), .D(Sin1[13]), .LD(n506), .CP(clk), .Q(
        Sin[13]) );
  FDS2L \Cos_reg[13]  ( .CR(1'b1), .D(Cos1[13]), .LD(n505), .CP(clk), .Q(
        Cos[13]) );
  FDS2L \Sin_reg[12]  ( .CR(1'b1), .D(Sin1[12]), .LD(n506), .CP(clk), .Q(
        Sin[12]) );
  FDS2L \Cos_reg[12]  ( .CR(1'b1), .D(Cos1[12]), .LD(n505), .CP(clk), .Q(
        Cos[12]) );
  FDS2L \Sin_reg[11]  ( .CR(1'b1), .D(Sin1[11]), .LD(n506), .CP(clk), .Q(
        Sin[11]) );
  FDS2L \Cos_reg[11]  ( .CR(1'b1), .D(Cos1[11]), .LD(n505), .CP(clk), .Q(
        Cos[11]) );
  FDS2L \Sin_reg[10]  ( .CR(1'b1), .D(Sin1[10]), .LD(n506), .CP(clk), .Q(
        Sin[10]) );
  FDS2L \Cos_reg[10]  ( .CR(1'b1), .D(Cos1[10]), .LD(n504), .CP(clk), .Q(
        Cos[10]) );
  FDS2L \Sin_reg[9]  ( .CR(1'b1), .D(Sin1[9]), .LD(n506), .CP(clk), .Q(Sin[9])
         );
  FDS2L \Cos_reg[9]  ( .CR(1'b1), .D(Cos1[9]), .LD(n504), .CP(clk), .Q(Cos[9])
         );
  FDS2L \LogOut2_reg[24]  ( .CR(1'b1), .D(LogOut[24]), .LD(n503), .CP(clk), 
        .Q(LogOut2[24]) );
  FDS2L \Sin_reg[8]  ( .CR(1'b1), .D(Sin1[8]), .LD(n506), .CP(clk), .Q(Sin[8])
         );
  FDS2L \Cos_reg[8]  ( .CR(1'b1), .D(Cos1[8]), .LD(n504), .CP(clk), .Q(Cos[8])
         );
  FDS2L \LogOut2_reg[23]  ( .CR(1'b1), .D(LogOut[23]), .LD(n503), .CP(clk), 
        .Q(LogOut2[23]) );
  FDS2L \LogOut2_reg[22]  ( .CR(1'b1), .D(LogOut[22]), .LD(n503), .CP(clk), 
        .Q(LogOut2[22]) );
  FDS2L \Sin_reg[7]  ( .CR(1'b1), .D(Sin1[7]), .LD(n506), .CP(clk), .Q(Sin[7])
         );
  FDS2L \Cos_reg[7]  ( .CR(1'b1), .D(Cos1[7]), .LD(n504), .CP(clk), .Q(Cos[7])
         );
  FDS2L \LogOut2_reg[21]  ( .CR(1'b1), .D(LogOut[21]), .LD(n503), .CP(clk), 
        .Q(LogOut2[21]) );
  FDS2L \Angle_reg[7]  ( .CR(1'b1), .D(Taus2[7]), .LD(n528), .CP(clk), .Q(
        Angle[7]) );
  FDS2L \Angle_reg[6]  ( .CR(1'b1), .D(Taus2[6]), .LD(n528), .CP(clk), .Q(
        Angle[6]) );
  FDS2L \Sin_reg[6]  ( .CR(1'b1), .D(Sin1[6]), .LD(n505), .CP(clk), .Q(Sin[6])
         );
  FDS2L \Cos_reg[6]  ( .CR(1'b1), .D(Cos1[6]), .LD(n504), .CP(clk), .Q(Cos[6])
         );
  FDS2L \Angle_reg[0]  ( .CR(1'b1), .D(Taus2[0]), .LD(n528), .CP(clk), .Q(
        Angle[0]) );
  FDS2L \LogOut2_reg[20]  ( .CR(1'b1), .D(LogOut[20]), .LD(n503), .CP(clk), 
        .Q(LogOut2[20]) );
  FDS2L \Angle_reg[5]  ( .CR(1'b1), .D(Taus2[5]), .LD(n528), .CP(clk), .Q(
        Angle[5]) );
  FDS2L \LogOut2_reg[19]  ( .CR(1'b1), .D(LogOut[19]), .LD(n503), .CP(clk), 
        .Q(LogOut2[19]) );
  FDS2L \LogOut2_reg[18]  ( .CR(1'b1), .D(LogOut[18]), .LD(n503), .CP(clk), 
        .Q(LogOut2[18]) );
  FDS2L \LogOut2_reg[17]  ( .CR(1'b1), .D(LogOut[17]), .LD(n502), .CP(clk), 
        .Q(LogOut2[17]) );
  FDS2L \Angle_reg[4]  ( .CR(1'b1), .D(Taus2[4]), .LD(n528), .CP(clk), .Q(
        Angle[4]) );
  FDS2L \Angle_reg[3]  ( .CR(1'b1), .D(Taus2[3]), .LD(n528), .CP(clk), .Q(
        Angle[3]) );
  FDS2L \Angle_reg[2]  ( .CR(1'b1), .D(Taus2[2]), .LD(n528), .CP(clk), .Q(
        Angle[2]) );
  FDS2L \Angle_reg[1]  ( .CR(1'b1), .D(Taus2[1]), .LD(n528), .CP(clk), .Q(
        Angle[1]) );
  FDS2L \LogOut2_reg[16]  ( .CR(1'b1), .D(LogOut[16]), .LD(n502), .CP(clk), 
        .Q(LogOut2[16]) );
  FDS2L \Sin_reg[5]  ( .CR(1'b1), .D(Sin1[5]), .LD(n505), .CP(clk), .Q(Sin[5])
         );
  FDS2L \Cos_reg[5]  ( .CR(1'b1), .D(Cos1[5]), .LD(n504), .CP(clk), .Q(Cos[5])
         );
  FDS2L \LogOut2_reg[15]  ( .CR(1'b1), .D(LogOut[15]), .LD(n502), .CP(clk), 
        .Q(LogOut2[15]) );
  FDS2L \Angle_reg[14]  ( .CR(1'b1), .D(Taus2[14]), .LD(n529), .CP(clk), .Q(
        Angle[14]) );
  FDS2L \LogOut2_reg[14]  ( .CR(1'b1), .D(LogOut[14]), .LD(n502), .CP(clk), 
        .Q(LogOut2[14]) );
  FDS2L \LogOut2_reg[13]  ( .CR(1'b1), .D(LogOut[13]), .LD(n502), .CP(clk), 
        .Q(LogOut2[13]) );
  FDS2L \LogOut2_reg[12]  ( .CR(1'b1), .D(LogOut[12]), .LD(n502), .CP(clk), 
        .Q(LogOut2[12]) );
  FDS2L \LogOut2_reg[11]  ( .CR(1'b1), .D(LogOut[11]), .LD(n502), .CP(clk), 
        .Q(LogOut2[11]) );
  FDS2L \LogOut2_reg[10]  ( .CR(1'b1), .D(LogOut[10]), .LD(n502), .CP(clk), 
        .Q(LogOut2[10]) );
  FDS2L \LogOut2_reg[9]  ( .CR(1'b1), .D(LogOut[9]), .LD(n502), .CP(clk), .Q(
        LogOut2[9]) );
  FDS2L \LogOut2_reg[8]  ( .CR(1'b1), .D(LogOut[8]), .LD(n502), .CP(clk), .Q(
        LogOut2[8]) );
  FDS2L \LogOut2_reg[7]  ( .CR(1'b1), .D(LogOut[7]), .LD(n502), .CP(clk), .Q(
        LogOut2[7]) );
  FDS2L \Sin_reg[4]  ( .CR(1'b1), .D(Sin1[4]), .LD(n505), .CP(clk), .Q(Sin[4])
         );
  FDS2L \Cos_reg[4]  ( .CR(1'b1), .D(Cos1[4]), .LD(n504), .CP(clk), .Q(Cos[4])
         );
  FDS2L \Angle_reg[11]  ( .CR(1'b1), .D(Taus2[11]), .LD(n529), .CP(clk), .Q(
        Angle[11]) );
  FDS2L \LogOut2_reg[6]  ( .CR(1'b1), .D(LogOut[6]), .LD(n502), .CP(clk), .Q(
        LogOut2[6]) );
  FDS2L \Sin_reg[3]  ( .CR(1'b1), .D(Sin1[3]), .LD(n505), .CP(clk), .Q(Sin[3])
         );
  FDS2L \Cos_reg[3]  ( .CR(1'b1), .D(Cos1[3]), .LD(n504), .CP(clk), .Q(Cos[3])
         );
  FDS2L \Angle_reg[12]  ( .CR(1'b1), .D(Taus2[12]), .LD(n529), .CP(clk), .Q(
        Angle[12]) );
  FDS2L \Angle_reg[13]  ( .CR(1'b1), .D(Taus2[13]), .LD(n529), .CP(clk), .Q(
        Angle[13]) );
  FDS2L \LogOut2_reg[5]  ( .CR(1'b1), .D(LogOut[5]), .LD(n501), .CP(clk), .Q(
        LogOut2[5]) );
  FDS2L \LogOut2_reg[0]  ( .CR(1'b1), .D(1'b0), .LD(n501), .CP(clk), .Q(
        LogOut2[0]) );
  FDS2L \LogOut2_reg[4]  ( .CR(1'b1), .D(LogOut[4]), .LD(n501), .CP(clk), .Q(
        LogOut2[4]) );
  FDS2L \LogOut2_reg[3]  ( .CR(1'b1), .D(LogOut[3]), .LD(n501), .CP(clk), .Q(
        LogOut2[3]) );
  FDS2L \LogOut2_reg[2]  ( .CR(1'b1), .D(LogOut[2]), .LD(n501), .CP(clk), .Q(
        LogOut2[2]) );
  FDS2L \LogOut2_reg[1]  ( .CR(1'b1), .D(LogOut[1]), .LD(n501), .CP(clk), .Q(
        LogOut2[1]) );
  FDS2L \Sin_reg[2]  ( .CR(1'b1), .D(Sin1[2]), .LD(n505), .CP(clk), .Q(Sin[2])
         );
  FDS2L \Cos_reg[2]  ( .CR(1'b1), .D(Cos1[2]), .LD(n504), .CP(clk), .Q(Cos[2])
         );
  FDS2L \Sin_reg[0]  ( .CR(1'b1), .D(Sin1[0]), .LD(n505), .CP(clk), .Q(Sin[0])
         );
  FDS2L \Cos_reg[0]  ( .CR(1'b1), .D(Cos1[0]), .LD(n504), .CP(clk), .Q(Cos[0])
         );
  FDS2L \Angle_reg[9]  ( .CR(1'b1), .D(Taus2[9]), .LD(n528), .CP(clk), .Q(
        Angle[9]) );
  FDS2L \Angle_reg[8]  ( .CR(1'b1), .D(Taus2[8]), .LD(n528), .CP(clk), .Q(
        Angle[8]) );
  FDS2L \Sin_reg[1]  ( .CR(1'b1), .D(Sin1[1]), .LD(n505), .CP(clk), .Q(Sin[1])
         );
  FDS2L \Cos_reg[1]  ( .CR(1'b1), .D(Cos1[1]), .LD(n504), .CP(clk), .Q(Cos[1])
         );
  FDS2L \Angle_reg[10]  ( .CR(1'b1), .D(Taus2[10]), .LD(n528), .CP(clk), .Q(
        Angle[10]) );
  FDS2L \LogOut2_reg[29]  ( .CR(1'b1), .D(LogOut[29]), .LD(n503), .CP(clk), 
        .Q(LogOut2[29]) );
  FDS2L \LogOut2_reg[28]  ( .CR(1'b1), .D(LogOut[28]), .LD(n503), .CP(clk), 
        .Q(LogOut2[28]) );
  FDS2L \LogOut2_reg[30]  ( .CR(1'b1), .D(LogOut[30]), .LD(n504), .CP(clk), 
        .Q(LogOut2[30]) );
  FDS2L \LogOut2_reg[25]  ( .CR(1'b1), .D(LogOut[25]), .LD(n503), .CP(clk), 
        .Q(LogOut2[25]) );
  FDS2L \LogOut2_reg[27]  ( .CR(1'b1), .D(LogOut[27]), .LD(n503), .CP(clk), 
        .Q(LogOut2[27]) );
  FDS2L \LogOut2_reg[26]  ( .CR(1'b1), .D(LogOut[26]), .LD(n503), .CP(clk), 
        .Q(LogOut2[26]) );
  FDS2 Valid_reg ( .CR(Valid15), .D(n529), .CP(clk), .Q(Valid) );
  FDS2 \X1_Out_reg[15]  ( .CR(X11[15]), .D(n494), .CP(clk), .Q(X1_Out[15]) );
  FDS2 \X1_Out_reg[14]  ( .CR(X11[14]), .D(n494), .CP(clk), .Q(X1_Out[14]) );
  FDS2 \X1_Out_reg[13]  ( .CR(X11[13]), .D(n494), .CP(clk), .Q(X1_Out[13]) );
  FDS2 \X1_Out_reg[12]  ( .CR(X11[12]), .D(n494), .CP(clk), .Q(X1_Out[12]) );
  FDS2 \X1_Out_reg[11]  ( .CR(X11[11]), .D(n494), .CP(clk), .Q(X1_Out[11]) );
  FDS2 \X1_Out_reg[10]  ( .CR(X11[10]), .D(n494), .CP(clk), .Q(X1_Out[10]) );
  FDS2 \X1_Out_reg[9]  ( .CR(X11[9]), .D(n493), .CP(clk), .Q(X1_Out[9]) );
  FDS2 \X1_Out_reg[8]  ( .CR(X11[8]), .D(n493), .CP(clk), .Q(X1_Out[8]) );
  FDS2 \X1_Out_reg[7]  ( .CR(X11[7]), .D(n493), .CP(clk), .Q(X1_Out[7]) );
  FDS2 \X1_Out_reg[6]  ( .CR(X11[6]), .D(n493), .CP(clk), .Q(X1_Out[6]) );
  FDS2 \X1_Out_reg[5]  ( .CR(X11[5]), .D(n493), .CP(clk), .Q(X1_Out[5]) );
  FDS2 \X1_Out_reg[4]  ( .CR(X11[4]), .D(n493), .CP(clk), .Q(X1_Out[4]) );
  FDS2 \X1_Out_reg[3]  ( .CR(X11[3]), .D(n492), .CP(clk), .Q(X1_Out[3]) );
  FDS2 \X1_Out_reg[2]  ( .CR(X11[2]), .D(n492), .CP(clk), .Q(X1_Out[2]) );
  FDS2 \X1_Out_reg[1]  ( .CR(X11[1]), .D(n492), .CP(clk), .Q(X1_Out[1]) );
  FDS2 \X1_Out_reg[0]  ( .CR(X11[0]), .D(n492), .CP(clk), .Q(X1_Out[0]) );
  FDS2 \X0_Out_reg[15]  ( .CR(X01[15]), .D(n492), .CP(clk), .Q(X0_Out[15]) );
  FDS2 \X0_Out_reg[14]  ( .CR(X01[14]), .D(n492), .CP(clk), .Q(X0_Out[14]) );
  FDS2 \X0_Out_reg[13]  ( .CR(X01[13]), .D(n492), .CP(clk), .Q(X0_Out[13]) );
  FDS2 \X0_Out_reg[12]  ( .CR(X01[12]), .D(n492), .CP(clk), .Q(X0_Out[12]) );
  FDS2 \X0_Out_reg[11]  ( .CR(X01[11]), .D(n491), .CP(clk), .Q(X0_Out[11]) );
  FDS2 \X0_Out_reg[10]  ( .CR(X01[10]), .D(n491), .CP(clk), .Q(X0_Out[10]) );
  FDS2 \X0_Out_reg[9]  ( .CR(X01[9]), .D(n491), .CP(clk), .Q(X0_Out[9]) );
  FDS2 \X0_Out_reg[8]  ( .CR(X01[8]), .D(n491), .CP(clk), .Q(X0_Out[8]) );
  FDS2 \X0_Out_reg[7]  ( .CR(X01[7]), .D(n491), .CP(clk), .Q(X0_Out[7]) );
  FDS2 \X0_Out_reg[6]  ( .CR(X01[6]), .D(n491), .CP(clk), .Q(X0_Out[6]) );
  FDS2 \X0_Out_reg[5]  ( .CR(X01[5]), .D(n491), .CP(clk), .Q(X0_Out[5]) );
  FDS2 \X0_Out_reg[4]  ( .CR(X01[4]), .D(n491), .CP(clk), .Q(X0_Out[4]) );
  FDS2 \X0_Out_reg[3]  ( .CR(X01[3]), .D(n491), .CP(clk), .Q(X0_Out[3]) );
  FDS2 \X0_Out_reg[2]  ( .CR(X01[2]), .D(n491), .CP(clk), .Q(X0_Out[2]) );
  FDS2 \X0_Out_reg[1]  ( .CR(X01[1]), .D(n491), .CP(clk), .Q(X0_Out[1]) );
  FDS2 \X0_Out_reg[0]  ( .CR(X01[0]), .D(n491), .CP(clk), .Q(X0_Out[0]) );
  FD1 Valid0_reg ( .D(n530), .CP(clk), .Q(Valid0) );
  FDS2 Valid1_reg ( .CR(Valid0), .D(n530), .CP(clk), .Q(Valid1) );
  FDS2 Valid2_reg ( .CR(Valid1), .D(n530), .CP(clk), .Q(Valid2) );
  FDS2 Valid3_reg ( .CR(Valid2), .D(n530), .CP(clk), .Q(Valid3) );
  FDS2 Valid4_reg ( .CR(Valid3), .D(n530), .CP(clk), .Q(Valid4) );
  FDS2 Valid5_reg ( .CR(Valid4), .D(n530), .CP(clk), .Q(Valid5) );
  FDS2 Valid6_reg ( .CR(Valid5), .D(n530), .CP(clk), .Q(Valid6) );
  FDS2 Valid7_reg ( .CR(Valid6), .D(n530), .CP(clk), .Q(Valid7) );
  FDS2 Valid8_reg ( .CR(Valid7), .D(n530), .CP(clk), .Q(Valid8) );
  FDS2 Valid9_reg ( .CR(Valid8), .D(n530), .CP(clk), .Q(Valid9) );
  FDS2 Valid10_reg ( .CR(Valid9), .D(n529), .CP(clk), .Q(Valid10) );
  FDS2 Valid11_reg ( .CR(Valid10), .D(n529), .CP(clk), .Q(Valid11) );
  FDS2 Valid12_reg ( .CR(Valid11), .D(n529), .CP(clk), .Q(Valid12) );
  FDS2 Valid13_reg ( .CR(Valid12), .D(n529), .CP(clk), .Q(Valid13) );
  FDS2 Valid14_reg ( .CR(Valid13), .D(n529), .CP(clk), .Q(Valid14) );
  FDS2 Valid15_reg ( .CR(Valid14), .D(n529), .CP(clk), .Q(Valid15) );
  FDS2L \Sin2_reg[15]  ( .CR(1'b1), .D(Sin11[15]), .LD(n528), .CP(clk), .Q(
        Sin2[15]) );
  FDS2L \Sin2_reg[14]  ( .CR(1'b1), .D(Sin11[14]), .LD(n527), .CP(clk), .Q(
        Sin2[14]) );
  FDS2L \Sin2_reg[13]  ( .CR(1'b1), .D(Sin11[13]), .LD(n527), .CP(clk), .Q(
        Sin2[13]) );
  FDS2L \Sin2_reg[12]  ( .CR(1'b1), .D(Sin11[12]), .LD(n527), .CP(clk), .Q(
        Sin2[12]) );
  FDS2L \Sin2_reg[11]  ( .CR(1'b1), .D(Sin11[11]), .LD(n527), .CP(clk), .Q(
        Sin2[11]) );
  FDS2L \Sin2_reg[10]  ( .CR(1'b1), .D(Sin11[10]), .LD(n527), .CP(clk), .Q(
        Sin2[10]) );
  FDS2L \Sin2_reg[9]  ( .CR(1'b1), .D(Sin11[9]), .LD(n527), .CP(clk), .Q(
        Sin2[9]) );
  FDS2L \Sin2_reg[8]  ( .CR(1'b1), .D(Sin11[8]), .LD(n527), .CP(clk), .Q(
        Sin2[8]) );
  FDS2L \Sin2_reg[7]  ( .CR(1'b1), .D(Sin11[7]), .LD(n527), .CP(clk), .Q(
        Sin2[7]) );
  FDS2L \Sin2_reg[6]  ( .CR(1'b1), .D(Sin11[6]), .LD(n527), .CP(clk), .Q(
        Sin2[6]) );
  FDS2L \Sin2_reg[5]  ( .CR(1'b1), .D(Sin11[5]), .LD(n527), .CP(clk), .Q(
        Sin2[5]) );
  FDS2L \Sin2_reg[4]  ( .CR(1'b1), .D(Sin11[4]), .LD(n527), .CP(clk), .Q(
        Sin2[4]) );
  FDS2L \Sin2_reg[3]  ( .CR(1'b1), .D(Sin11[3]), .LD(n527), .CP(clk), .Q(
        Sin2[3]) );
  FDS2L \Sin2_reg[2]  ( .CR(1'b1), .D(Sin11[2]), .LD(n526), .CP(clk), .Q(
        Sin2[2]) );
  FDS2L \Sin2_reg[1]  ( .CR(1'b1), .D(Sin11[1]), .LD(n526), .CP(clk), .Q(
        Sin2[1]) );
  FDS2L \Sin2_reg[0]  ( .CR(1'b1), .D(Sin11[0]), .LD(n526), .CP(clk), .Q(
        Sin2[0]) );
  FDS2L \Cos2_reg[15]  ( .CR(1'b1), .D(Cos11[15]), .LD(n526), .CP(clk), .Q(
        Cos2[15]) );
  FDS2L \Cos2_reg[14]  ( .CR(1'b1), .D(Cos11[14]), .LD(n526), .CP(clk), .Q(
        Cos2[14]) );
  FDS2L \Cos2_reg[13]  ( .CR(1'b1), .D(Cos11[13]), .LD(n526), .CP(clk), .Q(
        Cos2[13]) );
  FDS2L \Cos2_reg[12]  ( .CR(1'b1), .D(Cos11[12]), .LD(n526), .CP(clk), .Q(
        Cos2[12]) );
  FDS2L \Cos2_reg[11]  ( .CR(1'b1), .D(Cos11[11]), .LD(n526), .CP(clk), .Q(
        Cos2[11]) );
  FDS2L \Cos2_reg[10]  ( .CR(1'b1), .D(Cos11[10]), .LD(n526), .CP(clk), .Q(
        Cos2[10]) );
  FDS2L \Cos2_reg[9]  ( .CR(1'b1), .D(Cos11[9]), .LD(n526), .CP(clk), .Q(
        Cos2[9]) );
  FDS2L \Cos2_reg[8]  ( .CR(1'b1), .D(Cos11[8]), .LD(n526), .CP(clk), .Q(
        Cos2[8]) );
  FDS2L \Cos2_reg[7]  ( .CR(1'b1), .D(Cos11[7]), .LD(n526), .CP(clk), .Q(
        Cos2[7]) );
  FDS2L \Cos2_reg[6]  ( .CR(1'b1), .D(Cos11[6]), .LD(n525), .CP(clk), .Q(
        Cos2[6]) );
  FDS2L \Cos2_reg[5]  ( .CR(1'b1), .D(Cos11[5]), .LD(n525), .CP(clk), .Q(
        Cos2[5]) );
  FDS2L \Cos2_reg[4]  ( .CR(1'b1), .D(Cos11[4]), .LD(n525), .CP(clk), .Q(
        Cos2[4]) );
  FDS2L \Cos2_reg[3]  ( .CR(1'b1), .D(Cos11[3]), .LD(n525), .CP(clk), .Q(
        Cos2[3]) );
  FDS2L \Cos2_reg[2]  ( .CR(1'b1), .D(Cos11[2]), .LD(n525), .CP(clk), .Q(
        Cos2[2]) );
  FDS2L \Cos2_reg[1]  ( .CR(1'b1), .D(Cos11[1]), .LD(n525), .CP(clk), .Q(
        Cos2[1]) );
  FDS2L \Cos2_reg[0]  ( .CR(1'b1), .D(Cos11[0]), .LD(n525), .CP(clk), .Q(
        Cos2[0]) );
  FDS2L \Sin3_reg[15]  ( .CR(1'b1), .D(Sin2[15]), .LD(n525), .CP(clk), .Q(
        Sin3[15]) );
  FDS2L \Sin3_reg[14]  ( .CR(1'b1), .D(Sin2[14]), .LD(n525), .CP(clk), .Q(
        Sin3[14]) );
  FDS2L \Sin3_reg[13]  ( .CR(1'b1), .D(Sin2[13]), .LD(n525), .CP(clk), .Q(
        Sin3[13]) );
  FDS2L \Sin3_reg[12]  ( .CR(1'b1), .D(Sin2[12]), .LD(n525), .CP(clk), .Q(
        Sin3[12]) );
  FDS2L \Sin3_reg[11]  ( .CR(1'b1), .D(Sin2[11]), .LD(n525), .CP(clk), .Q(
        Sin3[11]) );
  FDS2L \Sin3_reg[10]  ( .CR(1'b1), .D(Sin2[10]), .LD(n524), .CP(clk), .Q(
        Sin3[10]) );
  FDS2L \Sin3_reg[9]  ( .CR(1'b1), .D(Sin2[9]), .LD(n524), .CP(clk), .Q(
        Sin3[9]) );
  FDS2L \Sin3_reg[8]  ( .CR(1'b1), .D(Sin2[8]), .LD(n524), .CP(clk), .Q(
        Sin3[8]) );
  FDS2L \Sin3_reg[7]  ( .CR(1'b1), .D(Sin2[7]), .LD(n524), .CP(clk), .Q(
        Sin3[7]) );
  FDS2L \Sin3_reg[6]  ( .CR(1'b1), .D(Sin2[6]), .LD(n524), .CP(clk), .Q(
        Sin3[6]) );
  FDS2L \Sin3_reg[5]  ( .CR(1'b1), .D(Sin2[5]), .LD(n524), .CP(clk), .Q(
        Sin3[5]) );
  FDS2L \Sin3_reg[4]  ( .CR(1'b1), .D(Sin2[4]), .LD(n524), .CP(clk), .Q(
        Sin3[4]) );
  FDS2L \Sin3_reg[3]  ( .CR(1'b1), .D(Sin2[3]), .LD(n524), .CP(clk), .Q(
        Sin3[3]) );
  FDS2L \Sin3_reg[2]  ( .CR(1'b1), .D(Sin2[2]), .LD(n524), .CP(clk), .Q(
        Sin3[2]) );
  FDS2L \Sin3_reg[1]  ( .CR(1'b1), .D(Sin2[1]), .LD(n524), .CP(clk), .Q(
        Sin3[1]) );
  FDS2L \Sin3_reg[0]  ( .CR(1'b1), .D(Sin2[0]), .LD(n524), .CP(clk), .Q(
        Sin3[0]) );
  FDS2L \Cos3_reg[15]  ( .CR(1'b1), .D(Cos2[15]), .LD(n524), .CP(clk), .Q(
        Cos3[15]) );
  FDS2L \Cos3_reg[14]  ( .CR(1'b1), .D(Cos2[14]), .LD(n523), .CP(clk), .Q(
        Cos3[14]) );
  FDS2L \Cos3_reg[13]  ( .CR(1'b1), .D(Cos2[13]), .LD(n523), .CP(clk), .Q(
        Cos3[13]) );
  FDS2L \Cos3_reg[12]  ( .CR(1'b1), .D(Cos2[12]), .LD(n523), .CP(clk), .Q(
        Cos3[12]) );
  FDS2L \Cos3_reg[11]  ( .CR(1'b1), .D(Cos2[11]), .LD(n523), .CP(clk), .Q(
        Cos3[11]) );
  FDS2L \Cos3_reg[10]  ( .CR(1'b1), .D(Cos2[10]), .LD(n523), .CP(clk), .Q(
        Cos3[10]) );
  FDS2L \Cos3_reg[9]  ( .CR(1'b1), .D(Cos2[9]), .LD(n523), .CP(clk), .Q(
        Cos3[9]) );
  FDS2L \Cos3_reg[8]  ( .CR(1'b1), .D(Cos2[8]), .LD(n523), .CP(clk), .Q(
        Cos3[8]) );
  FDS2L \Cos3_reg[7]  ( .CR(1'b1), .D(Cos2[7]), .LD(n523), .CP(clk), .Q(
        Cos3[7]) );
  FDS2L \Cos3_reg[6]  ( .CR(1'b1), .D(Cos2[6]), .LD(n523), .CP(clk), .Q(
        Cos3[6]) );
  FDS2L \Cos3_reg[5]  ( .CR(1'b1), .D(Cos2[5]), .LD(n523), .CP(clk), .Q(
        Cos3[5]) );
  FDS2L \Cos3_reg[4]  ( .CR(1'b1), .D(Cos2[4]), .LD(n523), .CP(clk), .Q(
        Cos3[4]) );
  FDS2L \Cos3_reg[3]  ( .CR(1'b1), .D(Cos2[3]), .LD(n523), .CP(clk), .Q(
        Cos3[3]) );
  FDS2L \Cos3_reg[2]  ( .CR(1'b1), .D(Cos2[2]), .LD(n522), .CP(clk), .Q(
        Cos3[2]) );
  FDS2L \Cos3_reg[1]  ( .CR(1'b1), .D(Cos2[1]), .LD(n522), .CP(clk), .Q(
        Cos3[1]) );
  FDS2L \Cos3_reg[0]  ( .CR(1'b1), .D(Cos2[0]), .LD(n522), .CP(clk), .Q(
        Cos3[0]) );
  FDS2L \Sin4_reg[15]  ( .CR(1'b1), .D(Sin3[15]), .LD(n522), .CP(clk), .Q(
        Sin4[15]) );
  FDS2L \Sin4_reg[14]  ( .CR(1'b1), .D(Sin3[14]), .LD(n522), .CP(clk), .Q(
        Sin4[14]) );
  FDS2L \Sin4_reg[13]  ( .CR(1'b1), .D(Sin3[13]), .LD(n522), .CP(clk), .Q(
        Sin4[13]) );
  FDS2L \Sin4_reg[12]  ( .CR(1'b1), .D(Sin3[12]), .LD(n522), .CP(clk), .Q(
        Sin4[12]) );
  FDS2L \Sin4_reg[11]  ( .CR(1'b1), .D(Sin3[11]), .LD(n522), .CP(clk), .Q(
        Sin4[11]) );
  FDS2L \Sin4_reg[10]  ( .CR(1'b1), .D(Sin3[10]), .LD(n522), .CP(clk), .Q(
        Sin4[10]) );
  FDS2L \Sin4_reg[9]  ( .CR(1'b1), .D(Sin3[9]), .LD(n522), .CP(clk), .Q(
        Sin4[9]) );
  FDS2L \Sin4_reg[8]  ( .CR(1'b1), .D(Sin3[8]), .LD(n522), .CP(clk), .Q(
        Sin4[8]) );
  FDS2L \Sin4_reg[7]  ( .CR(1'b1), .D(Sin3[7]), .LD(n522), .CP(clk), .Q(
        Sin4[7]) );
  FDS2L \Sin4_reg[6]  ( .CR(1'b1), .D(Sin3[6]), .LD(n521), .CP(clk), .Q(
        Sin4[6]) );
  FDS2L \Sin4_reg[5]  ( .CR(1'b1), .D(Sin3[5]), .LD(n521), .CP(clk), .Q(
        Sin4[5]) );
  FDS2L \Sin4_reg[4]  ( .CR(1'b1), .D(Sin3[4]), .LD(n521), .CP(clk), .Q(
        Sin4[4]) );
  FDS2L \Sin4_reg[3]  ( .CR(1'b1), .D(Sin3[3]), .LD(n521), .CP(clk), .Q(
        Sin4[3]) );
  FDS2L \Sin4_reg[2]  ( .CR(1'b1), .D(Sin3[2]), .LD(n521), .CP(clk), .Q(
        Sin4[2]) );
  FDS2L \Sin4_reg[1]  ( .CR(1'b1), .D(Sin3[1]), .LD(n521), .CP(clk), .Q(
        Sin4[1]) );
  FDS2L \Sin4_reg[0]  ( .CR(1'b1), .D(Sin3[0]), .LD(n521), .CP(clk), .Q(
        Sin4[0]) );
  FDS2L \Cos4_reg[15]  ( .CR(1'b1), .D(Cos3[15]), .LD(n521), .CP(clk), .Q(
        Cos4[15]) );
  FDS2L \Cos4_reg[14]  ( .CR(1'b1), .D(Cos3[14]), .LD(n521), .CP(clk), .Q(
        Cos4[14]) );
  FDS2L \Cos4_reg[13]  ( .CR(1'b1), .D(Cos3[13]), .LD(n521), .CP(clk), .Q(
        Cos4[13]) );
  FDS2L \Cos4_reg[12]  ( .CR(1'b1), .D(Cos3[12]), .LD(n521), .CP(clk), .Q(
        Cos4[12]) );
  FDS2L \Cos4_reg[11]  ( .CR(1'b1), .D(Cos3[11]), .LD(n521), .CP(clk), .Q(
        Cos4[11]) );
  FDS2L \Cos4_reg[10]  ( .CR(1'b1), .D(Cos3[10]), .LD(n520), .CP(clk), .Q(
        Cos4[10]) );
  FDS2L \Cos4_reg[9]  ( .CR(1'b1), .D(Cos3[9]), .LD(n520), .CP(clk), .Q(
        Cos4[9]) );
  FDS2L \Cos4_reg[8]  ( .CR(1'b1), .D(Cos3[8]), .LD(n520), .CP(clk), .Q(
        Cos4[8]) );
  FDS2L \Cos4_reg[7]  ( .CR(1'b1), .D(Cos3[7]), .LD(n520), .CP(clk), .Q(
        Cos4[7]) );
  FDS2L \Cos4_reg[6]  ( .CR(1'b1), .D(Cos3[6]), .LD(n520), .CP(clk), .Q(
        Cos4[6]) );
  FDS2L \Cos4_reg[5]  ( .CR(1'b1), .D(Cos3[5]), .LD(n520), .CP(clk), .Q(
        Cos4[5]) );
  FDS2L \Cos4_reg[4]  ( .CR(1'b1), .D(Cos3[4]), .LD(n520), .CP(clk), .Q(
        Cos4[4]) );
  FDS2L \Cos4_reg[3]  ( .CR(1'b1), .D(Cos3[3]), .LD(n520), .CP(clk), .Q(
        Cos4[3]) );
  FDS2L \Cos4_reg[2]  ( .CR(1'b1), .D(Cos3[2]), .LD(n520), .CP(clk), .Q(
        Cos4[2]) );
  FDS2L \Cos4_reg[1]  ( .CR(1'b1), .D(Cos3[1]), .LD(n520), .CP(clk), .Q(
        Cos4[1]) );
  FDS2L \Cos4_reg[0]  ( .CR(1'b1), .D(Cos3[0]), .LD(n520), .CP(clk), .Q(
        Cos4[0]) );
  FDS2L \Sin5_reg[15]  ( .CR(1'b1), .D(Sin4[15]), .LD(n520), .CP(clk), .Q(
        Sin5[15]) );
  FDS2L \Sin5_reg[14]  ( .CR(1'b1), .D(Sin4[14]), .LD(n519), .CP(clk), .Q(
        Sin5[14]) );
  FDS2L \Sin5_reg[13]  ( .CR(1'b1), .D(Sin4[13]), .LD(n519), .CP(clk), .Q(
        Sin5[13]) );
  FDS2L \Sin5_reg[12]  ( .CR(1'b1), .D(Sin4[12]), .LD(n519), .CP(clk), .Q(
        Sin5[12]) );
  FDS2L \Sin5_reg[11]  ( .CR(1'b1), .D(Sin4[11]), .LD(n519), .CP(clk), .Q(
        Sin5[11]) );
  FDS2L \Sin5_reg[10]  ( .CR(1'b1), .D(Sin4[10]), .LD(n519), .CP(clk), .Q(
        Sin5[10]) );
  FDS2L \Sin5_reg[9]  ( .CR(1'b1), .D(Sin4[9]), .LD(n519), .CP(clk), .Q(
        Sin5[9]) );
  FDS2L \Sin5_reg[8]  ( .CR(1'b1), .D(Sin4[8]), .LD(n519), .CP(clk), .Q(
        Sin5[8]) );
  FDS2L \Sin5_reg[7]  ( .CR(1'b1), .D(Sin4[7]), .LD(n519), .CP(clk), .Q(
        Sin5[7]) );
  FDS2L \Sin5_reg[6]  ( .CR(1'b1), .D(Sin4[6]), .LD(n519), .CP(clk), .Q(
        Sin5[6]) );
  FDS2L \Sin5_reg[5]  ( .CR(1'b1), .D(Sin4[5]), .LD(n519), .CP(clk), .Q(
        Sin5[5]) );
  FDS2L \Sin5_reg[4]  ( .CR(1'b1), .D(Sin4[4]), .LD(n519), .CP(clk), .Q(
        Sin5[4]) );
  FDS2L \Sin5_reg[3]  ( .CR(1'b1), .D(Sin4[3]), .LD(n519), .CP(clk), .Q(
        Sin5[3]) );
  FDS2L \Sin5_reg[2]  ( .CR(1'b1), .D(Sin4[2]), .LD(n518), .CP(clk), .Q(
        Sin5[2]) );
  FDS2L \Sin5_reg[1]  ( .CR(1'b1), .D(Sin4[1]), .LD(n518), .CP(clk), .Q(
        Sin5[1]) );
  FDS2L \Sin5_reg[0]  ( .CR(1'b1), .D(Sin4[0]), .LD(n518), .CP(clk), .Q(
        Sin5[0]) );
  FDS2L \Cos5_reg[15]  ( .CR(1'b1), .D(Cos4[15]), .LD(n518), .CP(clk), .Q(
        Cos5[15]) );
  FDS2L \Cos5_reg[14]  ( .CR(1'b1), .D(Cos4[14]), .LD(n518), .CP(clk), .Q(
        Cos5[14]) );
  FDS2L \Cos5_reg[13]  ( .CR(1'b1), .D(Cos4[13]), .LD(n518), .CP(clk), .Q(
        Cos5[13]) );
  FDS2L \Cos5_reg[12]  ( .CR(1'b1), .D(Cos4[12]), .LD(n518), .CP(clk), .Q(
        Cos5[12]) );
  FDS2L \Cos5_reg[11]  ( .CR(1'b1), .D(Cos4[11]), .LD(n518), .CP(clk), .Q(
        Cos5[11]) );
  FDS2L \Cos5_reg[10]  ( .CR(1'b1), .D(Cos4[10]), .LD(n518), .CP(clk), .Q(
        Cos5[10]) );
  FDS2L \Cos5_reg[9]  ( .CR(1'b1), .D(Cos4[9]), .LD(n518), .CP(clk), .Q(
        Cos5[9]) );
  FDS2L \Cos5_reg[8]  ( .CR(1'b1), .D(Cos4[8]), .LD(n518), .CP(clk), .Q(
        Cos5[8]) );
  FDS2L \Cos5_reg[7]  ( .CR(1'b1), .D(Cos4[7]), .LD(n518), .CP(clk), .Q(
        Cos5[7]) );
  FDS2L \Cos5_reg[6]  ( .CR(1'b1), .D(Cos4[6]), .LD(n517), .CP(clk), .Q(
        Cos5[6]) );
  FDS2L \Cos5_reg[5]  ( .CR(1'b1), .D(Cos4[5]), .LD(n517), .CP(clk), .Q(
        Cos5[5]) );
  FDS2L \Cos5_reg[4]  ( .CR(1'b1), .D(Cos4[4]), .LD(n517), .CP(clk), .Q(
        Cos5[4]) );
  FDS2L \Cos5_reg[3]  ( .CR(1'b1), .D(Cos4[3]), .LD(n517), .CP(clk), .Q(
        Cos5[3]) );
  FDS2L \Cos5_reg[2]  ( .CR(1'b1), .D(Cos4[2]), .LD(n517), .CP(clk), .Q(
        Cos5[2]) );
  FDS2L \Cos5_reg[1]  ( .CR(1'b1), .D(Cos4[1]), .LD(n517), .CP(clk), .Q(
        Cos5[1]) );
  FDS2L \Cos5_reg[0]  ( .CR(1'b1), .D(Cos4[0]), .LD(n517), .CP(clk), .Q(
        Cos5[0]) );
  FDS2L \Sin6_reg[15]  ( .CR(1'b1), .D(Sin5[15]), .LD(n517), .CP(clk), .Q(
        Sin6[15]) );
  FDS2L \Sin6_reg[14]  ( .CR(1'b1), .D(Sin5[14]), .LD(n517), .CP(clk), .Q(
        Sin6[14]) );
  FDS2L \Sin6_reg[13]  ( .CR(1'b1), .D(Sin5[13]), .LD(n517), .CP(clk), .Q(
        Sin6[13]) );
  FDS2L \Sin6_reg[12]  ( .CR(1'b1), .D(Sin5[12]), .LD(n517), .CP(clk), .Q(
        Sin6[12]) );
  FDS2L \Sin6_reg[11]  ( .CR(1'b1), .D(Sin5[11]), .LD(n517), .CP(clk), .Q(
        Sin6[11]) );
  FDS2L \Sin6_reg[10]  ( .CR(1'b1), .D(Sin5[10]), .LD(n516), .CP(clk), .Q(
        Sin6[10]) );
  FDS2L \Sin6_reg[9]  ( .CR(1'b1), .D(Sin5[9]), .LD(n516), .CP(clk), .Q(
        Sin6[9]) );
  FDS2L \Sin6_reg[8]  ( .CR(1'b1), .D(Sin5[8]), .LD(n516), .CP(clk), .Q(
        Sin6[8]) );
  FDS2L \Sin6_reg[7]  ( .CR(1'b1), .D(Sin5[7]), .LD(n516), .CP(clk), .Q(
        Sin6[7]) );
  FDS2L \Sin6_reg[6]  ( .CR(1'b1), .D(Sin5[6]), .LD(n516), .CP(clk), .Q(
        Sin6[6]) );
  FDS2L \Sin6_reg[5]  ( .CR(1'b1), .D(Sin5[5]), .LD(n516), .CP(clk), .Q(
        Sin6[5]) );
  FDS2L \Sin6_reg[4]  ( .CR(1'b1), .D(Sin5[4]), .LD(n516), .CP(clk), .Q(
        Sin6[4]) );
  FDS2L \Sin6_reg[3]  ( .CR(1'b1), .D(Sin5[3]), .LD(n516), .CP(clk), .Q(
        Sin6[3]) );
  FDS2L \Sin6_reg[2]  ( .CR(1'b1), .D(Sin5[2]), .LD(n516), .CP(clk), .Q(
        Sin6[2]) );
  FDS2L \Sin6_reg[1]  ( .CR(1'b1), .D(Sin5[1]), .LD(n516), .CP(clk), .Q(
        Sin6[1]) );
  FDS2L \Sin6_reg[0]  ( .CR(1'b1), .D(Sin5[0]), .LD(n516), .CP(clk), .Q(
        Sin6[0]) );
  FDS2L \Cos6_reg[15]  ( .CR(1'b1), .D(Cos5[15]), .LD(n516), .CP(clk), .Q(
        Cos6[15]) );
  FDS2L \Cos6_reg[14]  ( .CR(1'b1), .D(Cos5[14]), .LD(n515), .CP(clk), .Q(
        Cos6[14]) );
  FDS2L \Cos6_reg[13]  ( .CR(1'b1), .D(Cos5[13]), .LD(n515), .CP(clk), .Q(
        Cos6[13]) );
  FDS2L \Cos6_reg[12]  ( .CR(1'b1), .D(Cos5[12]), .LD(n515), .CP(clk), .Q(
        Cos6[12]) );
  FDS2L \Cos6_reg[11]  ( .CR(1'b1), .D(Cos5[11]), .LD(n515), .CP(clk), .Q(
        Cos6[11]) );
  FDS2L \Cos6_reg[10]  ( .CR(1'b1), .D(Cos5[10]), .LD(n515), .CP(clk), .Q(
        Cos6[10]) );
  FDS2L \Cos6_reg[9]  ( .CR(1'b1), .D(Cos5[9]), .LD(n515), .CP(clk), .Q(
        Cos6[9]) );
  FDS2L \Cos6_reg[8]  ( .CR(1'b1), .D(Cos5[8]), .LD(n515), .CP(clk), .Q(
        Cos6[8]) );
  FDS2L \Cos6_reg[7]  ( .CR(1'b1), .D(Cos5[7]), .LD(n515), .CP(clk), .Q(
        Cos6[7]) );
  FDS2L \Cos6_reg[6]  ( .CR(1'b1), .D(Cos5[6]), .LD(n515), .CP(clk), .Q(
        Cos6[6]) );
  FDS2L \Cos6_reg[5]  ( .CR(1'b1), .D(Cos5[5]), .LD(n515), .CP(clk), .Q(
        Cos6[5]) );
  FDS2L \Cos6_reg[4]  ( .CR(1'b1), .D(Cos5[4]), .LD(n515), .CP(clk), .Q(
        Cos6[4]) );
  FDS2L \Cos6_reg[3]  ( .CR(1'b1), .D(Cos5[3]), .LD(n515), .CP(clk), .Q(
        Cos6[3]) );
  FDS2L \Cos6_reg[2]  ( .CR(1'b1), .D(Cos5[2]), .LD(n514), .CP(clk), .Q(
        Cos6[2]) );
  FDS2L \Cos6_reg[1]  ( .CR(1'b1), .D(Cos5[1]), .LD(n514), .CP(clk), .Q(
        Cos6[1]) );
  FDS2L \Cos6_reg[0]  ( .CR(1'b1), .D(Cos5[0]), .LD(n514), .CP(clk), .Q(
        Cos6[0]) );
  FDS2L \Sin7_reg[15]  ( .CR(1'b1), .D(Sin6[15]), .LD(n514), .CP(clk), .Q(
        Sin7[15]) );
  FDS2L \Sin7_reg[14]  ( .CR(1'b1), .D(Sin6[14]), .LD(n514), .CP(clk), .Q(
        Sin7[14]) );
  FDS2L \Sin7_reg[13]  ( .CR(1'b1), .D(Sin6[13]), .LD(n514), .CP(clk), .Q(
        Sin7[13]) );
  FDS2L \Sin7_reg[12]  ( .CR(1'b1), .D(Sin6[12]), .LD(n514), .CP(clk), .Q(
        Sin7[12]) );
  FDS2L \Sin7_reg[11]  ( .CR(1'b1), .D(Sin6[11]), .LD(n514), .CP(clk), .Q(
        Sin7[11]) );
  FDS2L \Sin7_reg[10]  ( .CR(1'b1), .D(Sin6[10]), .LD(n514), .CP(clk), .Q(
        Sin7[10]) );
  FDS2L \Sin7_reg[9]  ( .CR(1'b1), .D(Sin6[9]), .LD(n514), .CP(clk), .Q(
        Sin7[9]) );
  FDS2L \Sin7_reg[8]  ( .CR(1'b1), .D(Sin6[8]), .LD(n514), .CP(clk), .Q(
        Sin7[8]) );
  FDS2L \Sin7_reg[7]  ( .CR(1'b1), .D(Sin6[7]), .LD(n514), .CP(clk), .Q(
        Sin7[7]) );
  FDS2L \Sin7_reg[6]  ( .CR(1'b1), .D(Sin6[6]), .LD(n513), .CP(clk), .Q(
        Sin7[6]) );
  FDS2L \Sin7_reg[5]  ( .CR(1'b1), .D(Sin6[5]), .LD(n513), .CP(clk), .Q(
        Sin7[5]) );
  FDS2L \Sin7_reg[4]  ( .CR(1'b1), .D(Sin6[4]), .LD(n513), .CP(clk), .Q(
        Sin7[4]) );
  FDS2L \Sin7_reg[3]  ( .CR(1'b1), .D(Sin6[3]), .LD(n513), .CP(clk), .Q(
        Sin7[3]) );
  FDS2L \Sin7_reg[2]  ( .CR(1'b1), .D(Sin6[2]), .LD(n513), .CP(clk), .Q(
        Sin7[2]) );
  FDS2L \Sin7_reg[1]  ( .CR(1'b1), .D(Sin6[1]), .LD(n513), .CP(clk), .Q(
        Sin7[1]) );
  FDS2L \Sin7_reg[0]  ( .CR(1'b1), .D(Sin6[0]), .LD(n513), .CP(clk), .Q(
        Sin7[0]) );
  FDS2L \Cos7_reg[15]  ( .CR(1'b1), .D(Cos6[15]), .LD(n513), .CP(clk), .Q(
        Cos7[15]) );
  FDS2L \Cos7_reg[14]  ( .CR(1'b1), .D(Cos6[14]), .LD(n513), .CP(clk), .Q(
        Cos7[14]) );
  FDS2L \Cos7_reg[13]  ( .CR(1'b1), .D(Cos6[13]), .LD(n513), .CP(clk), .Q(
        Cos7[13]) );
  FDS2L \Cos7_reg[12]  ( .CR(1'b1), .D(Cos6[12]), .LD(n513), .CP(clk), .Q(
        Cos7[12]) );
  FDS2L \Cos7_reg[11]  ( .CR(1'b1), .D(Cos6[11]), .LD(n513), .CP(clk), .Q(
        Cos7[11]) );
  FDS2L \Cos7_reg[10]  ( .CR(1'b1), .D(Cos6[10]), .LD(n512), .CP(clk), .Q(
        Cos7[10]) );
  FDS2L \Cos7_reg[9]  ( .CR(1'b1), .D(Cos6[9]), .LD(n512), .CP(clk), .Q(
        Cos7[9]) );
  FDS2L \Cos7_reg[8]  ( .CR(1'b1), .D(Cos6[8]), .LD(n512), .CP(clk), .Q(
        Cos7[8]) );
  FDS2L \Cos7_reg[7]  ( .CR(1'b1), .D(Cos6[7]), .LD(n512), .CP(clk), .Q(
        Cos7[7]) );
  FDS2L \Cos7_reg[6]  ( .CR(1'b1), .D(Cos6[6]), .LD(n512), .CP(clk), .Q(
        Cos7[6]) );
  FDS2L \Cos7_reg[5]  ( .CR(1'b1), .D(Cos6[5]), .LD(n512), .CP(clk), .Q(
        Cos7[5]) );
  FDS2L \Cos7_reg[4]  ( .CR(1'b1), .D(Cos6[4]), .LD(n512), .CP(clk), .Q(
        Cos7[4]) );
  FDS2L \Cos7_reg[3]  ( .CR(1'b1), .D(Cos6[3]), .LD(n512), .CP(clk), .Q(
        Cos7[3]) );
  FDS2L \Cos7_reg[2]  ( .CR(1'b1), .D(Cos6[2]), .LD(n512), .CP(clk), .Q(
        Cos7[2]) );
  FDS2L \Cos7_reg[1]  ( .CR(1'b1), .D(Cos6[1]), .LD(n512), .CP(clk), .Q(
        Cos7[1]) );
  FDS2L \Cos7_reg[0]  ( .CR(1'b1), .D(Cos6[0]), .LD(n512), .CP(clk), .Q(
        Cos7[0]) );
  FDS2L \Sin8_reg[15]  ( .CR(1'b1), .D(Sin7[15]), .LD(n512), .CP(clk), .Q(
        Sin8[15]) );
  FDS2L \Sin8_reg[14]  ( .CR(1'b1), .D(Sin7[14]), .LD(n511), .CP(clk), .Q(
        Sin8[14]) );
  FDS2L \Sin8_reg[13]  ( .CR(1'b1), .D(Sin7[13]), .LD(n511), .CP(clk), .Q(
        Sin8[13]) );
  FDS2L \Sin8_reg[12]  ( .CR(1'b1), .D(Sin7[12]), .LD(n511), .CP(clk), .Q(
        Sin8[12]) );
  FDS2L \Sin8_reg[11]  ( .CR(1'b1), .D(Sin7[11]), .LD(n511), .CP(clk), .Q(
        Sin8[11]) );
  FDS2L \Sin8_reg[10]  ( .CR(1'b1), .D(Sin7[10]), .LD(n511), .CP(clk), .Q(
        Sin8[10]) );
  FDS2L \Sin8_reg[9]  ( .CR(1'b1), .D(Sin7[9]), .LD(n511), .CP(clk), .Q(
        Sin8[9]) );
  FDS2L \Sin8_reg[8]  ( .CR(1'b1), .D(Sin7[8]), .LD(n511), .CP(clk), .Q(
        Sin8[8]) );
  FDS2L \Sin8_reg[7]  ( .CR(1'b1), .D(Sin7[7]), .LD(n511), .CP(clk), .Q(
        Sin8[7]) );
  FDS2L \Sin8_reg[6]  ( .CR(1'b1), .D(Sin7[6]), .LD(n511), .CP(clk), .Q(
        Sin8[6]) );
  FDS2L \Sin8_reg[5]  ( .CR(1'b1), .D(Sin7[5]), .LD(n511), .CP(clk), .Q(
        Sin8[5]) );
  FDS2L \Sin8_reg[4]  ( .CR(1'b1), .D(Sin7[4]), .LD(n511), .CP(clk), .Q(
        Sin8[4]) );
  FDS2L \Sin8_reg[3]  ( .CR(1'b1), .D(Sin7[3]), .LD(n511), .CP(clk), .Q(
        Sin8[3]) );
  FDS2L \Sin8_reg[2]  ( .CR(1'b1), .D(Sin7[2]), .LD(n510), .CP(clk), .Q(
        Sin8[2]) );
  FDS2L \Sin8_reg[1]  ( .CR(1'b1), .D(Sin7[1]), .LD(n510), .CP(clk), .Q(
        Sin8[1]) );
  FDS2L \Sin8_reg[0]  ( .CR(1'b1), .D(Sin7[0]), .LD(n510), .CP(clk), .Q(
        Sin8[0]) );
  FDS2L \Cos8_reg[15]  ( .CR(1'b1), .D(Cos7[15]), .LD(n510), .CP(clk), .Q(
        Cos8[15]) );
  FDS2L \Cos8_reg[14]  ( .CR(1'b1), .D(Cos7[14]), .LD(n510), .CP(clk), .Q(
        Cos8[14]) );
  FDS2L \Cos8_reg[13]  ( .CR(1'b1), .D(Cos7[13]), .LD(n510), .CP(clk), .Q(
        Cos8[13]) );
  FDS2L \Cos8_reg[12]  ( .CR(1'b1), .D(Cos7[12]), .LD(n510), .CP(clk), .Q(
        Cos8[12]) );
  FDS2L \Cos8_reg[11]  ( .CR(1'b1), .D(Cos7[11]), .LD(n510), .CP(clk), .Q(
        Cos8[11]) );
  FDS2L \Cos8_reg[10]  ( .CR(1'b1), .D(Cos7[10]), .LD(n510), .CP(clk), .Q(
        Cos8[10]) );
  FDS2L \Cos8_reg[9]  ( .CR(1'b1), .D(Cos7[9]), .LD(n510), .CP(clk), .Q(
        Cos8[9]) );
  FDS2L \Cos8_reg[8]  ( .CR(1'b1), .D(Cos7[8]), .LD(n510), .CP(clk), .Q(
        Cos8[8]) );
  FDS2L \Cos8_reg[7]  ( .CR(1'b1), .D(Cos7[7]), .LD(n510), .CP(clk), .Q(
        Cos8[7]) );
  FDS2L \Cos8_reg[6]  ( .CR(1'b1), .D(Cos7[6]), .LD(n509), .CP(clk), .Q(
        Cos8[6]) );
  FDS2L \Cos8_reg[5]  ( .CR(1'b1), .D(Cos7[5]), .LD(n509), .CP(clk), .Q(
        Cos8[5]) );
  FDS2L \Cos8_reg[4]  ( .CR(1'b1), .D(Cos7[4]), .LD(n509), .CP(clk), .Q(
        Cos8[4]) );
  FDS2L \Cos8_reg[3]  ( .CR(1'b1), .D(Cos7[3]), .LD(n509), .CP(clk), .Q(
        Cos8[3]) );
  FDS2L \Cos8_reg[2]  ( .CR(1'b1), .D(Cos7[2]), .LD(n509), .CP(clk), .Q(
        Cos8[2]) );
  FDS2L \Cos8_reg[1]  ( .CR(1'b1), .D(Cos7[1]), .LD(n509), .CP(clk), .Q(
        Cos8[1]) );
  FDS2L \Cos8_reg[0]  ( .CR(1'b1), .D(Cos7[0]), .LD(n509), .CP(clk), .Q(
        Cos8[0]) );
  FDS2L \Sin1_reg[15]  ( .CR(1'b1), .D(Sin8[15]), .LD(n509), .CP(clk), .Q(
        Sin1[15]) );
  FDS2L \Sin1_reg[14]  ( .CR(1'b1), .D(Sin8[14]), .LD(n509), .CP(clk), .Q(
        Sin1[14]) );
  FDS2L \Sin1_reg[13]  ( .CR(1'b1), .D(Sin8[13]), .LD(n509), .CP(clk), .Q(
        Sin1[13]) );
  FDS2L \Sin1_reg[12]  ( .CR(1'b1), .D(Sin8[12]), .LD(n509), .CP(clk), .Q(
        Sin1[12]) );
  FDS2L \Sin1_reg[11]  ( .CR(1'b1), .D(Sin8[11]), .LD(n509), .CP(clk), .Q(
        Sin1[11]) );
  FDS2L \Sin1_reg[10]  ( .CR(1'b1), .D(Sin8[10]), .LD(n508), .CP(clk), .Q(
        Sin1[10]) );
  FDS2L \Sin1_reg[9]  ( .CR(1'b1), .D(Sin8[9]), .LD(n508), .CP(clk), .Q(
        Sin1[9]) );
  FDS2L \Sin1_reg[8]  ( .CR(1'b1), .D(Sin8[8]), .LD(n508), .CP(clk), .Q(
        Sin1[8]) );
  FDS2L \Sin1_reg[7]  ( .CR(1'b1), .D(Sin8[7]), .LD(n508), .CP(clk), .Q(
        Sin1[7]) );
  FDS2L \Sin1_reg[6]  ( .CR(1'b1), .D(Sin8[6]), .LD(n508), .CP(clk), .Q(
        Sin1[6]) );
  FDS2L \Sin1_reg[5]  ( .CR(1'b1), .D(Sin8[5]), .LD(n508), .CP(clk), .Q(
        Sin1[5]) );
  FDS2L \Sin1_reg[4]  ( .CR(1'b1), .D(Sin8[4]), .LD(n508), .CP(clk), .Q(
        Sin1[4]) );
  FDS2L \Sin1_reg[3]  ( .CR(1'b1), .D(Sin8[3]), .LD(n508), .CP(clk), .Q(
        Sin1[3]) );
  FDS2L \Sin1_reg[2]  ( .CR(1'b1), .D(Sin8[2]), .LD(n508), .CP(clk), .Q(
        Sin1[2]) );
  FDS2L \Sin1_reg[1]  ( .CR(1'b1), .D(Sin8[1]), .LD(n508), .CP(clk), .Q(
        Sin1[1]) );
  FDS2L \Sin1_reg[0]  ( .CR(1'b1), .D(Sin8[0]), .LD(n508), .CP(clk), .Q(
        Sin1[0]) );
  FDS2L \Cos1_reg[15]  ( .CR(1'b1), .D(Cos8[15]), .LD(n508), .CP(clk), .Q(
        Cos1[15]) );
  FDS2L \Cos1_reg[14]  ( .CR(1'b1), .D(Cos8[14]), .LD(n507), .CP(clk), .Q(
        Cos1[14]) );
  FDS2L \Cos1_reg[13]  ( .CR(1'b1), .D(Cos8[13]), .LD(n507), .CP(clk), .Q(
        Cos1[13]) );
  FDS2L \Cos1_reg[12]  ( .CR(1'b1), .D(Cos8[12]), .LD(n507), .CP(clk), .Q(
        Cos1[12]) );
  FDS2L \Cos1_reg[11]  ( .CR(1'b1), .D(Cos8[11]), .LD(n507), .CP(clk), .Q(
        Cos1[11]) );
  FDS2L \Cos1_reg[10]  ( .CR(1'b1), .D(Cos8[10]), .LD(n507), .CP(clk), .Q(
        Cos1[10]) );
  FDS2L \Cos1_reg[9]  ( .CR(1'b1), .D(Cos8[9]), .LD(n507), .CP(clk), .Q(
        Cos1[9]) );
  FDS2L \Cos1_reg[8]  ( .CR(1'b1), .D(Cos8[8]), .LD(n507), .CP(clk), .Q(
        Cos1[8]) );
  FDS2L \Cos1_reg[7]  ( .CR(1'b1), .D(Cos8[7]), .LD(n507), .CP(clk), .Q(
        Cos1[7]) );
  FDS2L \Cos1_reg[6]  ( .CR(1'b1), .D(Cos8[6]), .LD(n507), .CP(clk), .Q(
        Cos1[6]) );
  FDS2L \Cos1_reg[5]  ( .CR(1'b1), .D(Cos8[5]), .LD(n507), .CP(clk), .Q(
        Cos1[5]) );
  FDS2L \Cos1_reg[4]  ( .CR(1'b1), .D(Cos8[4]), .LD(n507), .CP(clk), .Q(
        Cos1[4]) );
  FDS2L \Cos1_reg[3]  ( .CR(1'b1), .D(Cos8[3]), .LD(n507), .CP(clk), .Q(
        Cos1[3]) );
  FDS2L \Cos1_reg[2]  ( .CR(1'b1), .D(Cos8[2]), .LD(n506), .CP(clk), .Q(
        Cos1[2]) );
  FDS2L \Cos1_reg[1]  ( .CR(1'b1), .D(Cos8[1]), .LD(n506), .CP(clk), .Q(
        Cos1[1]) );
  FDS2L \Cos1_reg[0]  ( .CR(1'b1), .D(Cos8[0]), .LD(n506), .CP(clk), .Q(
        Cos1[0]) );
  FDS2L \Sin_reg[15]  ( .CR(1'b1), .D(Sin1[15]), .LD(n506), .CP(clk), .Q(
        Sin[15]) );
  FDS2L \Cos_reg[15]  ( .CR(1'b1), .D(Cos1[15]), .LD(n505), .CP(clk), .Q(
        Cos[15]) );
  FDS2L \X0_reg[15]  ( .CR(1'b1), .D(Sin[15]), .LD(n501), .CP(clk), .Q(X0[15])
         );
  FDS2L \X1_reg[15]  ( .CR(1'b1), .D(Cos[15]), .LD(n501), .CP(clk), .Q(X1[15])
         );
  FDS2L \RegX0_reg[31]  ( .CR(1'b1), .D(N19), .LD(n501), .CP(clk), .Q(
        RegX0[31]) );
  FDS2L \X0_reg[14]  ( .CR(1'b1), .D(RegX0[31]), .LD(n501), .CP(clk), .Q(
        X0[14]) );
  FDS2L \RegX0_reg[30]  ( .CR(1'b1), .D(N18), .LD(n501), .CP(clk), .Q(
        RegX0[30]) );
  FDS2L \X0_reg[13]  ( .CR(1'b1), .D(RegX0[30]), .LD(n501), .CP(clk), .Q(
        X0[13]) );
  FDS2L \RegX0_reg[29]  ( .CR(1'b1), .D(N17), .LD(n500), .CP(clk), .Q(
        RegX0[29]) );
  FDS2L \X0_reg[12]  ( .CR(1'b1), .D(RegX0[29]), .LD(n500), .CP(clk), .Q(
        X0[12]) );
  FDS2L \RegX0_reg[28]  ( .CR(1'b1), .D(N16), .LD(n500), .CP(clk), .Q(
        RegX0[28]) );
  FDS2L \X0_reg[11]  ( .CR(1'b1), .D(RegX0[28]), .LD(n500), .CP(clk), .Q(
        X0[11]) );
  FDS2L \RegX0_reg[27]  ( .CR(1'b1), .D(N15), .LD(n500), .CP(clk), .Q(
        RegX0[27]) );
  FDS2L \X0_reg[10]  ( .CR(1'b1), .D(RegX0[27]), .LD(n500), .CP(clk), .Q(
        X0[10]) );
  FDS2L \RegX0_reg[26]  ( .CR(1'b1), .D(N14), .LD(n500), .CP(clk), .Q(
        RegX0[26]) );
  FDS2L \X0_reg[9]  ( .CR(1'b1), .D(RegX0[26]), .LD(n500), .CP(clk), .Q(X0[9])
         );
  FDS2L \RegX0_reg[25]  ( .CR(1'b1), .D(N13), .LD(n500), .CP(clk), .Q(
        RegX0[25]) );
  FDS2L \X0_reg[8]  ( .CR(1'b1), .D(RegX0[25]), .LD(n500), .CP(clk), .Q(X0[8])
         );
  FDS2L \RegX0_reg[24]  ( .CR(1'b1), .D(N12), .LD(n500), .CP(clk), .Q(
        RegX0[24]) );
  FDS2L \X0_reg[7]  ( .CR(1'b1), .D(RegX0[24]), .LD(n500), .CP(clk), .Q(X0[7])
         );
  FDS2L \RegX0_reg[23]  ( .CR(1'b1), .D(N11), .LD(n499), .CP(clk), .Q(
        RegX0[23]) );
  FDS2L \X0_reg[6]  ( .CR(1'b1), .D(RegX0[23]), .LD(n499), .CP(clk), .Q(X0[6])
         );
  FDS2L \RegX0_reg[22]  ( .CR(1'b1), .D(N10), .LD(n499), .CP(clk), .Q(
        RegX0[22]) );
  FDS2L \X0_reg[5]  ( .CR(1'b1), .D(RegX0[22]), .LD(n499), .CP(clk), .Q(X0[5])
         );
  FDS2L \RegX0_reg[21]  ( .CR(1'b1), .D(N9), .LD(n499), .CP(clk), .Q(RegX0[21]) );
  FDS2L \X0_reg[4]  ( .CR(1'b1), .D(RegX0[21]), .LD(n499), .CP(clk), .Q(X0[4])
         );
  FDS2L \RegX0_reg[20]  ( .CR(1'b1), .D(N8), .LD(n499), .CP(clk), .Q(RegX0[20]) );
  FDS2L \X0_reg[3]  ( .CR(1'b1), .D(RegX0[20]), .LD(n499), .CP(clk), .Q(X0[3])
         );
  FDS2L \RegX0_reg[19]  ( .CR(1'b1), .D(N7), .LD(n499), .CP(clk), .Q(RegX0[19]) );
  FDS2L \X0_reg[2]  ( .CR(1'b1), .D(RegX0[19]), .LD(n499), .CP(clk), .Q(X0[2])
         );
  FDS2L \RegX0_reg[18]  ( .CR(1'b1), .D(N6), .LD(n499), .CP(clk), .Q(RegX0[18]) );
  FDS2L \X0_reg[1]  ( .CR(1'b1), .D(RegX0[18]), .LD(n499), .CP(clk), .Q(X0[1])
         );
  FDS2L \RegX0_reg[17]  ( .CR(1'b1), .D(N5), .LD(n498), .CP(clk), .Q(RegX0[17]) );
  FDS2L \X0_reg[0]  ( .CR(1'b1), .D(RegX0[17]), .LD(n498), .CP(clk), .Q(X0[0])
         );
  FDS2L \RegX1_reg[31]  ( .CR(1'b1), .D(N34), .LD(n498), .CP(clk), .Q(
        RegX1[31]) );
  FDS2L \X1_reg[14]  ( .CR(1'b1), .D(RegX1[31]), .LD(n498), .CP(clk), .Q(
        X1[14]) );
  FDS2L \RegX1_reg[30]  ( .CR(1'b1), .D(N33), .LD(n498), .CP(clk), .Q(
        RegX1[30]) );
  FDS2L \X1_reg[13]  ( .CR(1'b1), .D(RegX1[30]), .LD(n498), .CP(clk), .Q(
        X1[13]) );
  FDS2L \RegX1_reg[29]  ( .CR(1'b1), .D(N32), .LD(n498), .CP(clk), .Q(
        RegX1[29]) );
  FDS2L \X1_reg[12]  ( .CR(1'b1), .D(RegX1[29]), .LD(n498), .CP(clk), .Q(
        X1[12]) );
  FDS2L \RegX1_reg[28]  ( .CR(1'b1), .D(N31), .LD(n498), .CP(clk), .Q(
        RegX1[28]) );
  FDS2L \X1_reg[11]  ( .CR(1'b1), .D(RegX1[28]), .LD(n498), .CP(clk), .Q(
        X1[11]) );
  FDS2L \RegX1_reg[27]  ( .CR(1'b1), .D(N30), .LD(n498), .CP(clk), .Q(
        RegX1[27]) );
  FDS2L \X1_reg[10]  ( .CR(1'b1), .D(RegX1[27]), .LD(n498), .CP(clk), .Q(
        X1[10]) );
  FDS2L \RegX1_reg[26]  ( .CR(1'b1), .D(N29), .LD(n497), .CP(clk), .Q(
        RegX1[26]) );
  FDS2L \X1_reg[9]  ( .CR(1'b1), .D(RegX1[26]), .LD(n497), .CP(clk), .Q(X1[9])
         );
  FDS2L \RegX1_reg[25]  ( .CR(1'b1), .D(N28), .LD(n497), .CP(clk), .Q(
        RegX1[25]) );
  FDS2L \X1_reg[8]  ( .CR(1'b1), .D(RegX1[25]), .LD(n497), .CP(clk), .Q(X1[8])
         );
  FDS2L \RegX1_reg[24]  ( .CR(1'b1), .D(N27), .LD(n497), .CP(clk), .Q(
        RegX1[24]) );
  FDS2L \X1_reg[7]  ( .CR(1'b1), .D(RegX1[24]), .LD(n497), .CP(clk), .Q(X1[7])
         );
  FDS2L \RegX1_reg[23]  ( .CR(1'b1), .D(N26), .LD(n497), .CP(clk), .Q(
        RegX1[23]) );
  FDS2L \X1_reg[6]  ( .CR(1'b1), .D(RegX1[23]), .LD(n497), .CP(clk), .Q(X1[6])
         );
  FDS2L \RegX1_reg[22]  ( .CR(1'b1), .D(N25), .LD(n497), .CP(clk), .Q(
        RegX1[22]) );
  FDS2L \X1_reg[5]  ( .CR(1'b1), .D(RegX1[22]), .LD(n497), .CP(clk), .Q(X1[5])
         );
  FDS2L \RegX1_reg[21]  ( .CR(1'b1), .D(N24), .LD(n497), .CP(clk), .Q(
        RegX1[21]) );
  FDS2L \X1_reg[4]  ( .CR(1'b1), .D(RegX1[21]), .LD(n497), .CP(clk), .Q(X1[4])
         );
  FDS2L \RegX1_reg[20]  ( .CR(1'b1), .D(N23), .LD(n496), .CP(clk), .Q(
        RegX1[20]) );
  FDS2L \X1_reg[3]  ( .CR(1'b1), .D(RegX1[20]), .LD(n496), .CP(clk), .Q(X1[3])
         );
  FDS2L \RegX1_reg[19]  ( .CR(1'b1), .D(N22), .LD(n496), .CP(clk), .Q(
        RegX1[19]) );
  FDS2L \X1_reg[2]  ( .CR(1'b1), .D(RegX1[19]), .LD(n496), .CP(clk), .Q(X1[2])
         );
  FDS2L \RegX1_reg[18]  ( .CR(1'b1), .D(N21), .LD(n496), .CP(clk), .Q(
        RegX1[18]) );
  FDS2L \X1_reg[1]  ( .CR(1'b1), .D(RegX1[18]), .LD(n496), .CP(clk), .Q(X1[1])
         );
  FDS2L \RegX1_reg[17]  ( .CR(1'b1), .D(N20), .LD(n496), .CP(clk), .Q(
        RegX1[17]) );
  FDS2L \X1_reg[0]  ( .CR(1'b1), .D(RegX1[17]), .LD(n496), .CP(clk), .Q(X1[0])
         );
  FDS2L \X01_reg[15]  ( .CR(1'b1), .D(X0[15]), .LD(n496), .CP(clk), .Q(X01[15]) );
  FDS2L \X01_reg[14]  ( .CR(1'b1), .D(X0[14]), .LD(n496), .CP(clk), .Q(X01[14]) );
  FDS2L \X01_reg[13]  ( .CR(1'b1), .D(X0[13]), .LD(n496), .CP(clk), .Q(X01[13]) );
  FDS2L \X01_reg[12]  ( .CR(1'b1), .D(X0[12]), .LD(n496), .CP(clk), .Q(X01[12]) );
  FDS2L \X01_reg[11]  ( .CR(1'b1), .D(X0[11]), .LD(n495), .CP(clk), .Q(X01[11]) );
  FDS2L \X01_reg[10]  ( .CR(1'b1), .D(X0[10]), .LD(n495), .CP(clk), .Q(X01[10]) );
  FDS2L \X01_reg[9]  ( .CR(1'b1), .D(X0[9]), .LD(n495), .CP(clk), .Q(X01[9])
         );
  FDS2L \X01_reg[8]  ( .CR(1'b1), .D(X0[8]), .LD(n495), .CP(clk), .Q(X01[8])
         );
  FDS2L \X01_reg[7]  ( .CR(1'b1), .D(X0[7]), .LD(n495), .CP(clk), .Q(X01[7])
         );
  FDS2L \X01_reg[6]  ( .CR(1'b1), .D(X0[6]), .LD(n495), .CP(clk), .Q(X01[6])
         );
  FDS2L \X01_reg[5]  ( .CR(1'b1), .D(X0[5]), .LD(n495), .CP(clk), .Q(X01[5])
         );
  FDS2L \X01_reg[4]  ( .CR(1'b1), .D(X0[4]), .LD(n495), .CP(clk), .Q(X01[4])
         );
  FDS2L \X01_reg[3]  ( .CR(1'b1), .D(X0[3]), .LD(n495), .CP(clk), .Q(X01[3])
         );
  FDS2L \X01_reg[2]  ( .CR(1'b1), .D(X0[2]), .LD(n495), .CP(clk), .Q(X01[2])
         );
  FDS2L \X01_reg[1]  ( .CR(1'b1), .D(X0[1]), .LD(n495), .CP(clk), .Q(X01[1])
         );
  FDS2L \X01_reg[0]  ( .CR(1'b1), .D(X0[0]), .LD(n495), .CP(clk), .Q(X01[0])
         );
  FDS2L \X11_reg[15]  ( .CR(1'b1), .D(X1[15]), .LD(n494), .CP(clk), .Q(X11[15]) );
  FDS2L \X11_reg[14]  ( .CR(1'b1), .D(X1[14]), .LD(n494), .CP(clk), .Q(X11[14]) );
  FDS2L \X11_reg[13]  ( .CR(1'b1), .D(X1[13]), .LD(n494), .CP(clk), .Q(X11[13]) );
  FDS2L \X11_reg[12]  ( .CR(1'b1), .D(X1[12]), .LD(n494), .CP(clk), .Q(X11[12]) );
  FDS2L \X11_reg[11]  ( .CR(1'b1), .D(X1[11]), .LD(n494), .CP(clk), .Q(X11[11]) );
  FDS2L \X11_reg[10]  ( .CR(1'b1), .D(X1[10]), .LD(n494), .CP(clk), .Q(X11[10]) );
  FDS2L \X11_reg[9]  ( .CR(1'b1), .D(X1[9]), .LD(n493), .CP(clk), .Q(X11[9])
         );
  FDS2L \X11_reg[8]  ( .CR(1'b1), .D(X1[8]), .LD(n493), .CP(clk), .Q(X11[8])
         );
  FDS2L \X11_reg[7]  ( .CR(1'b1), .D(X1[7]), .LD(n493), .CP(clk), .Q(X11[7])
         );
  FDS2L \X11_reg[6]  ( .CR(1'b1), .D(X1[6]), .LD(n493), .CP(clk), .Q(X11[6])
         );
  FDS2L \X11_reg[5]  ( .CR(1'b1), .D(X1[5]), .LD(n493), .CP(clk), .Q(X11[5])
         );
  FDS2L \X11_reg[4]  ( .CR(1'b1), .D(X1[4]), .LD(n493), .CP(clk), .Q(X11[4])
         );
  FDS2L \X11_reg[3]  ( .CR(1'b1), .D(X1[3]), .LD(n492), .CP(clk), .Q(X11[3])
         );
  FDS2L \X11_reg[2]  ( .CR(1'b1), .D(X1[2]), .LD(n492), .CP(clk), .Q(X11[2])
         );
  FDS2L \X11_reg[1]  ( .CR(1'b1), .D(X1[1]), .LD(n492), .CP(clk), .Q(X11[1])
         );
  FDS2L \X11_reg[0]  ( .CR(1'b1), .D(X1[0]), .LD(n492), .CP(clk), .Q(X11[0])
         );
  FDS2L \LogIn_reg[43]  ( .CR(1'b1), .D(Taus1[27]), .LD(n490), .CP(clk), .Q(
        LogIn[43]) );
  FDS2L \LogIn_reg[34]  ( .CR(1'b1), .D(Taus1[18]), .LD(n489), .CP(clk), .Q(
        LogIn[34]) );
  FDS2L \LogIn_reg[22]  ( .CR(1'b1), .D(Taus1[6]), .LD(n488), .CP(clk), .Q(
        LogIn[22]) );
  FDS2L \LogIn_reg[21]  ( .CR(1'b1), .D(Taus1[5]), .LD(n488), .CP(clk), .Q(
        LogIn[21]) );
  FDS2L \LogIn_reg[17]  ( .CR(1'b1), .D(Taus1[1]), .LD(n488), .CP(clk), .Q(
        LogIn[17]) );
  FDS2L \LogIn_reg[40]  ( .CR(1'b1), .D(Taus1[24]), .LD(n490), .CP(clk), .Q(
        LogIn[40]) );
  FDS2L \LogIn_reg[42]  ( .CR(1'b1), .D(Taus1[26]), .LD(n490), .CP(clk), .Q(
        LogIn[42]) );
  FDS2L \LogIn_reg[13]  ( .CR(1'b1), .D(Taus2[29]), .LD(n488), .CP(clk), .Q(
        LogIn[13]) );
  FDS2L \LogIn_reg[10]  ( .CR(1'b1), .D(Taus2[26]), .LD(n487), .CP(clk), .Q(
        LogIn[10]) );
  FDS2L \LogIn_reg[9]  ( .CR(1'b1), .D(Taus2[25]), .LD(n487), .CP(clk), .Q(
        LogIn[9]) );
  FDS2L \LogIn_reg[7]  ( .CR(1'b1), .D(Taus2[23]), .LD(n487), .CP(clk), .Q(
        LogIn[7]) );
  FDS2L \LogIn_reg[6]  ( .CR(1'b1), .D(Taus2[22]), .LD(n487), .CP(clk), .Q(
        LogIn[6]) );
  FDS2L \LogIn_reg[8]  ( .CR(1'b1), .D(Taus2[24]), .LD(n487), .CP(clk), .Q(
        LogIn[8]) );
  FDS2L \LogIn_reg[5]  ( .CR(1'b1), .D(Taus2[21]), .LD(n487), .CP(clk), .Q(
        LogIn[5]) );
  FDS2L \LogIn_reg[4]  ( .CR(1'b1), .D(Taus2[20]), .LD(n487), .CP(clk), .Q(
        LogIn[4]) );
  FDS2L \LogIn_reg[3]  ( .CR(1'b1), .D(Taus2[19]), .LD(n487), .CP(clk), .Q(
        LogIn[3]) );
  FDS2L \LogIn_reg[35]  ( .CR(1'b1), .D(Taus1[19]), .LD(n489), .CP(clk), .Q(
        LogIn[35]) );
  FDS2L \LogIn_reg[44]  ( .CR(1'b1), .D(Taus1[28]), .LD(n490), .CP(clk), .Q(
        LogIn[44]) );
  FDS2L \LogIn_reg[23]  ( .CR(1'b1), .D(Taus1[7]), .LD(n488), .CP(clk), .Q(
        LogIn[23]) );
  FDS2L \LogIn_reg[24]  ( .CR(1'b1), .D(Taus1[8]), .LD(n489), .CP(clk), .Q(
        LogIn[24]) );
  FD1 \LogIn_reg[12]  ( .D(n483), .CP(clk), .Q(LogIn[12]) );
  FDS2L \LogIn_reg[45]  ( .CR(1'b1), .D(Taus1[29]), .LD(n490), .CP(clk), .Q(
        LogIn[45]) );
  FDS2L \LogIn_reg[14]  ( .CR(1'b1), .D(Taus2[30]), .LD(n488), .CP(clk), .Q(
        LogIn[14]) );
  FD1 \LogIn_reg[18]  ( .D(n482), .CP(clk), .Q(LogIn[18]) );
  FDS2L \LogIn_reg[46]  ( .CR(1'b1), .D(Taus1[30]), .LD(n490), .CP(clk), .Q(
        LogIn[46]) );
  FDS2L \LogIn_reg[36]  ( .CR(1'b1), .D(Taus1[20]), .LD(n490), .CP(clk), .Q(
        LogIn[36]) );
  FDS2L \LogIn_reg[19]  ( .CR(1'b1), .D(Taus1[3]), .LD(n488), .CP(clk), .Q(
        LogIn[19]) );
  FDS2L \LogIn_reg[25]  ( .CR(1'b1), .D(Taus1[9]), .LD(n489), .CP(clk), .Q(
        LogIn[25]) );
  FD1 \LogIn_reg[20]  ( .D(n481), .CP(clk), .Q(LogIn[20]) );
  FDS2L \LogIn_reg[41]  ( .CR(1'b1), .D(Taus1[25]), .LD(n490), .CP(clk), .Q(
        LogIn[41]) );
  FDS2L \LogIn_reg[39]  ( .CR(1'b1), .D(Taus1[23]), .LD(n490), .CP(clk), .Q(
        LogIn[39]) );
  FDS2L \LogIn_reg[38]  ( .CR(1'b1), .D(Taus1[22]), .LD(n490), .CP(clk), .Q(
        LogIn[38]) );
  FDS2L \LogIn_reg[37]  ( .CR(1'b1), .D(Taus1[21]), .LD(n490), .CP(clk), .Q(
        LogIn[37]) );
  FDS2L \LogIn_reg[33]  ( .CR(1'b1), .D(Taus1[17]), .LD(n489), .CP(clk), .Q(
        LogIn[33]) );
  FDS2L \LogIn_reg[31]  ( .CR(1'b1), .D(Taus1[15]), .LD(n489), .CP(clk), .Q(
        LogIn[31]) );
  FDS2L \LogIn_reg[30]  ( .CR(1'b1), .D(Taus1[14]), .LD(n489), .CP(clk), .Q(
        LogIn[30]) );
  FDS2L \LogIn_reg[29]  ( .CR(1'b1), .D(Taus1[13]), .LD(n489), .CP(clk), .Q(
        LogIn[29]) );
  FDS2L \LogIn_reg[28]  ( .CR(1'b1), .D(Taus1[12]), .LD(n489), .CP(clk), .Q(
        LogIn[28]) );
  FDS2L \LogIn_reg[16]  ( .CR(1'b1), .D(Taus1[0]), .LD(n488), .CP(clk), .Q(
        LogIn[16]) );
  FDS2L \LogIn_reg[15]  ( .CR(1'b1), .D(Taus2[31]), .LD(n488), .CP(clk), .Q(
        LogIn[15]) );
  FD1 \LogIn_reg[11]  ( .D(n485), .CP(clk), .Q(LogIn[11]) );
  IVP U481 ( .A(n534), .Z(n488) );
  IVP U482 ( .A(n534), .Z(n487) );
  IVP U483 ( .A(n534), .Z(n489) );
  IVP U484 ( .A(n534), .Z(n492) );
  IVP U485 ( .A(n534), .Z(n493) );
  IVP U486 ( .A(n534), .Z(n494) );
  IVP U487 ( .A(n533), .Z(n495) );
  IVP U488 ( .A(n533), .Z(n496) );
  IVP U489 ( .A(n533), .Z(n497) );
  IVP U490 ( .A(n533), .Z(n498) );
  IVP U491 ( .A(n533), .Z(n499) );
  IVP U492 ( .A(n533), .Z(n500) );
  IVP U493 ( .A(n533), .Z(n501) );
  IVP U494 ( .A(n533), .Z(n502) );
  IVP U495 ( .A(n533), .Z(n503) );
  IVP U496 ( .A(n533), .Z(n504) );
  IVP U497 ( .A(n533), .Z(n505) );
  IVP U498 ( .A(n533), .Z(n506) );
  IVP U499 ( .A(n532), .Z(n507) );
  IVP U500 ( .A(n532), .Z(n508) );
  IVP U501 ( .A(n532), .Z(n509) );
  IVP U502 ( .A(n532), .Z(n510) );
  IVP U503 ( .A(n532), .Z(n511) );
  IVP U504 ( .A(n532), .Z(n512) );
  IVP U505 ( .A(n532), .Z(n513) );
  IVP U506 ( .A(n532), .Z(n514) );
  IVP U507 ( .A(n532), .Z(n515) );
  IVP U508 ( .A(n532), .Z(n516) );
  IVP U509 ( .A(n532), .Z(n517) );
  IVP U510 ( .A(n532), .Z(n518) );
  IVP U511 ( .A(n531), .Z(n519) );
  IVP U512 ( .A(n531), .Z(n520) );
  IVP U513 ( .A(n531), .Z(n521) );
  IVP U514 ( .A(n531), .Z(n522) );
  IVP U515 ( .A(n531), .Z(n523) );
  IVP U516 ( .A(n531), .Z(n524) );
  IVP U517 ( .A(n531), .Z(n525) );
  IVP U518 ( .A(n531), .Z(n526) );
  IVP U519 ( .A(n531), .Z(n527) );
  IVP U520 ( .A(n531), .Z(n528) );
  IVP U521 ( .A(n534), .Z(n490) );
  IVP U522 ( .A(n531), .Z(n529) );
  IVP U523 ( .A(n534), .Z(n491) );
  IVP U524 ( .A(n531), .Z(n530) );
  IVP U525 ( .A(n535), .Z(n533) );
  IVP U526 ( .A(n535), .Z(n532) );
  IVP U527 ( .A(n535), .Z(n531) );
  IVP U528 ( .A(n535), .Z(n534) );
  MUX21H U529 ( .A(LogIn[20]), .B(Taus1[4]), .S(n488), .Z(n481) );
  MUX21H U530 ( .A(LogIn[18]), .B(Taus1[2]), .S(n488), .Z(n482) );
  MUX21H U531 ( .A(LogIn[12]), .B(Taus2[28]), .S(n488), .Z(n483) );
  MUX21H U532 ( .A(LogIn[2]), .B(Taus2[18]), .S(n487), .Z(n484) );
  MUX21H U533 ( .A(LogIn[11]), .B(Taus2[27]), .S(n487), .Z(n485) );
  MUX21H U534 ( .A(LogIn[27]), .B(Taus1[11]), .S(n489), .Z(n486) );
  IVA U535 ( .A(reset), .Z(n535) );
endmodule

