
module Taus ( clk, reset, Tout );
  output [31:0] Tout;
  input clk, reset;
  wire   N44, N46, N77, N108, N109, N110, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n88, n108, n110, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158;
  wire   [31:0] s0;
  wire   [31:0] s1;
  wire   [31:0] s2;

  FD1 \s0_reg[1]  ( .D(N77), .CP(clk), .Q(s0[1]) );
  FDS2 \s0_reg[13]  ( .CR(n153), .D(s0[1]), .CP(clk), .Q(s0[13]), .QN(n42) );
  FDS2 \s0_reg[25]  ( .CR(n153), .D(s0[13]), .CP(clk), .Q(s0[25]) );
  FDS2 \s0_reg[7]  ( .CR(n153), .D(n152), .CP(clk), .Q(s0[7]) );
  FDS2 \s0_reg[19]  ( .CR(n153), .D(s0[7]), .CP(clk), .Q(s0[19]), .QN(n36) );
  FDS2 \s0_reg[31]  ( .CR(n153), .D(s0[19]), .CP(clk), .Q(s0[31]) );
  FDS2 \s0_reg[12]  ( .CR(n153), .D(n151), .CP(clk), .Q(s0[12]), .QN(n43) );
  FDS2 \s0_reg[24]  ( .CR(n153), .D(s0[12]), .CP(clk), .Q(s0[24]) );
  FDS2 \s0_reg[6]  ( .CR(n153), .D(n150), .CP(clk), .Q(s0[6]) );
  FDS2 \s0_reg[18]  ( .CR(n153), .D(s0[6]), .CP(clk), .Q(s0[18]), .QN(n37) );
  FDS2 \s0_reg[30]  ( .CR(n153), .D(s0[18]), .CP(clk), .Q(s0[30]) );
  FDS2 \s0_reg[11]  ( .CR(n153), .D(n149), .CP(clk), .Q(s0[11]) );
  FDS2 \s0_reg[23]  ( .CR(n153), .D(s0[11]), .CP(clk), .Q(s0[23]) );
  FDS2 \s0_reg[5]  ( .CR(n154), .D(n148), .CP(clk), .Q(s0[5]) );
  FDS2 \s0_reg[17]  ( .CR(n154), .D(s0[5]), .CP(clk), .Q(s0[17]), .QN(n38) );
  FDS2 \s0_reg[29]  ( .CR(n154), .D(s0[17]), .CP(clk), .Q(s0[29]) );
  FDS2 \s0_reg[10]  ( .CR(n154), .D(n147), .CP(clk), .Q(s0[10]) );
  FDS2 \s0_reg[22]  ( .CR(n154), .D(s0[10]), .CP(clk), .Q(s0[22]) );
  FDS2 \s0_reg[4]  ( .CR(n154), .D(n146), .CP(clk), .Q(s0[4]) );
  FDS2 \s0_reg[16]  ( .CR(n154), .D(s0[4]), .CP(clk), .Q(s0[16]), .QN(n39) );
  FDS2 \s0_reg[28]  ( .CR(n154), .D(s0[16]), .CP(clk), .Q(s0[28]) );
  FDS2 \s0_reg[9]  ( .CR(n154), .D(n145), .CP(clk), .Q(s0[9]) );
  FDS2 \s0_reg[21]  ( .CR(n154), .D(s0[9]), .CP(clk), .Q(s0[21]) );
  FDS2 \s0_reg[3]  ( .CR(n154), .D(n144), .CP(clk), .Q(s0[3]) );
  FDS2 \s0_reg[15]  ( .CR(n154), .D(s0[3]), .CP(clk), .Q(s0[15]), .QN(n40) );
  FDS2 \s0_reg[27]  ( .CR(n154), .D(s0[15]), .CP(clk), .Q(s0[27]) );
  FDS2 \s0_reg[8]  ( .CR(n154), .D(n143), .CP(clk), .Q(s0[8]) );
  FDS2 \s0_reg[20]  ( .CR(n154), .D(s0[8]), .CP(clk), .Q(s0[20]) );
  FDS2 \s0_reg[2]  ( .CR(n154), .D(n142), .CP(clk), .Q(s0[2]) );
  FDS2 \s0_reg[14]  ( .CR(n154), .D(s0[2]), .CP(clk), .Q(s0[14]), .QN(n41) );
  FDS2 \s0_reg[26]  ( .CR(n154), .D(s0[14]), .CP(clk), .Q(s0[26]) );
  FDS2 \s0_reg[0]  ( .CR(n154), .D(n141), .CP(clk), .Q(s0[0]) );
  FDS2 \s2_reg[4]  ( .CR(n154), .D(n124), .CP(clk), .Q(s2[4]) );
  FDS2 \s2_reg[21]  ( .CR(n154), .D(s2[4]), .CP(clk), .Q(s2[21]) );
  FDS2 \s2_reg[10]  ( .CR(n154), .D(n140), .CP(clk), .Q(s2[10]) );
  FDS2 \s2_reg[27]  ( .CR(n154), .D(s2[10]), .CP(clk), .Q(s2[27]) );
  FDS2 \s2_reg[16]  ( .CR(n154), .D(n139), .CP(clk), .Q(s2[16]) );
  FDS2 \s2_reg[5]  ( .CR(n155), .D(n123), .CP(clk), .Q(s2[5]) );
  FDS2 \s2_reg[22]  ( .CR(n155), .D(s2[5]), .CP(clk), .Q(s2[22]) );
  FDS2 \s2_reg[11]  ( .CR(n155), .D(n138), .CP(clk), .Q(s2[11]) );
  FDS2 \s2_reg[28]  ( .CR(n155), .D(s2[11]), .CP(clk), .Q(s2[28]) );
  FDS2 \s2_reg[17]  ( .CR(n155), .D(n137), .CP(clk), .Q(s2[17]) );
  FDS2 \s2_reg[6]  ( .CR(n155), .D(n122), .CP(clk), .Q(s2[6]) );
  FDS2 \s2_reg[23]  ( .CR(n155), .D(s2[6]), .CP(clk), .Q(s2[23]) );
  FDS2 \s2_reg[12]  ( .CR(n155), .D(n136), .CP(clk), .Q(s2[12]) );
  FDS2 \s2_reg[29]  ( .CR(n155), .D(s2[12]), .CP(clk), .Q(s2[29]) );
  FDS2 \s2_reg[18]  ( .CR(n155), .D(n135), .CP(clk), .Q(s2[18]) );
  FDS2 \s2_reg[7]  ( .CR(n155), .D(n134), .CP(clk), .Q(s2[7]) );
  FDS2 \s2_reg[24]  ( .CR(n155), .D(s2[7]), .CP(clk), .Q(s2[24]) );
  FDS2 \s2_reg[13]  ( .CR(n155), .D(n133), .CP(clk), .Q(s2[13]) );
  FDS2 \s2_reg[30]  ( .CR(n155), .D(s2[13]), .CP(clk), .Q(s2[30]) );
  FDS2 \s2_reg[19]  ( .CR(n155), .D(n132), .CP(clk), .Q(s2[19]) );
  FDS2 \s2_reg[8]  ( .CR(n155), .D(n131), .CP(clk), .Q(s2[8]) );
  FDS2 \s2_reg[25]  ( .CR(n155), .D(s2[8]), .CP(clk), .Q(s2[25]) );
  FDS2 \s2_reg[14]  ( .CR(n155), .D(n130), .CP(clk), .Q(s2[14]) );
  FDS2 \s2_reg[31]  ( .CR(n155), .D(s2[14]), .CP(clk), .Q(s2[31]) );
  FDS2 \s2_reg[20]  ( .CR(n155), .D(n129), .CP(clk), .Q(s2[20]) );
  FDS2 \s2_reg[9]  ( .CR(n155), .D(n128), .CP(clk), .Q(s2[9]) );
  FDS2 \s2_reg[26]  ( .CR(n155), .D(s2[9]), .CP(clk), .Q(s2[26]) );
  FDS2 \s2_reg[15]  ( .CR(n155), .D(n127), .CP(clk), .Q(s2[15]) );
  FDS2 \s2_reg[3]  ( .CR(n155), .D(n121), .CP(clk), .Q(s2[3]) );
  FD1 \s2_reg[2]  ( .D(N46), .CP(clk), .Q(s2[2]) );
  FDS2 \s2_reg[1]  ( .CR(n156), .D(n120), .CP(clk), .Q(s2[1]) );
  FD1 \s2_reg[0]  ( .D(N44), .CP(clk), .Q(s2[0]) );
  FDS2 \s1_reg[3]  ( .CR(n156), .D(n119), .CP(clk), .Q(s1[3]) );
  FDS2 \s1_reg[7]  ( .CR(n156), .D(s1[3]), .CP(clk), .Q(s1[7]) );
  FDS2 \s1_reg[11]  ( .CR(n156), .D(s1[7]), .CP(clk), .Q(s1[11]) );
  FDS2 \s1_reg[15]  ( .CR(n156), .D(s1[11]), .CP(clk), .Q(s1[15]) );
  FDS2 \s1_reg[19]  ( .CR(n156), .D(s1[15]), .CP(clk), .Q(s1[19]) );
  FDS2 \s1_reg[23]  ( .CR(n156), .D(s1[19]), .CP(clk), .Q(s1[23]) );
  FDS2 \s1_reg[27]  ( .CR(n156), .D(s1[23]), .CP(clk), .Q(s1[27]) );
  FDS2 \s1_reg[31]  ( .CR(n156), .D(s1[27]), .CP(clk), .Q(s1[31]) );
  FDS2 \s1_reg[4]  ( .CR(n156), .D(n118), .CP(clk), .Q(s1[4]) );
  FDS2 \s1_reg[8]  ( .CR(n156), .D(s1[4]), .CP(clk), .Q(s1[8]) );
  FDS2 \s1_reg[12]  ( .CR(n156), .D(s1[8]), .CP(clk), .Q(s1[12]) );
  FDS2 \s1_reg[16]  ( .CR(n156), .D(s1[12]), .CP(clk), .Q(s1[16]) );
  FDS2 \s1_reg[20]  ( .CR(n156), .D(s1[16]), .CP(clk), .Q(s1[20]) );
  FDS2 \s1_reg[24]  ( .CR(n156), .D(s1[20]), .CP(clk), .Q(s1[24]) );
  FDS2 \s1_reg[28]  ( .CR(n156), .D(s1[24]), .CP(clk), .Q(s1[28]) );
  FDS2 \s1_reg[5]  ( .CR(n156), .D(n126), .CP(clk), .Q(s1[5]) );
  FDS2 \s1_reg[9]  ( .CR(n156), .D(s1[5]), .CP(clk), .Q(s1[9]) );
  FDS2 \s1_reg[13]  ( .CR(n156), .D(s1[9]), .CP(clk), .Q(s1[13]) );
  FDS2 \s1_reg[17]  ( .CR(n156), .D(s1[13]), .CP(clk), .Q(s1[17]) );
  FDS2 \s1_reg[21]  ( .CR(n156), .D(s1[17]), .CP(clk), .Q(s1[21]) );
  FDS2 \s1_reg[25]  ( .CR(n156), .D(s1[21]), .CP(clk), .Q(s1[25]) );
  FDS2 \s1_reg[29]  ( .CR(n156), .D(s1[25]), .CP(clk), .Q(s1[29]) );
  FDS2 \s1_reg[6]  ( .CR(n156), .D(n125), .CP(clk), .Q(s1[6]) );
  FDS2 \s1_reg[10]  ( .CR(n157), .D(s1[6]), .CP(clk), .Q(s1[10]) );
  FDS2 \s1_reg[14]  ( .CR(n157), .D(s1[10]), .CP(clk), .Q(s1[14]) );
  FDS2 \s1_reg[18]  ( .CR(n157), .D(s1[14]), .CP(clk), .Q(s1[18]) );
  FDS2 \s1_reg[22]  ( .CR(n157), .D(s1[18]), .CP(clk), .Q(s1[22]) );
  FDS2 \s1_reg[26]  ( .CR(n157), .D(s1[22]), .CP(clk), .Q(s1[26]) );
  FDS2 \s1_reg[30]  ( .CR(n157), .D(s1[26]), .CP(clk), .Q(s1[30]) );
  FD1 \s1_reg[2]  ( .D(N110), .CP(clk), .Q(s1[2]) );
  FD1 \s1_reg[1]  ( .D(N109), .CP(clk), .Q(s1[1]) );
  FD1 \s1_reg[0]  ( .D(N108), .CP(clk), .Q(s1[0]) );
  IVP U150 ( .A(n158), .Z(n156) );
  IVP U151 ( .A(n158), .Z(n155) );
  IVP U152 ( .A(n158), .Z(n154) );
  IVP U153 ( .A(n158), .Z(n153) );
  EO U154 ( .A(s0[11]), .B(n74), .Z(Tout[11]) );
  EO U155 ( .A(s2[11]), .B(s1[11]), .Z(n74) );
  ND2 U156 ( .A(n110), .B(n153), .Z(N44) );
  EN U157 ( .A(s2[8]), .B(s2[11]), .Z(n110) );
  EO U158 ( .A(s1[29]), .B(s1[27]), .Z(n118) );
  EO U159 ( .A(s1[28]), .B(s1[26]), .Z(n119) );
  EO U160 ( .A(s2[9]), .B(s2[12]), .Z(n120) );
  EO U161 ( .A(s2[11]), .B(s2[14]), .Z(n121) );
  EO U162 ( .A(s2[17]), .B(s2[14]), .Z(n122) );
  EO U163 ( .A(s2[16]), .B(s2[13]), .Z(n123) );
  EO U164 ( .A(s2[15]), .B(s2[12]), .Z(n124) );
  ND2 U165 ( .A(n117), .B(n153), .Z(N108) );
  EN U166 ( .A(s1[23]), .B(s1[25]), .Z(n117) );
  ND2 U167 ( .A(n116), .B(n153), .Z(N109) );
  EN U168 ( .A(s1[24]), .B(s1[26]), .Z(n116) );
  ND2 U169 ( .A(n115), .B(n153), .Z(N110) );
  EN U170 ( .A(s1[25]), .B(s1[27]), .Z(n115) );
  ND2 U171 ( .A(n108), .B(n153), .Z(N46) );
  EN U172 ( .A(s2[10]), .B(s2[13]), .Z(n108) );
  ND2 U173 ( .A(n88), .B(n153), .Z(N77) );
  EN U174 ( .A(s0[20]), .B(s0[7]), .Z(n88) );
  EN U175 ( .A(n43), .B(n73), .Z(Tout[12]) );
  EO U176 ( .A(s2[12]), .B(s1[12]), .Z(n73) );
  EN U177 ( .A(n42), .B(n72), .Z(Tout[13]) );
  EO U178 ( .A(s2[13]), .B(s1[13]), .Z(n72) );
  EN U179 ( .A(n41), .B(n71), .Z(Tout[14]) );
  EO U180 ( .A(s2[14]), .B(s1[14]), .Z(n71) );
  EO U181 ( .A(s0[25]), .B(n59), .Z(Tout[25]) );
  EO U182 ( .A(s2[25]), .B(s1[25]), .Z(n59) );
  EO U183 ( .A(s0[26]), .B(n58), .Z(Tout[26]) );
  EO U184 ( .A(s2[26]), .B(s1[26]), .Z(n58) );
  EO U185 ( .A(s0[27]), .B(n57), .Z(Tout[27]) );
  EO U186 ( .A(s2[27]), .B(s1[27]), .Z(n57) );
  IVP U187 ( .A(n44), .Z(n158) );
  IVP U188 ( .A(reset), .Z(n44) );
  EO U189 ( .A(s1[29]), .B(s1[31]), .Z(n125) );
  EO U190 ( .A(s1[28]), .B(s1[30]), .Z(n126) );
  EO U191 ( .A(s2[23]), .B(s2[26]), .Z(n127) );
  EO U192 ( .A(s2[17]), .B(s2[20]), .Z(n128) );
  EO U193 ( .A(s2[28]), .B(s2[31]), .Z(n129) );
  EO U194 ( .A(s2[22]), .B(s2[25]), .Z(n130) );
  EO U195 ( .A(s2[16]), .B(s2[19]), .Z(n131) );
  EO U196 ( .A(s2[27]), .B(s2[30]), .Z(n132) );
  EO U197 ( .A(s2[21]), .B(s2[24]), .Z(n133) );
  EO U198 ( .A(s2[15]), .B(s2[18]), .Z(n134) );
  EO U199 ( .A(s2[26]), .B(s2[29]), .Z(n135) );
  EO U200 ( .A(s2[20]), .B(s2[23]), .Z(n136) );
  EO U201 ( .A(s2[25]), .B(s2[28]), .Z(n137) );
  EO U202 ( .A(s2[19]), .B(s2[22]), .Z(n138) );
  EO U203 ( .A(s2[24]), .B(s2[27]), .Z(n139) );
  EO U204 ( .A(s2[18]), .B(s2[21]), .Z(n140) );
  EO U205 ( .A(s0[19]), .B(s0[6]), .Z(n141) );
  EO U206 ( .A(s0[21]), .B(s0[8]), .Z(n142) );
  EO U207 ( .A(s0[14]), .B(s0[27]), .Z(n143) );
  EO U208 ( .A(s0[22]), .B(s0[9]), .Z(n144) );
  EO U209 ( .A(s0[15]), .B(s0[28]), .Z(n145) );
  EO U210 ( .A(s0[10]), .B(s0[23]), .Z(n146) );
  EO U211 ( .A(s0[16]), .B(s0[29]), .Z(n147) );
  EO U212 ( .A(s0[11]), .B(s0[24]), .Z(n148) );
  EO U213 ( .A(s0[17]), .B(s0[30]), .Z(n149) );
  EO U214 ( .A(s0[12]), .B(s0[25]), .Z(n150) );
  EO U215 ( .A(s0[18]), .B(s0[31]), .Z(n151) );
  EO U216 ( .A(s0[13]), .B(s0[26]), .Z(n152) );
  EO U217 ( .A(s0[0]), .B(n76), .Z(Tout[0]) );
  EO U218 ( .A(s2[0]), .B(s1[0]), .Z(n76) );
  EO U219 ( .A(s0[1]), .B(n65), .Z(Tout[1]) );
  EO U220 ( .A(s2[1]), .B(s1[1]), .Z(n65) );
  EO U221 ( .A(s0[2]), .B(n54), .Z(Tout[2]) );
  EO U222 ( .A(s2[2]), .B(s1[2]), .Z(n54) );
  EO U223 ( .A(s0[3]), .B(n51), .Z(Tout[3]) );
  EO U224 ( .A(s2[3]), .B(s1[3]), .Z(n51) );
  EO U225 ( .A(s0[4]), .B(n50), .Z(Tout[4]) );
  EO U226 ( .A(s2[4]), .B(s1[4]), .Z(n50) );
  EO U227 ( .A(s0[5]), .B(n49), .Z(Tout[5]) );
  EO U228 ( .A(s2[5]), .B(s1[5]), .Z(n49) );
  EO U229 ( .A(s0[6]), .B(n48), .Z(Tout[6]) );
  EO U230 ( .A(s2[6]), .B(s1[6]), .Z(n48) );
  EO U231 ( .A(s0[7]), .B(n47), .Z(Tout[7]) );
  EO U232 ( .A(s2[7]), .B(s1[7]), .Z(n47) );
  EO U233 ( .A(s0[8]), .B(n46), .Z(Tout[8]) );
  EO U234 ( .A(s2[8]), .B(s1[8]), .Z(n46) );
  EO U235 ( .A(s0[9]), .B(n45), .Z(Tout[9]) );
  EO U236 ( .A(s2[9]), .B(s1[9]), .Z(n45) );
  EO U237 ( .A(s0[10]), .B(n75), .Z(Tout[10]) );
  EO U238 ( .A(s2[10]), .B(s1[10]), .Z(n75) );
  EN U239 ( .A(n40), .B(n70), .Z(Tout[15]) );
  EO U240 ( .A(s2[15]), .B(s1[15]), .Z(n70) );
  EN U241 ( .A(n39), .B(n69), .Z(Tout[16]) );
  EO U242 ( .A(s2[16]), .B(s1[16]), .Z(n69) );
  EN U243 ( .A(n38), .B(n68), .Z(Tout[17]) );
  EO U244 ( .A(s2[17]), .B(s1[17]), .Z(n68) );
  EN U245 ( .A(n37), .B(n67), .Z(Tout[18]) );
  EO U246 ( .A(s2[18]), .B(s1[18]), .Z(n67) );
  EN U247 ( .A(n36), .B(n66), .Z(Tout[19]) );
  EO U248 ( .A(s2[19]), .B(s1[19]), .Z(n66) );
  EO U249 ( .A(s0[20]), .B(n64), .Z(Tout[20]) );
  EO U250 ( .A(s2[20]), .B(s1[20]), .Z(n64) );
  EO U251 ( .A(s0[21]), .B(n63), .Z(Tout[21]) );
  EO U252 ( .A(s2[21]), .B(s1[21]), .Z(n63) );
  EO U253 ( .A(s0[22]), .B(n62), .Z(Tout[22]) );
  EO U254 ( .A(s2[22]), .B(s1[22]), .Z(n62) );
  EO U255 ( .A(s0[23]), .B(n61), .Z(Tout[23]) );
  EO U256 ( .A(s2[23]), .B(s1[23]), .Z(n61) );
  EO U257 ( .A(s0[24]), .B(n60), .Z(Tout[24]) );
  EO U258 ( .A(s2[24]), .B(s1[24]), .Z(n60) );
  EO U259 ( .A(s0[28]), .B(n56), .Z(Tout[28]) );
  EO U260 ( .A(s2[28]), .B(s1[28]), .Z(n56) );
  EO U261 ( .A(s0[29]), .B(n55), .Z(Tout[29]) );
  EO U262 ( .A(s2[29]), .B(s1[29]), .Z(n55) );
  EO U263 ( .A(s0[30]), .B(n53), .Z(Tout[30]) );
  EO U264 ( .A(s2[30]), .B(s1[30]), .Z(n53) );
  EO U265 ( .A(s0[31]), .B(n52), .Z(Tout[31]) );
  EO U266 ( .A(s2[31]), .B(s1[31]), .Z(n52) );
  IVA U267 ( .A(n158), .Z(n157) );
endmodule

