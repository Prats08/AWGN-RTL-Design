
module SQRT_POLY_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;

  wire   [13:1] carry;

  FA1A U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA1A U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(SUM[13]), .S(SUM[12])
         );
  FA1A U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA1A U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  FA1A U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA1A U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA1A U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA1A U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA1A U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA1A U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA1A U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA1A U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  EO U1 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
  AN2P U2 ( .A(A[0]), .B(B[0]), .Z(carry[1]) );
endmodule


module SQRT_POLY_DW01_add_2 ( A, B, CI, SUM, CO );
  input [40:0] A;
  input [40:0] B;
  output [40:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271;

  AO7P U2 ( .A(n238), .B(n239), .C(n240), .Z(n237) );
  IVDA U3 ( .A(n175), .Z(n1) );
  AO7P U4 ( .A(n47), .B(n48), .C(n49), .Z(n45) );
  B4I U5 ( .A(n85), .Z(n47) );
  IVP U6 ( .A(B[16]), .Z(n265) );
  B2I U7 ( .A(n132), .Z2(n2) );
  AO6 U8 ( .A(n162), .B(n141), .C(n144), .Z(n151) );
  ND5 U9 ( .A(B[11]), .B(A[11]), .C(n254), .D(n20), .E(n256), .Z(n30) );
  ND2 U10 ( .A(n65), .B(n66), .Z(n56) );
  ND2 U11 ( .A(n86), .B(n87), .Z(n75) );
  ND2 U12 ( .A(B[32]), .B(A[32]), .Z(n68) );
  ND2 U13 ( .A(n116), .B(n166), .Z(n141) );
  ND2 U14 ( .A(n59), .B(n60), .Z(n51) );
  ND2 U15 ( .A(B[33]), .B(A[33]), .Z(n80) );
  IVP U16 ( .A(B[29]), .Z(n129) );
  ND2 U17 ( .A(n268), .B(n269), .Z(n262) );
  ND2 U18 ( .A(n270), .B(n271), .Z(n261) );
  IVDA U19 ( .A(A[12]), .Y(n44), .Z(n43) );
  ND2 U20 ( .A(n224), .B(n225), .Z(n219) );
  NR3 U21 ( .A(n116), .B(n112), .C(n117), .Z(n109) );
  EN U22 ( .A(n64), .B(n40), .Z(SUM[35]) );
  EN U23 ( .A(n246), .B(n247), .Z(SUM[21]) );
  EO U24 ( .A(n194), .B(n195), .Z(SUM[26]) );
  EN U25 ( .A(n187), .B(n188), .Z(SUM[27]) );
  EO U26 ( .A(n148), .B(n149), .Z(SUM[30]) );
  AO6 U27 ( .A(n140), .B(n141), .C(n142), .Z(n139) );
  IVDA U28 ( .A(n101), .Z(n3) );
  AN2P U29 ( .A(n56), .B(n51), .Z(n4) );
  AN3 U30 ( .A(n189), .B(n190), .C(n177), .Z(n5) );
  IVDA U31 ( .A(n126), .Y(n6), .Z(n7) );
  AN2P U32 ( .A(n260), .B(n131), .Z(n8) );
  AN2P U33 ( .A(n260), .B(n131), .Z(n9) );
  OR2 U34 ( .A(A[22]), .B(B[22]), .Z(n31) );
  IVDA U35 ( .A(n216), .Y(n233) );
  IVDA U36 ( .A(n174), .Z(n10) );
  ND2P U37 ( .A(n170), .B(n171), .Z(n106) );
  IVDAP U38 ( .A(A[28]), .Y(n12), .Z(n11) );
  ND2 U39 ( .A(n260), .B(n131), .Z(n13) );
  IVDA U40 ( .A(n222), .Y(n15) );
  NR2P U41 ( .A(A[21]), .B(B[21]), .Z(n222) );
  OR2 U42 ( .A(A[21]), .B(B[21]), .Z(n217) );
  IV U43 ( .A(n130), .Z(n16) );
  IV U44 ( .A(A[24]), .Z(n182) );
  B3I U45 ( .A(n245), .Z1(n18), .Z2(n17) );
  IV U46 ( .A(B[14]), .Z(n258) );
  IV U47 ( .A(B[12]), .Z(n257) );
  IV U48 ( .A(A[26]), .Z(n197) );
  AO3 U49 ( .A(n207), .B(n208), .C(n161), .D(n8), .Z(n202) );
  ND4P U50 ( .A(n178), .B(n179), .C(n180), .D(n175), .Z(n19) );
  AO3P U51 ( .A(n118), .B(n119), .C(n120), .D(n121), .Z(n88) );
  NR3P U52 ( .A(n19), .B(n22), .C(n98), .Z(n121) );
  OR2 U53 ( .A(A[22]), .B(B[22]), .Z(n216) );
  IV U54 ( .A(A[18]), .Z(n269) );
  IV U55 ( .A(A[25]), .Z(n184) );
  OR2 U56 ( .A(B[13]), .B(A[13]), .Z(n20) );
  AN2 U57 ( .A(n213), .B(n214), .Z(n212) );
  IVDA U58 ( .A(n214), .Y(n232), .Z(n14) );
  AN3P U59 ( .A(n156), .B(n157), .C(n23), .Z(n21) );
  ND4 U60 ( .A(n261), .B(n262), .C(n263), .D(n264), .Z(n22) );
  AO3P U61 ( .A(n207), .B(n160), .C(n161), .D(n9), .Z(n23) );
  IV U62 ( .A(n47), .Z(n24) );
  IVDA U63 ( .A(n3), .Y(n25) );
  IVAP U64 ( .A(n97), .Z(n101) );
  IV U65 ( .A(n93), .Z(n241) );
  NR2P U66 ( .A(n236), .B(n237), .Z(n235) );
  IVDAP U67 ( .A(A[31]), .Y(n27), .Z(n26) );
  IV U68 ( .A(B[17]), .Z(n270) );
  ND2P U69 ( .A(n129), .B(n130), .Z(n28) );
  B5I U70 ( .A(A[29]), .Z(n130) );
  ND2P U71 ( .A(n2), .B(n133), .Z(n208) );
  IVAP U72 ( .A(n122), .Z(n260) );
  ND3 U73 ( .A(n156), .B(n157), .C(n202), .Z(n29) );
  EN U74 ( .A(n24), .B(n36), .Z(SUM[32]) );
  ND3 U75 ( .A(n92), .B(n93), .C(n94), .Z(n91) );
  IV U76 ( .A(n63), .Z(n55) );
  ND4P U77 ( .A(n101), .B(n102), .C(n103), .D(n104), .Z(n100) );
  AN2 U78 ( .A(A[21]), .B(B[21]), .Z(n215) );
  ND2P U79 ( .A(n265), .B(n42), .Z(n264) );
  IVDAP U80 ( .A(A[16]), .Y(n42), .Z(n41) );
  AO3P U81 ( .A(n172), .B(n173), .C(n174), .D(n175), .Z(n171) );
  AO7P U82 ( .A(n47), .B(n63), .C(n67), .Z(n64) );
  ND5 U83 ( .A(B[11]), .B(A[11]), .C(n254), .D(n255), .E(n256), .Z(n133) );
  IVP U84 ( .A(n193), .Z(n172) );
  ND2P U85 ( .A(n31), .B(n217), .Z(n209) );
  ND2P U86 ( .A(n215), .B(n216), .Z(n211) );
  OR2P U87 ( .A(A[29]), .B(B[29]), .Z(n146) );
  IV U88 ( .A(n52), .Z(n67) );
  AO2P U89 ( .A(n50), .B(n51), .C(n4), .D(n52), .Z(n49) );
  ND4P U90 ( .A(n124), .B(n125), .C(n126), .D(n111), .Z(n32) );
  NR2P U91 ( .A(n107), .B(n96), .Z(n105) );
  IVA U92 ( .A(B[36]), .Z(n59) );
  ND2P U93 ( .A(n127), .B(n128), .Z(n125) );
  AO3 U94 ( .A(n153), .B(n154), .C(n145), .D(n146), .Z(n152) );
  ND3 U95 ( .A(n75), .B(n73), .C(n74), .Z(n63) );
  NR2P U96 ( .A(A[23]), .B(B[23]), .Z(n223) );
  ND2 U97 ( .A(B[22]), .B(A[22]), .Z(n214) );
  EO U98 ( .A(B[37]), .B(A[37]), .Z(n46) );
  ENP U99 ( .A(n136), .B(n33), .Z(SUM[31]) );
  ENP U100 ( .A(n203), .B(n204), .Z(SUM[25]) );
  ENP U101 ( .A(n167), .B(n34), .Z(SUM[28]) );
  EOP U102 ( .A(n163), .B(n164), .Z(SUM[29]) );
  ENP U103 ( .A(n227), .B(n228), .Z(SUM[23]) );
  ND2P U104 ( .A(n183), .B(n184), .Z(n179) );
  ND2P U105 ( .A(n185), .B(n186), .Z(n178) );
  ND2P U106 ( .A(n74), .B(n73), .Z(n69) );
  AN2 U107 ( .A(n146), .B(n147), .Z(n35) );
  AN2 U108 ( .A(n1), .B(n10), .Z(n37) );
  IV U109 ( .A(B[31]), .Z(n137) );
  OR2P U110 ( .A(B[34]), .B(A[34]), .Z(n73) );
  IVA U111 ( .A(B[33]), .Z(n82) );
  IVA U112 ( .A(A[33]), .Z(n83) );
  AO3P U113 ( .A(n209), .B(n210), .C(n211), .D(n212), .Z(n103) );
  IVA U114 ( .A(B[27]), .Z(n185) );
  ND2P U115 ( .A(n257), .B(n44), .Z(n256) );
  EOP U116 ( .A(n45), .B(n46), .Z(SUM[37]) );
  EO U117 ( .A(n29), .B(n206), .Z(SUM[24]) );
  NR2 U118 ( .A(n205), .B(n173), .Z(n206) );
  ND2 U119 ( .A(n156), .B(n157), .Z(n154) );
  AO3 U120 ( .A(n112), .B(n113), .C(n114), .D(n115), .Z(n110) );
  AO3 U121 ( .A(n47), .B(n61), .C(n54), .D(n62), .Z(n57) );
  ND2 U122 ( .A(n55), .B(n56), .Z(n61) );
  ND2 U123 ( .A(n52), .B(n56), .Z(n62) );
  AO7 U124 ( .A(n47), .B(n84), .C(n68), .Z(n81) );
  AO7 U125 ( .A(n47), .B(n77), .C(n78), .Z(n76) );
  ND2 U126 ( .A(n75), .B(n74), .Z(n77) );
  AO6 U127 ( .A(n79), .B(n74), .C(n72), .Z(n78) );
  ND2 U128 ( .A(n114), .B(n111), .Z(n33) );
  ND2 U129 ( .A(n10), .B(n193), .Z(n204) );
  ND2 U130 ( .A(n7), .B(n116), .Z(n34) );
  NR2 U131 ( .A(n144), .B(n117), .Z(n164) );
  ND2 U132 ( .A(n176), .B(n108), .Z(n188) );
  ND2 U133 ( .A(n198), .B(n193), .Z(n194) );
  AO3 U134 ( .A(n199), .B(n200), .C(n10), .D(n192), .Z(n198) );
  NR2 U135 ( .A(n150), .B(n112), .Z(n149) );
  ND2 U136 ( .A(n151), .B(n152), .Z(n148) );
  ND2 U137 ( .A(n134), .B(n135), .Z(n118) );
  ND2 U138 ( .A(n134), .B(n135), .Z(n159) );
  AO7 U139 ( .A(n248), .B(n17), .C(n239), .Z(n246) );
  ND2 U140 ( .A(n218), .B(n93), .Z(n156) );
  IVA U141 ( .A(A[36]), .Z(n60) );
  NR2 U142 ( .A(n117), .B(n6), .Z(n162) );
  ND2 U143 ( .A(n234), .B(n235), .Z(n230) );
  ND2 U144 ( .A(n242), .B(n243), .Z(n234) );
  ND3 U145 ( .A(n201), .B(n157), .C(n156), .Z(n200) );
  ND2 U146 ( .A(n143), .B(n115), .Z(n142) );
  ND2 U147 ( .A(n35), .B(n144), .Z(n143) );
  ND2 U148 ( .A(n53), .B(n54), .Z(n50) );
  ND2 U149 ( .A(n104), .B(n213), .Z(n228) );
  ND2 U150 ( .A(n14), .B(n229), .Z(n227) );
  ND2 U151 ( .A(n230), .B(n31), .Z(n229) );
  ND2 U152 ( .A(n68), .B(n75), .Z(n36) );
  EO U153 ( .A(n230), .B(n231), .Z(SUM[22]) );
  NR2 U154 ( .A(n232), .B(n233), .Z(n231) );
  ND2 U155 ( .A(B[36]), .B(A[36]), .Z(n53) );
  ND4 U156 ( .A(B[12]), .B(n43), .C(n20), .D(n254), .Z(n135) );
  ND2 U157 ( .A(n134), .B(n135), .Z(n207) );
  ND2 U158 ( .A(B[20]), .B(A[20]), .Z(n210) );
  IVA U159 ( .A(B[35]), .Z(n65) );
  IVA U160 ( .A(A[35]), .Z(n66) );
  IVA U161 ( .A(B[32]), .Z(n86) );
  IVP U162 ( .A(A[32]), .Z(n87) );
  ND2 U163 ( .A(B[30]), .B(A[30]), .Z(n115) );
  ND2 U164 ( .A(B[20]), .B(A[20]), .Z(n239) );
  ND2 U165 ( .A(B[35]), .B(A[35]), .Z(n54) );
  ND4 U166 ( .A(n135), .B(n134), .C(n2), .D(n30), .Z(n243) );
  OR2 U167 ( .A(B[15]), .B(A[15]), .Z(n131) );
  ND2 U168 ( .A(B[29]), .B(n16), .Z(n113) );
  OR2 U169 ( .A(B[13]), .B(A[13]), .Z(n255) );
  ND2 U170 ( .A(B[23]), .B(A[23]), .Z(n213) );
  ND2 U171 ( .A(B[34]), .B(A[34]), .Z(n71) );
  ND2 U172 ( .A(B[16]), .B(n41), .Z(n250) );
  IV U173 ( .A(A[22]), .Z(n225) );
  IV U174 ( .A(B[22]), .Z(n224) );
  IVP U175 ( .A(A[19]), .Z(n267) );
  IV U176 ( .A(B[18]), .Z(n268) );
  IV U177 ( .A(B[25]), .Z(n183) );
  IVP U178 ( .A(A[27]), .Z(n186) );
  ND2 U179 ( .A(B[28]), .B(n11), .Z(n116) );
  ND2 U180 ( .A(B[24]), .B(A[24]), .Z(n201) );
  ND2 U181 ( .A(B[26]), .B(A[26]), .Z(n177) );
  ND2 U182 ( .A(B[27]), .B(A[27]), .Z(n176) );
  ND2 U183 ( .A(B[21]), .B(A[21]), .Z(n240) );
  ND2 U184 ( .A(n53), .B(n51), .Z(n58) );
  ENP U185 ( .A(n81), .B(n38), .Z(SUM[33]) );
  ND2 U186 ( .A(n80), .B(n74), .Z(n38) );
  ND2 U187 ( .A(n3), .B(n126), .Z(n155) );
  IV U188 ( .A(n23), .Z(n199) );
  ND2 U189 ( .A(n103), .B(n104), .Z(n157) );
  NR2 U190 ( .A(n19), .B(n98), .Z(n92) );
  NR2 U191 ( .A(n95), .B(n98), .Z(n218) );
  ND2 U192 ( .A(n106), .B(n108), .Z(n166) );
  ND2 U193 ( .A(n106), .B(n108), .Z(n169) );
  NR2 U194 ( .A(n123), .B(n32), .Z(n120) );
  AN2 U195 ( .A(n35), .B(n7), .Z(n140) );
  ND2 U196 ( .A(n141), .B(n7), .Z(n165) );
  AO7 U197 ( .A(n21), .B(n138), .C(n139), .Z(n136) );
  AO7 U198 ( .A(n21), .B(n155), .C(n165), .Z(n163) );
  AO7 U199 ( .A(n21), .B(n25), .C(n169), .Z(n167) );
  AO7 U200 ( .A(n205), .B(n21), .C(n201), .Z(n203) );
  ENP U201 ( .A(n76), .B(n39), .Z(SUM[34]) );
  ND2 U202 ( .A(n73), .B(n71), .Z(n39) );
  ND2 U203 ( .A(n54), .B(n56), .Z(n40) );
  OR2P U204 ( .A(A[20]), .B(B[20]), .Z(n220) );
  NR2 U205 ( .A(n241), .B(n238), .Z(n236) );
  NR2 U206 ( .A(n95), .B(n96), .Z(n94) );
  IVA U207 ( .A(B[19]), .Z(n266) );
  IVA U208 ( .A(B[26]), .Z(n196) );
  ND2 U209 ( .A(n191), .B(n5), .Z(n187) );
  ND2 U210 ( .A(n173), .B(n37), .Z(n189) );
  ND2 U211 ( .A(n172), .B(n37), .Z(n190) );
  ND3 U212 ( .A(n37), .B(n192), .C(n29), .Z(n191) );
  AO7 U213 ( .A(A[17]), .B(B[17]), .C(n253), .Z(n249) );
  ND3 U214 ( .A(A[17]), .B(B[17]), .C(n253), .Z(n252) );
  AO2 U215 ( .A(B[19]), .B(A[19]), .C(B[18]), .D(A[18]), .Z(n251) );
  IV U216 ( .A(A[30]), .Z(n128) );
  IVA U217 ( .A(B[30]), .Z(n127) );
  AN2P U218 ( .A(n99), .B(n100), .Z(n90) );
  ND2 U219 ( .A(B[31]), .B(n26), .Z(n114) );
  IV U220 ( .A(A[17]), .Z(n271) );
  AO2 U221 ( .A(B[14]), .B(A[14]), .C(B[15]), .D(A[15]), .Z(n132) );
  ND2 U222 ( .A(n240), .B(n15), .Z(n247) );
  IVA U223 ( .A(B[24]), .Z(n181) );
  ND2 U224 ( .A(n105), .B(n106), .Z(n99) );
  AO7 U225 ( .A(n109), .B(n110), .C(n111), .Z(n89) );
  AO6 U226 ( .A(n9), .B(n243), .C(n93), .Z(n248) );
  AO3 U227 ( .A(n159), .B(n208), .C(n161), .D(n8), .Z(n158) );
  OR2P U228 ( .A(A[25]), .B(B[25]), .Z(n174) );
  NR2 U229 ( .A(n238), .B(n13), .Z(n242) );
  ND2 U230 ( .A(n2), .B(n133), .Z(n160) );
  ND2 U231 ( .A(n2), .B(n30), .Z(n119) );
  ND3 U232 ( .A(A[13]), .B(B[13]), .C(n254), .Z(n134) );
  IVA U233 ( .A(B[28]), .Z(n168) );
  IV U234 ( .A(A[14]), .Z(n259) );
  ND2 U235 ( .A(n4), .B(n55), .Z(n48) );
  ENP U236 ( .A(n57), .B(n58), .Z(SUM[36]) );
  AO3P U237 ( .A(n68), .B(n69), .C(n70), .D(n71), .Z(n52) );
  ND2P U238 ( .A(n72), .B(n73), .Z(n70) );
  IVA U239 ( .A(n80), .Z(n72) );
  IVA U240 ( .A(n68), .Z(n79) );
  ND2P U241 ( .A(n82), .B(n83), .Z(n74) );
  IVA U242 ( .A(n75), .Z(n84) );
  ND4P U243 ( .A(n88), .B(n89), .C(n90), .D(n91), .Z(n85) );
  IVA U244 ( .A(n32), .Z(n102) );
  IVA U245 ( .A(n108), .Z(n107) );
  ND4P U246 ( .A(n28), .B(n125), .C(n126), .D(n111), .Z(n96) );
  ND2P U247 ( .A(n129), .B(n130), .Z(n124) );
  IVA U248 ( .A(n131), .Z(n123) );
  ND2P U249 ( .A(n137), .B(n27), .Z(n111) );
  ND2 U250 ( .A(n35), .B(n145), .Z(n138) );
  IVA U251 ( .A(n147), .Z(n112) );
  OR2 U252 ( .A(A[30]), .B(B[30]), .Z(n147) );
  IVA U253 ( .A(n115), .Z(n150) );
  IVA U254 ( .A(n155), .Z(n145) );
  IVA U255 ( .A(n158), .Z(n153) );
  IVA U256 ( .A(n146), .Z(n117) );
  IVA U257 ( .A(n113), .Z(n144) );
  ND2P U258 ( .A(n168), .B(n12), .Z(n126) );
  AN2P U259 ( .A(B[24]), .B(A[24]), .Z(n173) );
  AN2P U260 ( .A(n176), .B(n177), .Z(n170) );
  ND4P U261 ( .A(n178), .B(n179), .C(n180), .D(n175), .Z(n97) );
  ND2P U262 ( .A(n181), .B(n182), .Z(n180) );
  OR2 U263 ( .A(A[27]), .B(B[27]), .Z(n108) );
  AN2P U264 ( .A(n1), .B(n177), .Z(n195) );
  ND2P U265 ( .A(n196), .B(n197), .Z(n175) );
  ND2P U266 ( .A(B[25]), .B(A[25]), .Z(n193) );
  IVA U267 ( .A(n192), .Z(n205) );
  OR2 U268 ( .A(A[24]), .B(B[24]), .Z(n192) );
  IVA U269 ( .A(n98), .Z(n161) );
  ND3P U270 ( .A(n219), .B(n220), .C(n221), .Z(n98) );
  NR2P U271 ( .A(n222), .B(n223), .Z(n221) );
  IVA U272 ( .A(n226), .Z(n95) );
  OR2 U273 ( .A(A[23]), .B(B[23]), .Z(n104) );
  AO7P U274 ( .A(n244), .B(n18), .C(n15), .Z(n238) );
  IVA U275 ( .A(n239), .Z(n244) );
  ND2P U276 ( .A(n220), .B(n226), .Z(n245) );
  OR2 U277 ( .A(A[19]), .B(B[19]), .Z(n226) );
  AO3P U278 ( .A(n249), .B(n250), .C(n251), .D(n252), .Z(n93) );
  OR2 U279 ( .A(A[18]), .B(B[18]), .Z(n253) );
  ND2P U280 ( .A(n258), .B(n259), .Z(n254) );
  ND4P U281 ( .A(n261), .B(n262), .C(n263), .D(n264), .Z(n122) );
  ND2P U282 ( .A(n266), .B(n267), .Z(n263) );
endmodule


module SQRT_POLY_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [11:0] A;
  input [30:0] B;
  output [42:0] PRODUCT;
  input TC;
  wire   \ab[11][30] , \ab[11][29] , \ab[11][28] , \ab[11][27] , \ab[11][26] ,
         \ab[11][25] , \ab[11][24] , \ab[11][23] , \ab[11][22] , \ab[11][21] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][30] , \ab[10][29] , \ab[10][28] , \ab[10][27] ,
         \ab[10][26] , \ab[10][25] , \ab[10][24] , \ab[10][23] , \ab[10][22] ,
         \ab[10][21] , \ab[10][20] , \ab[10][19] , \ab[10][18] , \ab[10][17] ,
         \ab[10][16] , \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] ,
         \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] ,
         \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] ,
         \ab[10][1] , \ab[10][0] , \ab[9][30] , \ab[9][29] , \ab[9][28] ,
         \ab[9][27] , \ab[9][26] , \ab[9][25] , \ab[9][24] , \ab[9][23] ,
         \ab[9][22] , \ab[9][21] , \ab[9][20] , \ab[9][19] , \ab[9][18] ,
         \ab[9][17] , \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] ,
         \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] ,
         \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] ,
         \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][30] , \ab[8][29] ,
         \ab[8][28] , \ab[8][27] , \ab[8][26] , \ab[8][25] , \ab[8][24] ,
         \ab[8][23] , \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] ,
         \ab[8][18] , \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][30] ,
         \ab[7][29] , \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][30] , \ab[6][29] , \ab[6][28] , \ab[6][27] , \ab[6][26] ,
         \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] , \ab[6][21] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] ,
         \ab[5][26] , \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] ,
         \ab[5][21] , \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] ,
         \ab[5][16] , \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] ,
         \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] ,
         \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] ,
         \ab[5][1] , \ab[5][0] , \ab[4][30] , \ab[4][29] , \ab[4][28] ,
         \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] , \ab[4][23] ,
         \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][30] , \ab[3][29] ,
         \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] , \ab[3][24] ,
         \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] ,
         \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][30] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] , \ab[1][26] ,
         \ab[1][25] , \ab[1][24] , \ab[1][23] , \ab[1][22] , \ab[1][21] ,
         \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[0][30] , \ab[0][29] ,
         \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] ,
         \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] ,
         \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][23] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][29] , \CARRYB[10][28] , \CARRYB[10][27] ,
         \CARRYB[10][26] , \CARRYB[10][25] , \CARRYB[10][24] ,
         \CARRYB[10][23] , \CARRYB[10][22] , \CARRYB[10][21] ,
         \CARRYB[10][20] , \CARRYB[10][19] , \CARRYB[10][18] ,
         \CARRYB[10][17] , \CARRYB[10][16] , \CARRYB[10][15] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][29] , \CARRYB[9][28] , \CARRYB[9][27] , \CARRYB[9][26] ,
         \CARRYB[9][25] , \CARRYB[9][24] , \CARRYB[9][23] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][29] , \CARRYB[8][28] ,
         \CARRYB[8][27] , \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] ,
         \CARRYB[8][23] , \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] ,
         \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] ,
         \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] ,
         \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] ,
         \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] ,
         \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][29] , \CARRYB[6][28] ,
         \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] ,
         \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] ,
         \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] ,
         \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][29] , \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][29] , \CARRYB[4][28] ,
         \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] ,
         \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] ,
         \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] ,
         \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][29] , \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][29] , \CARRYB[2][28] ,
         \CARRYB[2][27] , \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] ,
         \CARRYB[2][23] , \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] ,
         \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] ,
         \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[1][29] , \CARRYB[1][28] , \CARRYB[1][27] , \CARRYB[1][26] ,
         \CARRYB[1][25] , \CARRYB[1][24] , \CARRYB[1][23] , \CARRYB[1][22] ,
         \CARRYB[1][21] , \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] ,
         \CARRYB[1][17] , \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] ,
         \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] ,
         \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] ,
         \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] ,
         \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[11][29] , \SUMB[11][28] ,
         \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] ,
         \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[11][0] ,
         \SUMB[10][29] , \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] ,
         \SUMB[10][25] , \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] ,
         \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] ,
         \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] ,
         \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] ,
         \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] ,
         \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] ,
         \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] ,
         \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] , \SUMB[8][26] ,
         \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] , \SUMB[8][22] ,
         \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] ,
         \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][29] ,
         \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] , \SUMB[7][25] ,
         \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] , \SUMB[7][21] ,
         \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] , \SUMB[7][17] ,
         \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] ,
         \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] ,
         \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][29] ,
         \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] , \SUMB[6][25] ,
         \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] , \SUMB[6][21] ,
         \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] ,
         \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] ,
         \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] ,
         \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][29] ,
         \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] , \SUMB[4][25] ,
         \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] , \SUMB[4][21] ,
         \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] , \SUMB[4][17] ,
         \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] ,
         \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] ,
         \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][29] ,
         \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] , \SUMB[3][25] ,
         \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] , \SUMB[3][21] ,
         \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] , \SUMB[3][17] ,
         \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][29] ,
         \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] , \SUMB[2][25] ,
         \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] , \SUMB[2][21] ,
         \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] , \SUMB[2][17] ,
         \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] ,
         \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] ,
         \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][29] ,
         \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] , \SUMB[1][25] ,
         \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] , \SUMB[1][21] ,
         \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] , \SUMB[1][17] ,
         \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] , \SUMB[1][13] ,
         \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] , \SUMB[1][9] ,
         \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[39] , \A1[38] ,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] ,
         \A1[1] , \A1[0] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] ,
         \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , \A2[29] ,
         \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] ,
         \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] ,
         \A2[14] , \A2[13] , \A2[12] , \A2[11] , n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  FA1AP S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  SQRT_POLY_DW01_add_2 FS_1 ( .A({1'b0, \A1[39] , \A1[38] , \A1[37] , \A1[36] , 
        \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , 
        \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , 
        \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \SUMB[11][0] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , 
        \A1[0] }), .B({\A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , 
        \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , \A2[29] , 
        \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] , 
        \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , 
        \A2[14] , \A2[13] , \A2[12] , \A2[11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, PRODUCT[39:23], SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}) );
  FA1P S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1P S2_7_10 ( .A(\CARRYB[6][10] ), .B(\ab[7][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1P S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1P S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1P S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1P S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1P S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1P S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1P S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1P S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1A S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1P S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1P S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1P S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1P S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1P S4_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(
        \CARRYB[11][0] ), .S(\SUMB[11][0] ) );
  FA1P S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1P S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1P S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1P S4_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(
        \CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1P S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1P S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1P S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA1P S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA1P S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1P S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1AP S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1P S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S4_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1P S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1P S2_5_14 ( .A(\CARRYB[4][14] ), .B(\ab[5][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1P S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1P S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1P S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1AP S4_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1AP S4_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(
        \CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_4_15 ( .A(\CARRYB[3][15] ), .B(\ab[4][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA1A S2_10_15 ( .A(\CARRYB[9][15] ), .B(\ab[10][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1AP S4_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(
        \CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S5_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\ab[10][30] ), .CO(
        \CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1A S3_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\ab[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1A S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S3_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\ab[8][30] ), .CO(
        \CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1A S3_2_29 ( .A(\ab[2][29] ), .B(\CARRYB[1][29] ), .CI(\ab[1][30] ), .CO(
        \CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1A S4_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1A S2_2_27 ( .A(\ab[2][27] ), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1A S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1AP S4_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1A S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1A S3_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\ab[7][30] ), .CO(
        \CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1A S3_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\ab[2][30] ), .CO(
        \CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1A S3_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\ab[5][30] ), .CO(
        \CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA1A S3_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\ab[3][30] ), .CO(
        \CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1A S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA1A S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA1A S2_2_28 ( .A(\ab[2][28] ), .B(\CARRYB[1][28] ), .CI(\SUMB[1][29] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FA1A S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA1A S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA1A S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA1A S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1A S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1A S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1 S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA1AP S4_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1P S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1 S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA1 S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1P S3_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\ab[4][30] ), .CO(
        \CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA1AP S4_15 ( .A(\CARRYB[10][15] ), .B(\ab[11][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1P S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1AP S2_2_10 ( .A(\CARRYB[1][10] ), .B(\ab[2][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1A S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA1 S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), .CO(
        \CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA1A S3_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\ab[6][30] ), .CO(
        \CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1A S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1 S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), .CO(
        \CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), .CO(
        \CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA1P S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1P S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1A S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA1AP S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1AP S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1P S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1 S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), .CO(
        \CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1A S2_10_21 ( .A(\CARRYB[9][21] ), .B(\ab[10][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1P S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1P S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1P S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1 S2_10_20 ( .A(\SUMB[9][21] ), .B(\CARRYB[9][20] ), .CI(\ab[10][20] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1P S2_5_15 ( .A(\CARRYB[4][15] ), .B(\ab[5][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_10_13 ( .A(\CARRYB[9][13] ), .B(\ab[10][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1P S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1P S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1P S2_2_25 ( .A(\ab[2][25] ), .B(\CARRYB[1][25] ), .CI(\SUMB[1][26] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1P S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA1AP S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1AP S4_21 ( .A(\CARRYB[10][21] ), .B(\ab[11][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA1A S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1P S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1P S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1 S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), .CO(
        \CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA1AP S2_5_17 ( .A(\CARRYB[4][17] ), .B(\ab[5][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1AP S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA1P S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1AP S2_8_11 ( .A(\CARRYB[7][11] ), .B(\ab[8][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_2_13 ( .A(\CARRYB[1][13] ), .B(\ab[2][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1AP S4_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1P S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1P S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1AP S2_5_12 ( .A(\CARRYB[4][12] ), .B(\ab[5][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1P S2_6_12 ( .A(\CARRYB[5][12] ), .B(\ab[6][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1P S4_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1P S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA1P S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1AP S4_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1P S2_6_20 ( .A(\CARRYB[5][20] ), .B(\ab[6][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1P S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1P S2_2_9 ( .A(\SUMB[1][10] ), .B(\CARRYB[1][9] ), .CI(\ab[2][9] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), .CO(
        \CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), .CO(
        \CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1P S2_2_17 ( .A(\CARRYB[1][17] ), .B(\ab[2][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1P S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1AP S4_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1AP S4_13 ( .A(\CARRYB[10][13] ), .B(\ab[11][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1P S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1P S2_2_20 ( .A(\SUMB[1][21] ), .B(\CARRYB[1][20] ), .CI(\ab[2][20] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1P S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1AP S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1P S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1P S2_3_17 ( .A(\CARRYB[2][17] ), .B(\ab[3][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1 S2_3_15 ( .A(\CARRYB[2][15] ), .B(\ab[3][15] ), .CI(\SUMB[2][16] ), .CO(
        \CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1AP S4_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1P S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1P S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1AP S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1P S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA1A S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1P S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), .CO(
        \CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1P S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1P S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1P S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1P S2_6_17 ( .A(\CARRYB[5][17] ), .B(\ab[6][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1P S4_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(
        \CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1P S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1A S4_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1P S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1AP S2_6_15 ( .A(\CARRYB[5][15] ), .B(\ab[6][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1AP S4_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1P S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), .CO(
        \CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA1P S2_7_14 ( .A(\CARRYB[6][14] ), .B(\ab[7][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1P S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_9 ( .A(\CARRYB[5][9] ), .B(\ab[6][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), .CO(
        \CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1P S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1P S4_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(
        \CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1 S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1P S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1 S2_7_4 ( .A(\CARRYB[6][4] ), .B(\ab[7][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1P S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA1P S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1P S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1AP S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_3_9 ( .A(\CARRYB[2][9] ), .B(\ab[3][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), .CO(
        \CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA1AP S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1AP S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), .CO(
        \CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1AP S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1AP S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1P S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA1A S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S4_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(
        \CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1 S2_10_17 ( .A(\CARRYB[9][17] ), .B(\ab[10][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), .CO(
        \CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S4_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1A S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1A S4_3 ( .A(\CARRYB[10][3] ), .B(\ab[11][3] ), .CI(\SUMB[10][4] ), .CO(
        \CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1A S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA1A S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA1AP S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA1P S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1P S4_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(
        \CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1AP S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1AP S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1AP S2_2_16 ( .A(\CARRYB[1][16] ), .B(\ab[2][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1A S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), .CO(
        \CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S4_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1AP S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1AP S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1AP S2_8_16 ( .A(\CARRYB[7][16] ), .B(\ab[8][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1 S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1AP S2_8_14 ( .A(\CARRYB[7][14] ), .B(\ab[8][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), .CO(
        \CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  IVDAP U2 ( .A(n237), .Y(n139), .Z(n141) );
  EO3 U3 ( .A(\CARRYB[8][21] ), .B(\ab[9][21] ), .C(\SUMB[8][22] ), .Z(
        \SUMB[9][21] ) );
  EO3P U4 ( .A(\CARRYB[6][9] ), .B(\ab[7][9] ), .C(\SUMB[6][10] ), .Z(
        \SUMB[7][9] ) );
  ND2 U5 ( .A(\CARRYB[6][9] ), .B(\SUMB[6][10] ), .Z(n3) );
  ND2 U6 ( .A(\CARRYB[6][9] ), .B(\ab[7][9] ), .Z(n4) );
  ND2 U7 ( .A(\SUMB[6][10] ), .B(\ab[7][9] ), .Z(n5) );
  ND3 U8 ( .A(n3), .B(n4), .C(n5), .Z(\CARRYB[7][9] ) );
  EO U9 ( .A(\CARRYB[7][9] ), .B(\ab[8][9] ), .Z(n131) );
  EO U10 ( .A(\SUMB[9][12] ), .B(\ab[10][11] ), .Z(n6) );
  EO U11 ( .A(\CARRYB[9][11] ), .B(n6), .Z(\SUMB[10][11] ) );
  ND2 U12 ( .A(\CARRYB[9][11] ), .B(\SUMB[9][12] ), .Z(n7) );
  ND2 U13 ( .A(\CARRYB[9][11] ), .B(\ab[10][11] ), .Z(n8) );
  ND2 U14 ( .A(\SUMB[9][12] ), .B(\ab[10][11] ), .Z(n9) );
  ND3 U15 ( .A(n7), .B(n8), .C(n9), .Z(\CARRYB[10][11] ) );
  EOP U16 ( .A(\SUMB[3][24] ), .B(\ab[4][23] ), .Z(n10) );
  EO U17 ( .A(\CARRYB[3][23] ), .B(n10), .Z(\SUMB[4][23] ) );
  ND2 U18 ( .A(\CARRYB[3][23] ), .B(\SUMB[3][24] ), .Z(n11) );
  ND2 U19 ( .A(\CARRYB[3][23] ), .B(\ab[4][23] ), .Z(n12) );
  ND2 U20 ( .A(\SUMB[3][24] ), .B(\ab[4][23] ), .Z(n13) );
  ND3 U21 ( .A(n11), .B(n12), .C(n13), .Z(\CARRYB[4][23] ) );
  EO U22 ( .A(\SUMB[5][28] ), .B(\ab[6][27] ), .Z(n14) );
  EO U23 ( .A(\CARRYB[5][27] ), .B(n14), .Z(\SUMB[6][27] ) );
  ND2 U24 ( .A(\CARRYB[5][27] ), .B(\SUMB[5][28] ), .Z(n15) );
  ND2 U25 ( .A(\CARRYB[5][27] ), .B(\ab[6][27] ), .Z(n16) );
  ND2 U26 ( .A(\SUMB[5][28] ), .B(\ab[6][27] ), .Z(n17) );
  ND3 U27 ( .A(n15), .B(n16), .C(n17), .Z(\CARRYB[6][27] ) );
  ND2 U28 ( .A(\CARRYB[3][17] ), .B(n19), .Z(n20) );
  ND2 U29 ( .A(n18), .B(\ab[4][17] ), .Z(n21) );
  ND2P U30 ( .A(n20), .B(n21), .Z(n102) );
  IVA U31 ( .A(\CARRYB[3][17] ), .Z(n18) );
  IVP U32 ( .A(\ab[4][17] ), .Z(n19) );
  EOP U33 ( .A(\SUMB[3][18] ), .B(n102), .Z(\SUMB[4][17] ) );
  EO U34 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .Z(n22) );
  EO U35 ( .A(\SUMB[6][6] ), .B(n22), .Z(\SUMB[7][5] ) );
  ND2 U36 ( .A(\SUMB[6][6] ), .B(\CARRYB[6][5] ), .Z(n23) );
  ND2 U37 ( .A(\SUMB[6][6] ), .B(\ab[7][5] ), .Z(n24) );
  ND2 U38 ( .A(\CARRYB[6][5] ), .B(\ab[7][5] ), .Z(n25) );
  ND3 U39 ( .A(n23), .B(n24), .C(n25), .Z(\CARRYB[7][5] ) );
  EO U40 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .Z(n146) );
  ND2 U41 ( .A(\SUMB[1][22] ), .B(n27), .Z(n28) );
  ND2 U42 ( .A(n26), .B(n106), .Z(n29) );
  ND2P U43 ( .A(n28), .B(n29), .Z(\SUMB[2][21] ) );
  IVDA U44 ( .A(\SUMB[1][22] ), .Y(n26) );
  IV U45 ( .A(n106), .Z(n27) );
  EO3P U46 ( .A(\CARRYB[2][16] ), .B(\ab[3][16] ), .C(\SUMB[2][17] ), .Z(
        \SUMB[3][16] ) );
  ND2 U47 ( .A(\CARRYB[2][16] ), .B(\SUMB[2][17] ), .Z(n30) );
  ND2 U48 ( .A(\CARRYB[2][16] ), .B(\ab[3][16] ), .Z(n31) );
  ND2 U49 ( .A(\SUMB[2][17] ), .B(\ab[3][16] ), .Z(n32) );
  ND3P U50 ( .A(n30), .B(n31), .C(n32), .Z(\CARRYB[3][16] ) );
  EOP U51 ( .A(\CARRYB[9][5] ), .B(\ab[10][5] ), .Z(n33) );
  EOP U52 ( .A(\SUMB[9][6] ), .B(n33), .Z(\SUMB[10][5] ) );
  ND2 U53 ( .A(\SUMB[9][6] ), .B(\CARRYB[9][5] ), .Z(n34) );
  ND2 U54 ( .A(\SUMB[9][6] ), .B(\ab[10][5] ), .Z(n35) );
  ND2 U55 ( .A(\CARRYB[9][5] ), .B(\ab[10][5] ), .Z(n36) );
  ND3 U56 ( .A(n34), .B(n35), .C(n36), .Z(\CARRYB[10][5] ) );
  EO3P U57 ( .A(\SUMB[9][7] ), .B(\ab[10][6] ), .C(\CARRYB[9][6] ), .Z(
        \SUMB[10][6] ) );
  ND2 U58 ( .A(\SUMB[9][7] ), .B(\CARRYB[9][6] ), .Z(n37) );
  ND2 U59 ( .A(\SUMB[9][7] ), .B(\ab[10][6] ), .Z(n38) );
  ND2 U60 ( .A(\CARRYB[9][6] ), .B(\ab[10][6] ), .Z(n39) );
  ND3 U61 ( .A(n37), .B(n38), .C(n39), .Z(\CARRYB[10][6] ) );
  EO U62 ( .A(\SUMB[8][1] ), .B(\ab[9][0] ), .Z(n40) );
  EO U63 ( .A(\CARRYB[8][0] ), .B(n40), .Z(\A1[7] ) );
  ND2 U64 ( .A(\CARRYB[8][0] ), .B(\SUMB[8][1] ), .Z(n41) );
  ND2 U65 ( .A(\CARRYB[8][0] ), .B(\ab[9][0] ), .Z(n42) );
  ND2 U66 ( .A(\SUMB[8][1] ), .B(\ab[9][0] ), .Z(n43) );
  ND3 U67 ( .A(n41), .B(n42), .C(n43), .Z(\CARRYB[9][0] ) );
  EO3P U68 ( .A(\CARRYB[4][4] ), .B(\ab[5][4] ), .C(\SUMB[4][5] ), .Z(
        \SUMB[5][4] ) );
  ND2 U69 ( .A(\CARRYB[4][4] ), .B(\SUMB[4][5] ), .Z(n44) );
  ND2 U70 ( .A(\CARRYB[4][4] ), .B(\ab[5][4] ), .Z(n45) );
  ND2 U71 ( .A(\SUMB[4][5] ), .B(\ab[5][4] ), .Z(n46) );
  ND3 U72 ( .A(n44), .B(n45), .C(n46), .Z(\CARRYB[5][4] ) );
  ND3 U73 ( .A(n73), .B(n74), .C(n75), .Z(\CARRYB[4][4] ) );
  EOP U74 ( .A(\CARRYB[3][19] ), .B(\ab[4][19] ), .Z(n47) );
  EOP U75 ( .A(\SUMB[3][20] ), .B(n47), .Z(\SUMB[4][19] ) );
  ND2 U76 ( .A(\SUMB[3][20] ), .B(\CARRYB[3][19] ), .Z(n48) );
  ND2 U77 ( .A(\SUMB[3][20] ), .B(\ab[4][19] ), .Z(n49) );
  ND2 U78 ( .A(\CARRYB[3][19] ), .B(\ab[4][19] ), .Z(n50) );
  ND3 U79 ( .A(n48), .B(n49), .C(n50), .Z(\CARRYB[4][19] ) );
  ND3P U80 ( .A(n52), .B(n53), .C(n54), .Z(\CARRYB[3][19] ) );
  EO U81 ( .A(\CARRYB[2][19] ), .B(\ab[3][19] ), .Z(n51) );
  EO U82 ( .A(\SUMB[2][20] ), .B(n51), .Z(\SUMB[3][19] ) );
  ND2 U83 ( .A(\SUMB[2][20] ), .B(\CARRYB[2][19] ), .Z(n52) );
  ND2 U84 ( .A(\SUMB[2][20] ), .B(\ab[3][19] ), .Z(n53) );
  ND2 U85 ( .A(\CARRYB[2][19] ), .B(\ab[3][19] ), .Z(n54) );
  EOP U86 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A1[17] ) );
  EOP U87 ( .A(\SUMB[4][11] ), .B(n190), .Z(\SUMB[5][10] ) );
  EOP U88 ( .A(\SUMB[9][8] ), .B(n68), .Z(\SUMB[10][7] ) );
  AN2 U89 ( .A(n215), .B(B[8]), .Z(\ab[3][8] ) );
  ND3 U90 ( .A(n143), .B(n144), .C(n145), .Z(\CARRYB[2][8] ) );
  EOP U91 ( .A(\SUMB[8][6] ), .B(n179), .Z(\SUMB[9][5] ) );
  B3IP U92 ( .A(A[0]), .Z1(n57), .Z2(n58) );
  EO U93 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Z(\SUMB[1][27] ) );
  ND2 U94 ( .A(\CARRYB[8][3] ), .B(\ab[9][3] ), .Z(n137) );
  EO U95 ( .A(\CARRYB[8][5] ), .B(\ab[9][5] ), .Z(n179) );
  ND3 U96 ( .A(n169), .B(n170), .C(n171), .Z(\CARRYB[7][22] ) );
  EO U97 ( .A(\CARRYB[7][19] ), .B(\ab[8][19] ), .Z(n86) );
  EO U98 ( .A(\CARRYB[11][23] ), .B(\SUMB[11][24] ), .Z(\A1[33] ) );
  EO U99 ( .A(\CARRYB[11][24] ), .B(\SUMB[11][25] ), .Z(\A1[34] ) );
  EO U100 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Z(\SUMB[1][29] ) );
  EO U101 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Z(\SUMB[1][24] ) );
  ND2 U102 ( .A(\SUMB[1][9] ), .B(\ab[2][8] ), .Z(n144) );
  EO U103 ( .A(\CARRYB[1][15] ), .B(\ab[2][15] ), .Z(n94) );
  EO U104 ( .A(\SUMB[5][15] ), .B(n110), .Z(\SUMB[6][14] ) );
  EO U105 ( .A(\CARRYB[7][21] ), .B(\ab[8][21] ), .Z(n127) );
  EO U106 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U107 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U108 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U109 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U110 ( .A(\CARRYB[5][11] ), .B(\ab[6][11] ), .Z(n154) );
  ND3 U111 ( .A(n128), .B(n129), .C(n130), .Z(\CARRYB[8][21] ) );
  ND2 U112 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Z(n128) );
  ND2 U113 ( .A(\SUMB[7][22] ), .B(\ab[8][21] ), .Z(n129) );
  ND2 U114 ( .A(\CARRYB[8][21] ), .B(\ab[9][21] ), .Z(n209) );
  ND3 U115 ( .A(n172), .B(n173), .C(n174), .Z(\CARRYB[10][9] ) );
  ND2 U116 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .Z(n172) );
  ND2 U117 ( .A(\CARRYB[9][9] ), .B(\SUMB[9][10] ), .Z(n174) );
  ND3 U118 ( .A(n198), .B(n199), .C(n200), .Z(\CARRYB[9][22] ) );
  EO U119 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A1[12] ) );
  ND2 U120 ( .A(\SUMB[9][19] ), .B(\ab[10][18] ), .Z(n122) );
  EO U121 ( .A(\SUMB[9][19] ), .B(n120), .Z(\SUMB[10][18] ) );
  ND2 U122 ( .A(\SUMB[7][4] ), .B(\ab[8][3] ), .Z(n118) );
  EO U123 ( .A(\CARRYB[5][2] ), .B(n211), .Z(\SUMB[6][2] ) );
  EO U124 ( .A(\SUMB[7][4] ), .B(n116), .Z(\SUMB[8][3] ) );
  EO U125 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .Z(n116) );
  EO U126 ( .A(\SUMB[11][7] ), .B(\CARRYB[11][6] ), .Z(\A1[16] ) );
  IVDAP U127 ( .A(A[2]), .Y(n55), .Z(n56) );
  B2I U128 ( .A(A[4]), .Z2(n59) );
  IVDA U129 ( .A(B[28]), .Y(n60), .Z(n61) );
  B2I U130 ( .A(A[3]), .Z2(n215) );
  IVP U131 ( .A(n55), .Z(n188) );
  IVDA U132 ( .A(B[29]), .Y(n62), .Z(n63) );
  ND3 U133 ( .A(n212), .B(n213), .C(n214), .Z(\CARRYB[6][2] ) );
  ND3P U134 ( .A(n195), .B(n196), .C(n197), .Z(\CARRYB[9][5] ) );
  EO U135 ( .A(\CARRYB[9][18] ), .B(\ab[10][18] ), .Z(n120) );
  ND2 U136 ( .A(\SUMB[9][19] ), .B(\CARRYB[9][18] ), .Z(n121) );
  ND3 U137 ( .A(n121), .B(n122), .C(n123), .Z(\CARRYB[10][18] ) );
  EO U138 ( .A(\CARRYB[5][22] ), .B(\ab[6][22] ), .Z(n64) );
  EO U139 ( .A(\SUMB[5][23] ), .B(n64), .Z(\SUMB[6][22] ) );
  ND2 U140 ( .A(\SUMB[5][23] ), .B(\CARRYB[5][22] ), .Z(n65) );
  ND2 U141 ( .A(\SUMB[5][23] ), .B(\ab[6][22] ), .Z(n66) );
  ND2 U142 ( .A(\CARRYB[5][22] ), .B(\ab[6][22] ), .Z(n67) );
  ND3 U143 ( .A(n65), .B(n66), .C(n67), .Z(\CARRYB[6][22] ) );
  EO U144 ( .A(\CARRYB[6][22] ), .B(\ab[7][22] ), .Z(n168) );
  EO U145 ( .A(\CARRYB[9][7] ), .B(\ab[10][7] ), .Z(n68) );
  ND2 U146 ( .A(\SUMB[9][8] ), .B(\CARRYB[9][7] ), .Z(n69) );
  ND2 U147 ( .A(\SUMB[9][8] ), .B(\ab[10][7] ), .Z(n70) );
  ND2 U148 ( .A(\CARRYB[9][7] ), .B(\ab[10][7] ), .Z(n71) );
  ND3 U149 ( .A(n69), .B(n70), .C(n71), .Z(\CARRYB[10][7] ) );
  EO U150 ( .A(\CARRYB[3][4] ), .B(\ab[4][4] ), .Z(n72) );
  EO U151 ( .A(\SUMB[3][5] ), .B(n72), .Z(\SUMB[4][4] ) );
  ND2 U152 ( .A(\SUMB[3][5] ), .B(\CARRYB[3][4] ), .Z(n73) );
  ND2 U153 ( .A(\SUMB[3][5] ), .B(\ab[4][4] ), .Z(n74) );
  ND2 U154 ( .A(\CARRYB[3][4] ), .B(\ab[4][4] ), .Z(n75) );
  EO3 U155 ( .A(\CARRYB[2][5] ), .B(\ab[3][5] ), .C(\SUMB[2][6] ), .Z(
        \SUMB[3][5] ) );
  ND2 U156 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Z(n76) );
  ND2 U157 ( .A(\CARRYB[2][5] ), .B(\ab[3][5] ), .Z(n77) );
  ND2 U158 ( .A(\SUMB[2][6] ), .B(\ab[3][5] ), .Z(n78) );
  ND3 U159 ( .A(n76), .B(n77), .C(n78), .Z(\CARRYB[3][5] ) );
  EO U160 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  AN2P U161 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\CARRYB[1][26] ) );
  EO3P U162 ( .A(\SUMB[4][12] ), .B(\ab[5][11] ), .C(\CARRYB[4][11] ), .Z(
        \SUMB[5][11] ) );
  ND2 U163 ( .A(\SUMB[4][12] ), .B(\CARRYB[4][11] ), .Z(n79) );
  ND2 U164 ( .A(\SUMB[4][12] ), .B(\ab[5][11] ), .Z(n80) );
  ND2 U165 ( .A(\CARRYB[4][11] ), .B(\ab[5][11] ), .Z(n81) );
  ND3P U166 ( .A(n79), .B(n80), .C(n81), .Z(\CARRYB[5][11] ) );
  EO U167 ( .A(\CARRYB[3][12] ), .B(\ab[4][12] ), .Z(n82) );
  EOP U168 ( .A(\SUMB[3][13] ), .B(n82), .Z(\SUMB[4][12] ) );
  ND2 U169 ( .A(\SUMB[3][13] ), .B(\CARRYB[3][12] ), .Z(n83) );
  ND2 U170 ( .A(\SUMB[3][13] ), .B(\ab[4][12] ), .Z(n84) );
  ND2 U171 ( .A(\CARRYB[3][12] ), .B(\ab[4][12] ), .Z(n85) );
  ND3 U172 ( .A(n83), .B(n84), .C(n85), .Z(\CARRYB[4][12] ) );
  ND3 U173 ( .A(n132), .B(n133), .C(n134), .Z(\CARRYB[8][9] ) );
  AN2 U174 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  EO U175 ( .A(\SUMB[7][20] ), .B(n86), .Z(\SUMB[8][19] ) );
  ND2 U176 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Z(n87) );
  ND2 U177 ( .A(\SUMB[7][20] ), .B(\ab[8][19] ), .Z(n88) );
  ND2 U178 ( .A(\CARRYB[7][19] ), .B(\ab[8][19] ), .Z(n89) );
  ND3P U179 ( .A(n87), .B(n88), .C(n89), .Z(\CARRYB[8][19] ) );
  EOP U180 ( .A(\SUMB[3][10] ), .B(\ab[4][9] ), .Z(n90) );
  EOP U181 ( .A(\CARRYB[3][9] ), .B(n90), .Z(\SUMB[4][9] ) );
  ND2 U182 ( .A(\CARRYB[3][9] ), .B(\SUMB[3][10] ), .Z(n91) );
  ND2 U183 ( .A(\CARRYB[3][9] ), .B(\ab[4][9] ), .Z(n92) );
  ND2 U184 ( .A(\SUMB[3][10] ), .B(\ab[4][9] ), .Z(n93) );
  ND3P U185 ( .A(n91), .B(n92), .C(n93), .Z(\CARRYB[4][9] ) );
  ND3 U186 ( .A(n191), .B(n192), .C(n193), .Z(\CARRYB[5][10] ) );
  EOP U187 ( .A(\SUMB[1][16] ), .B(n94), .Z(\SUMB[2][15] ) );
  ND2 U188 ( .A(\SUMB[1][16] ), .B(\CARRYB[1][15] ), .Z(n95) );
  ND2 U189 ( .A(\SUMB[1][16] ), .B(\ab[2][15] ), .Z(n96) );
  ND2 U190 ( .A(\CARRYB[1][15] ), .B(\ab[2][15] ), .Z(n97) );
  ND3 U191 ( .A(n95), .B(n96), .C(n97), .Z(\CARRYB[2][15] ) );
  EO U192 ( .A(\ab[0][17] ), .B(n115), .Z(\SUMB[1][16] ) );
  AN2P U193 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  EOP U194 ( .A(\CARRYB[4][16] ), .B(\ab[5][16] ), .Z(n98) );
  EOP U195 ( .A(\SUMB[4][17] ), .B(n98), .Z(\SUMB[5][16] ) );
  ND2 U196 ( .A(\SUMB[4][17] ), .B(\CARRYB[4][16] ), .Z(n99) );
  ND2 U197 ( .A(\SUMB[4][17] ), .B(\ab[5][16] ), .Z(n100) );
  ND2 U198 ( .A(\CARRYB[4][16] ), .B(\ab[5][16] ), .Z(n101) );
  ND3 U199 ( .A(n99), .B(n100), .C(n101), .Z(\CARRYB[5][16] ) );
  ND2 U200 ( .A(\SUMB[3][18] ), .B(\CARRYB[3][17] ), .Z(n103) );
  ND2 U201 ( .A(\SUMB[3][18] ), .B(\ab[4][17] ), .Z(n104) );
  ND2 U202 ( .A(\CARRYB[3][17] ), .B(\ab[4][17] ), .Z(n105) );
  ND3 U203 ( .A(n103), .B(n104), .C(n105), .Z(\CARRYB[4][17] ) );
  AN2 U204 ( .A(n140), .B(B[4]), .Z(\ab[1][4] ) );
  EOP U205 ( .A(\CARRYB[1][21] ), .B(\ab[2][21] ), .Z(n106) );
  ND2 U206 ( .A(\SUMB[1][22] ), .B(\CARRYB[1][21] ), .Z(n107) );
  ND2 U207 ( .A(\SUMB[1][22] ), .B(\ab[2][21] ), .Z(n108) );
  ND2 U208 ( .A(\CARRYB[1][21] ), .B(\ab[2][21] ), .Z(n109) );
  ND3 U209 ( .A(n107), .B(n108), .C(n109), .Z(\CARRYB[2][21] ) );
  EOP U210 ( .A(\CARRYB[5][14] ), .B(\ab[6][14] ), .Z(n110) );
  ND2 U211 ( .A(\SUMB[5][15] ), .B(\CARRYB[5][14] ), .Z(n111) );
  ND2 U212 ( .A(\SUMB[5][15] ), .B(\ab[6][14] ), .Z(n112) );
  ND2 U213 ( .A(\CARRYB[5][14] ), .B(\ab[6][14] ), .Z(n113) );
  ND3P U214 ( .A(n111), .B(n112), .C(n113), .Z(\CARRYB[6][14] ) );
  ND3 U215 ( .A(n165), .B(n166), .C(n167), .Z(\CARRYB[3][4] ) );
  IVDA U216 ( .A(\SUMB[10][10] ), .Z(n114) );
  ND2 U217 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Z(n117) );
  AN2P U218 ( .A(n189), .B(B[16]), .Z(n115) );
  ND2P U219 ( .A(\CARRYB[5][11] ), .B(\ab[6][11] ), .Z(n157) );
  ND2 U220 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .Z(n119) );
  ND3P U221 ( .A(n117), .B(n118), .C(n119), .Z(\CARRYB[8][3] ) );
  ND2 U222 ( .A(\CARRYB[9][18] ), .B(\ab[10][18] ), .Z(n123) );
  EOP U223 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Z(\SUMB[1][21] ) );
  AN2P U224 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\CARRYB[1][19] ) );
  ND2 U225 ( .A(\CARRYB[4][16] ), .B(\SUMB[4][17] ), .Z(n124) );
  ND2 U226 ( .A(\CARRYB[4][16] ), .B(\ab[5][16] ), .Z(n125) );
  ND2 U227 ( .A(\SUMB[4][17] ), .B(\ab[5][16] ), .Z(n126) );
  ND3 U228 ( .A(n124), .B(n125), .C(n126), .Z(n138) );
  ND2 U229 ( .A(\SUMB[1][9] ), .B(\CARRYB[1][8] ), .Z(n143) );
  EO U230 ( .A(\SUMB[7][22] ), .B(n127), .Z(\SUMB[8][21] ) );
  ND2 U231 ( .A(\CARRYB[7][21] ), .B(\ab[8][21] ), .Z(n130) );
  AN2P U232 ( .A(n58), .B(B[20]), .Z(\ab[0][20] ) );
  EOP U233 ( .A(\SUMB[7][10] ), .B(n131), .Z(\SUMB[8][9] ) );
  ND2 U234 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Z(n132) );
  ND2 U235 ( .A(\SUMB[7][10] ), .B(\ab[8][9] ), .Z(n133) );
  ND2 U236 ( .A(\CARRYB[7][9] ), .B(\ab[8][9] ), .Z(n134) );
  EOP U237 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Z(\SUMB[1][22] ) );
  EOP U238 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\SUMB[1][19] ) );
  EO3P U239 ( .A(\SUMB[8][4] ), .B(\ab[9][3] ), .C(\CARRYB[8][3] ), .Z(
        \SUMB[9][3] ) );
  ND2 U240 ( .A(\SUMB[8][4] ), .B(\CARRYB[8][3] ), .Z(n135) );
  ND2 U241 ( .A(\SUMB[8][4] ), .B(\ab[9][3] ), .Z(n136) );
  ND3 U242 ( .A(n135), .B(n136), .C(n137), .Z(\CARRYB[9][3] ) );
  B4IP U243 ( .A(n235), .Z(n233) );
  AN2P U244 ( .A(n233), .B(B[8]), .Z(\ab[0][8] ) );
  IV U245 ( .A(n139), .Z(n140) );
  EOP U246 ( .A(\CARRYB[1][8] ), .B(\ab[2][8] ), .Z(n142) );
  EOP U247 ( .A(\SUMB[1][9] ), .B(n142), .Z(\SUMB[2][8] ) );
  ND2 U248 ( .A(\CARRYB[1][8] ), .B(\ab[2][8] ), .Z(n145) );
  EOP U249 ( .A(n146), .B(\SUMB[7][6] ), .Z(\SUMB[8][5] ) );
  ND2 U250 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Z(n147) );
  ND2 U251 ( .A(\SUMB[7][6] ), .B(\ab[8][5] ), .Z(n148) );
  ND2 U252 ( .A(\CARRYB[7][5] ), .B(\ab[8][5] ), .Z(n149) );
  ND3P U253 ( .A(n147), .B(n148), .C(n149), .Z(\CARRYB[8][5] ) );
  EOP U254 ( .A(\SUMB[9][17] ), .B(\ab[10][16] ), .Z(n150) );
  EOP U255 ( .A(\CARRYB[9][16] ), .B(n150), .Z(\SUMB[10][16] ) );
  ND2 U256 ( .A(\CARRYB[9][16] ), .B(\SUMB[9][17] ), .Z(n151) );
  ND2 U257 ( .A(\CARRYB[9][16] ), .B(\ab[10][16] ), .Z(n152) );
  ND2 U258 ( .A(\SUMB[9][17] ), .B(\ab[10][16] ), .Z(n153) );
  ND3P U259 ( .A(n151), .B(n152), .C(n153), .Z(\CARRYB[10][16] ) );
  IVA U260 ( .A(n55), .Z(n239) );
  AN2P U261 ( .A(n58), .B(B[16]), .Z(\ab[0][16] ) );
  AN2P U262 ( .A(n58), .B(B[18]), .Z(\ab[0][18] ) );
  AN2 U263 ( .A(n58), .B(B[12]), .Z(\ab[0][12] ) );
  AN2P U264 ( .A(n58), .B(B[19]), .Z(\ab[0][19] ) );
  IVAP U265 ( .A(n238), .Z(n189) );
  EOP U266 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\SUMB[1][10] ) );
  AN2P U267 ( .A(n233), .B(B[11]), .Z(\ab[0][11] ) );
  EOP U268 ( .A(\SUMB[5][12] ), .B(n154), .Z(\SUMB[6][11] ) );
  ND2P U269 ( .A(\SUMB[5][12] ), .B(\CARRYB[5][11] ), .Z(n155) );
  ND2P U270 ( .A(\SUMB[5][12] ), .B(\ab[6][11] ), .Z(n156) );
  ND3P U271 ( .A(n155), .B(n156), .C(n157), .Z(\CARRYB[6][11] ) );
  EOP U272 ( .A(\CARRYB[8][10] ), .B(\ab[9][10] ), .Z(n158) );
  EOP U273 ( .A(\SUMB[8][11] ), .B(n158), .Z(\SUMB[9][10] ) );
  ND2 U274 ( .A(\SUMB[8][11] ), .B(\CARRYB[8][10] ), .Z(n159) );
  ND2 U275 ( .A(\SUMB[8][11] ), .B(\ab[9][10] ), .Z(n160) );
  ND2 U276 ( .A(\CARRYB[8][10] ), .B(\ab[9][10] ), .Z(n161) );
  ND3 U277 ( .A(n159), .B(n160), .C(n161), .Z(\CARRYB[9][10] ) );
  IVA U278 ( .A(n238), .Z(n237) );
  AN2P U279 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\CARRYB[1][20] ) );
  EOP U280 ( .A(\CARRYB[11][16] ), .B(\SUMB[11][17] ), .Z(\A1[26] ) );
  EO U281 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO3P U282 ( .A(\SUMB[5][17] ), .B(\ab[6][16] ), .C(n138), .Z(\SUMB[6][16] )
         );
  ND2 U283 ( .A(\SUMB[5][17] ), .B(\CARRYB[5][16] ), .Z(n162) );
  ND2 U284 ( .A(\SUMB[5][17] ), .B(\ab[6][16] ), .Z(n163) );
  ND2 U285 ( .A(\CARRYB[5][16] ), .B(\ab[6][16] ), .Z(n164) );
  ND3 U286 ( .A(n162), .B(n163), .C(n164), .Z(\CARRYB[6][16] ) );
  EO U287 ( .A(\CARRYB[6][23] ), .B(n180), .Z(\SUMB[7][23] ) );
  EO3P U288 ( .A(\CARRYB[2][4] ), .B(\ab[3][4] ), .C(\SUMB[2][5] ), .Z(
        \SUMB[3][4] ) );
  ND2 U289 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Z(n165) );
  ND2 U290 ( .A(\CARRYB[2][4] ), .B(\ab[3][4] ), .Z(n166) );
  ND2 U291 ( .A(\SUMB[2][5] ), .B(\ab[3][4] ), .Z(n167) );
  AN2P U292 ( .A(n236), .B(n256), .Z(\ab[1][25] ) );
  EOP U293 ( .A(\SUMB[6][23] ), .B(n168), .Z(\SUMB[7][22] ) );
  ND2 U294 ( .A(\SUMB[6][23] ), .B(\CARRYB[6][22] ), .Z(n169) );
  ND2 U295 ( .A(\SUMB[6][23] ), .B(\ab[7][22] ), .Z(n170) );
  ND2 U296 ( .A(\CARRYB[6][22] ), .B(\ab[7][22] ), .Z(n171) );
  EO3 U297 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .C(\SUMB[9][10] ), .Z(
        \SUMB[10][9] ) );
  ND2 U298 ( .A(\ab[10][9] ), .B(\SUMB[9][10] ), .Z(n173) );
  EOP U299 ( .A(\SUMB[10][10] ), .B(\ab[11][9] ), .Z(n175) );
  EOP U300 ( .A(n175), .B(\CARRYB[10][9] ), .Z(\SUMB[11][9] ) );
  ND2 U301 ( .A(\ab[11][9] ), .B(n114), .Z(n176) );
  ND2 U302 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .Z(n177) );
  ND2 U303 ( .A(n114), .B(\CARRYB[10][9] ), .Z(n178) );
  ND3 U304 ( .A(n176), .B(n177), .C(n178), .Z(\CARRYB[11][9] ) );
  IVA U305 ( .A(n238), .Z(n236) );
  EOP U306 ( .A(\SUMB[6][24] ), .B(\ab[7][23] ), .Z(n180) );
  ND2P U307 ( .A(\CARRYB[6][23] ), .B(\SUMB[6][24] ), .Z(n181) );
  ND2P U308 ( .A(\CARRYB[6][23] ), .B(\ab[7][23] ), .Z(n182) );
  ND2 U309 ( .A(\SUMB[6][24] ), .B(\ab[7][23] ), .Z(n183) );
  ND3P U310 ( .A(n181), .B(n182), .C(n183), .Z(\CARRYB[7][23] ) );
  EOP U311 ( .A(\CARRYB[7][20] ), .B(\ab[8][20] ), .Z(n184) );
  EOP U312 ( .A(\SUMB[7][21] ), .B(n184), .Z(\SUMB[8][20] ) );
  ND2 U313 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Z(n185) );
  ND2 U314 ( .A(\SUMB[7][21] ), .B(\ab[8][20] ), .Z(n186) );
  ND2 U315 ( .A(\CARRYB[7][20] ), .B(\ab[8][20] ), .Z(n187) );
  ND3 U316 ( .A(n185), .B(n186), .C(n187), .Z(\CARRYB[8][20] ) );
  EOP U317 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A1[13] ) );
  EOP U318 ( .A(\CARRYB[4][10] ), .B(\ab[5][10] ), .Z(n190) );
  ND2 U319 ( .A(\SUMB[4][11] ), .B(\CARRYB[4][10] ), .Z(n191) );
  ND2 U320 ( .A(\SUMB[4][11] ), .B(\ab[5][10] ), .Z(n192) );
  ND2 U321 ( .A(\CARRYB[4][10] ), .B(\ab[5][10] ), .Z(n193) );
  IVP U322 ( .A(n57), .Z(n234) );
  ND2 U323 ( .A(\CARRYB[8][22] ), .B(n194), .Z(n198) );
  ND2 U324 ( .A(\CARRYB[8][22] ), .B(\ab[9][22] ), .Z(n199) );
  FA1A U325 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), .S(
        n194) );
  EO U326 ( .A(\SUMB[3][4] ), .B(\ab[4][3] ), .Z(n201) );
  EO U327 ( .A(\CARRYB[3][3] ), .B(n201), .Z(\SUMB[4][3] ) );
  IVAP U328 ( .A(A[1]), .Z(n238) );
  ND2 U329 ( .A(\CARRYB[8][5] ), .B(\SUMB[8][6] ), .Z(n195) );
  ND2 U330 ( .A(\CARRYB[8][5] ), .B(\ab[9][5] ), .Z(n196) );
  ND2 U331 ( .A(\SUMB[8][6] ), .B(\ab[9][5] ), .Z(n197) );
  EO3 U332 ( .A(\CARRYB[8][22] ), .B(\ab[9][22] ), .C(\SUMB[8][23] ), .Z(
        \SUMB[9][22] ) );
  ND2 U333 ( .A(n194), .B(\ab[9][22] ), .Z(n200) );
  EOP U334 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Z(\SUMB[1][26] ) );
  EO U335 ( .A(\SUMB[5][3] ), .B(\ab[6][2] ), .Z(n211) );
  ND2 U336 ( .A(\CARRYB[3][3] ), .B(\SUMB[3][4] ), .Z(n202) );
  ND2 U337 ( .A(\CARRYB[3][3] ), .B(\ab[4][3] ), .Z(n203) );
  ND2 U338 ( .A(\SUMB[3][4] ), .B(\ab[4][3] ), .Z(n204) );
  ND3P U339 ( .A(n202), .B(n203), .C(n204), .Z(\CARRYB[4][3] ) );
  EO3P U340 ( .A(\CARRYB[10][20] ), .B(\ab[11][20] ), .C(\SUMB[10][21] ), .Z(
        \SUMB[11][20] ) );
  ND2 U341 ( .A(\CARRYB[10][20] ), .B(\SUMB[10][21] ), .Z(n205) );
  ND2 U342 ( .A(\CARRYB[10][20] ), .B(\ab[11][20] ), .Z(n206) );
  ND2 U343 ( .A(\SUMB[10][21] ), .B(\ab[11][20] ), .Z(n207) );
  ND3 U344 ( .A(n205), .B(n206), .C(n207), .Z(\CARRYB[11][20] ) );
  IVP U345 ( .A(n232), .Z(n231) );
  IVP U346 ( .A(n259), .Z(n258) );
  IVP U347 ( .A(n257), .Z(n256) );
  EO U348 ( .A(\CARRYB[11][22] ), .B(\SUMB[11][23] ), .Z(\A1[32] ) );
  IVA U349 ( .A(n238), .Z(n217) );
  EOP U350 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\SUMB[1][18] ) );
  AN2P U351 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  ND2 U352 ( .A(\CARRYB[8][21] ), .B(\SUMB[8][22] ), .Z(n208) );
  ND2 U353 ( .A(\SUMB[8][22] ), .B(\ab[9][21] ), .Z(n210) );
  ND3 U354 ( .A(n208), .B(n209), .C(n210), .Z(\CARRYB[9][21] ) );
  ND2 U355 ( .A(\CARRYB[5][2] ), .B(\SUMB[5][3] ), .Z(n212) );
  ND2 U356 ( .A(\CARRYB[5][2] ), .B(\ab[6][2] ), .Z(n213) );
  ND2 U357 ( .A(\SUMB[5][3] ), .B(\ab[6][2] ), .Z(n214) );
  EOP U358 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A1[14] ) );
  EOP U359 ( .A(\CARRYB[11][21] ), .B(\SUMB[11][22] ), .Z(\A1[31] ) );
  EOP U360 ( .A(\CARRYB[11][15] ), .B(\SUMB[11][16] ), .Z(\A1[25] ) );
  EOP U361 ( .A(\CARRYB[11][17] ), .B(\SUMB[11][18] ), .Z(\A1[27] ) );
  EOP U362 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A1[18] ) );
  IVP U363 ( .A(n230), .Z(n227) );
  IVP U364 ( .A(n230), .Z(n228) );
  EO U365 ( .A(\CARRYB[11][25] ), .B(\SUMB[11][26] ), .Z(\A1[35] ) );
  IVP U366 ( .A(n222), .Z(n219) );
  IVP U367 ( .A(n222), .Z(n220) );
  EO U368 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Z(\SUMB[1][28] ) );
  EO U369 ( .A(\CARRYB[11][27] ), .B(\SUMB[11][28] ), .Z(\A1[37] ) );
  IVP U370 ( .A(n243), .Z(n240) );
  IVP U371 ( .A(n243), .Z(n241) );
  IVP U372 ( .A(n247), .Z(n245) );
  IVP U373 ( .A(n247), .Z(n244) );
  IVP U374 ( .A(n251), .Z(n248) );
  IVP U375 ( .A(n251), .Z(n249) );
  IVP U376 ( .A(n255), .Z(n252) );
  IVP U377 ( .A(n255), .Z(n253) );
  IVP U378 ( .A(n226), .Z(n224) );
  IVP U379 ( .A(n226), .Z(n223) );
  IVP U380 ( .A(A[11]), .Z(n267) );
  EO U381 ( .A(\CARRYB[11][28] ), .B(\SUMB[11][29] ), .Z(\A1[38] ) );
  EO U382 ( .A(\CARRYB[11][29] ), .B(\ab[11][30] ), .Z(\A1[39] ) );
  EO U383 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A1[11] ) );
  IVP U384 ( .A(n261), .Z(n260) );
  IVP U385 ( .A(A[9]), .Z(n265) );
  EO U386 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A1[10] ) );
  EO U387 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Z(\SUMB[1][23] ) );
  EO U388 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\SUMB[1][17] ) );
  EO U389 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Z(\SUMB[1][25] ) );
  EO U390 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  IVP U391 ( .A(B[9]), .Z(n218) );
  EO U392 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U393 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U394 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U395 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  AN2P U396 ( .A(n236), .B(B[1]), .Z(n216) );
  EO U397 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Z(\SUMB[1][20] ) );
  EO U398 ( .A(\ab[0][2] ), .B(n216), .Z(\SUMB[1][1] ) );
  EO U399 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  IVP U400 ( .A(A[10]), .Z(n266) );
  AN2P U401 ( .A(\CARRYB[11][2] ), .B(\SUMB[11][3] ), .Z(\A2[13] ) );
  AN2P U402 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(\A2[14] ) );
  AN2P U403 ( .A(\CARRYB[11][4] ), .B(\SUMB[11][5] ), .Z(\A2[15] ) );
  AN2P U404 ( .A(\CARRYB[11][7] ), .B(\SUMB[11][8] ), .Z(\A2[18] ) );
  AN2P U405 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A2[20] ) );
  EOP U406 ( .A(\CARRYB[11][9] ), .B(\SUMB[11][10] ), .Z(\A1[19] ) );
  AN2P U407 ( .A(\CARRYB[11][16] ), .B(\SUMB[11][17] ), .Z(\A2[27] ) );
  AN2P U408 ( .A(\CARRYB[11][17] ), .B(\SUMB[11][18] ), .Z(\A2[28] ) );
  AN2P U409 ( .A(\CARRYB[11][19] ), .B(\SUMB[11][20] ), .Z(\A2[30] ) );
  EOP U410 ( .A(\CARRYB[11][19] ), .B(\SUMB[11][20] ), .Z(\A1[29] ) );
  AN2P U411 ( .A(\CARRYB[11][20] ), .B(\SUMB[11][21] ), .Z(\A2[31] ) );
  EOP U412 ( .A(\CARRYB[11][20] ), .B(\SUMB[11][21] ), .Z(\A1[30] ) );
  AN2P U413 ( .A(\CARRYB[11][22] ), .B(\SUMB[11][23] ), .Z(\A2[33] ) );
  AN2P U414 ( .A(\CARRYB[11][23] ), .B(\SUMB[11][24] ), .Z(\A2[34] ) );
  AN2P U415 ( .A(\CARRYB[11][26] ), .B(\SUMB[11][27] ), .Z(\A2[37] ) );
  EOP U416 ( .A(\CARRYB[11][26] ), .B(\SUMB[11][27] ), .Z(\A1[36] ) );
  AN2P U417 ( .A(\CARRYB[11][27] ), .B(\SUMB[11][28] ), .Z(\A2[38] ) );
  AN2P U418 ( .A(\CARRYB[11][28] ), .B(\SUMB[11][29] ), .Z(\A2[39] ) );
  AN2P U419 ( .A(\CARRYB[11][29] ), .B(\ab[11][30] ), .Z(\A2[40] ) );
  AN2P U420 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U421 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(\CARRYB[1][25] ) );
  AN2P U422 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(\CARRYB[1][28] ) );
  AN2P U423 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(\CARRYB[1][29] ) );
  AN2P U424 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A2[16] ) );
  EOP U425 ( .A(\CARRYB[11][5] ), .B(\SUMB[11][6] ), .Z(\A1[15] ) );
  AN2P U426 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U427 ( .A(\CARRYB[11][15] ), .B(\SUMB[11][16] ), .Z(\A2[26] ) );
  AN2P U428 ( .A(\CARRYB[11][12] ), .B(\SUMB[11][13] ), .Z(\A2[23] ) );
  EOP U429 ( .A(\CARRYB[11][12] ), .B(\SUMB[11][13] ), .Z(\A1[22] ) );
  AN2P U430 ( .A(n115), .B(\ab[0][17] ), .Z(\CARRYB[1][16] ) );
  AN2P U431 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U432 ( .A(\CARRYB[11][1] ), .B(\SUMB[11][2] ), .Z(\A2[12] ) );
  AN2P U433 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\CARRYB[1][17] ) );
  AN2P U434 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\CARRYB[1][21] ) );
  AN2P U435 ( .A(\CARRYB[11][21] ), .B(\SUMB[11][22] ), .Z(\A2[32] ) );
  AN2P U436 ( .A(\CARRYB[11][13] ), .B(\SUMB[11][14] ), .Z(\A2[24] ) );
  EOP U437 ( .A(\CARRYB[11][13] ), .B(\SUMB[11][14] ), .Z(\A1[23] ) );
  AN2P U438 ( .A(\CARRYB[11][6] ), .B(\SUMB[11][7] ), .Z(\A2[17] ) );
  AN2P U439 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U440 ( .A(\CARRYB[11][14] ), .B(\SUMB[11][15] ), .Z(\A2[25] ) );
  EOP U441 ( .A(\CARRYB[11][14] ), .B(\SUMB[11][15] ), .Z(\A1[24] ) );
  AN2P U442 ( .A(\CARRYB[11][24] ), .B(\SUMB[11][25] ), .Z(\A2[35] ) );
  AN2P U443 ( .A(\CARRYB[11][8] ), .B(\SUMB[11][9] ), .Z(\A2[19] ) );
  AN2P U444 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\CARRYB[1][18] ) );
  AN2P U445 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  EOP U446 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  AN2P U447 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A2[22] ) );
  EOP U448 ( .A(\CARRYB[11][11] ), .B(\SUMB[11][12] ), .Z(\A1[21] ) );
  AN2P U449 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U450 ( .A(\CARRYB[11][0] ), .B(\SUMB[11][1] ), .Z(\A2[11] ) );
  AN2P U451 ( .A(\CARRYB[11][25] ), .B(\SUMB[11][26] ), .Z(\A2[36] ) );
  AN2P U452 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U453 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(\CARRYB[1][24] ) );
  AN2P U454 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U455 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(\CARRYB[1][27] ) );
  AN2P U456 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U457 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A2[21] ) );
  EOP U458 ( .A(\CARRYB[11][10] ), .B(\SUMB[11][11] ), .Z(\A1[20] ) );
  AN2P U459 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U460 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U461 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(\CARRYB[1][22] ) );
  AN2P U462 ( .A(n216), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U463 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(\CARRYB[1][23] ) );
  AN2P U464 ( .A(\CARRYB[11][18] ), .B(\SUMB[11][19] ), .Z(\A2[29] ) );
  EOP U465 ( .A(\CARRYB[11][18] ), .B(\SUMB[11][19] ), .Z(\A1[28] ) );
  AN2P U466 ( .A(A[0]), .B(B[23]), .Z(\ab[0][23] ) );
  AN2 U467 ( .A(n233), .B(B[10]), .Z(\ab[0][10] ) );
  AN2 U468 ( .A(n58), .B(B[14]), .Z(\ab[0][14] ) );
  AN2 U469 ( .A(n234), .B(B[7]), .Z(\ab[0][7] ) );
  AN2 U470 ( .A(n233), .B(B[2]), .Z(\ab[0][2] ) );
  AN2 U471 ( .A(n234), .B(B[6]), .Z(\ab[0][6] ) );
  AN2P U472 ( .A(n58), .B(B[5]), .Z(\ab[0][5] ) );
  NR2 U473 ( .A(n235), .B(n218), .Z(\ab[0][9] ) );
  AN2P U474 ( .A(n189), .B(B[10]), .Z(\ab[1][10] ) );
  AN2P U475 ( .A(n189), .B(n258), .Z(\ab[1][26] ) );
  AN2P U476 ( .A(n189), .B(B[18]), .Z(\ab[1][18] ) );
  AN2P U477 ( .A(n217), .B(B[3]), .Z(\ab[1][3] ) );
  AN2P U478 ( .A(n189), .B(B[19]), .Z(\ab[1][19] ) );
  AN2P U479 ( .A(n189), .B(B[15]), .Z(\ab[1][15] ) );
  AN2P U480 ( .A(n237), .B(B[23]), .Z(\ab[1][23] ) );
  AN2P U481 ( .A(n236), .B(B[14]), .Z(\ab[1][14] ) );
  AN2P U482 ( .A(n217), .B(B[21]), .Z(\ab[1][21] ) );
  AN2 U483 ( .A(n233), .B(B[3]), .Z(\ab[0][3] ) );
  AN2 U484 ( .A(n233), .B(B[4]), .Z(\ab[0][4] ) );
  AN2P U485 ( .A(n189), .B(B[12]), .Z(\ab[1][12] ) );
  AN2P U486 ( .A(n217), .B(B[17]), .Z(\ab[1][17] ) );
  AN2P U487 ( .A(n236), .B(B[22]), .Z(\ab[1][22] ) );
  IVAP U488 ( .A(A[0]), .Z(n235) );
  AN2P U489 ( .A(n189), .B(B[20]), .Z(\ab[1][20] ) );
  AN2P U490 ( .A(n237), .B(B[13]), .Z(\ab[1][13] ) );
  AN2 U491 ( .A(n234), .B(B[24]), .Z(\ab[0][24] ) );
  AN2 U492 ( .A(n58), .B(B[13]), .Z(\ab[0][13] ) );
  AN2 U493 ( .A(n233), .B(B[21]), .Z(\ab[0][21] ) );
  AN2 U494 ( .A(n233), .B(B[22]), .Z(\ab[0][22] ) );
  AN2 U495 ( .A(n233), .B(B[15]), .Z(\ab[0][15] ) );
  IVA U496 ( .A(n222), .Z(n221) );
  IVA U497 ( .A(n262), .Z(n222) );
  IVA U498 ( .A(n226), .Z(n225) );
  IVA U499 ( .A(n263), .Z(n226) );
  IVA U500 ( .A(n230), .Z(n229) );
  IVA U501 ( .A(n264), .Z(n230) );
  IVA U502 ( .A(B[30]), .Z(n232) );
  IVA U503 ( .A(n243), .Z(n242) );
  IVA U504 ( .A(A[5]), .Z(n243) );
  IVA U505 ( .A(n247), .Z(n246) );
  IVA U506 ( .A(A[6]), .Z(n247) );
  IVA U507 ( .A(n251), .Z(n250) );
  IVA U508 ( .A(A[7]), .Z(n251) );
  IVA U509 ( .A(n255), .Z(n254) );
  IVA U510 ( .A(A[8]), .Z(n255) );
  IVA U511 ( .A(B[25]), .Z(n257) );
  IVA U512 ( .A(B[26]), .Z(n259) );
  IVA U513 ( .A(B[27]), .Z(n261) );
  AN2P U514 ( .A(n233), .B(n231), .Z(\ab[0][30] ) );
  AN2P U515 ( .A(n140), .B(n63), .Z(\ab[1][29] ) );
  AN2P U516 ( .A(n58), .B(n63), .Z(\ab[0][29] ) );
  AN2P U517 ( .A(n141), .B(n61), .Z(\ab[1][28] ) );
  AN2P U518 ( .A(n58), .B(n61), .Z(\ab[0][28] ) );
  AN2P U519 ( .A(n217), .B(n260), .Z(\ab[1][27] ) );
  AN2P U520 ( .A(n58), .B(n260), .Z(\ab[0][27] ) );
  AN2P U521 ( .A(n58), .B(n258), .Z(\ab[0][26] ) );
  AN2P U522 ( .A(n233), .B(n256), .Z(\ab[0][25] ) );
  AN2P U523 ( .A(n236), .B(B[24]), .Z(\ab[1][24] ) );
  AN2P U524 ( .A(n233), .B(B[17]), .Z(\ab[0][17] ) );
  AN2P U525 ( .A(n217), .B(B[11]), .Z(\ab[1][11] ) );
  AN2P U526 ( .A(n189), .B(B[9]), .Z(\ab[1][9] ) );
  AN2P U527 ( .A(n237), .B(B[8]), .Z(\ab[1][8] ) );
  AN2P U528 ( .A(n217), .B(B[7]), .Z(\ab[1][7] ) );
  AN2P U529 ( .A(n189), .B(B[6]), .Z(\ab[1][6] ) );
  AN2P U530 ( .A(n236), .B(B[5]), .Z(\ab[1][5] ) );
  AN2P U531 ( .A(n141), .B(B[2]), .Z(\ab[1][2] ) );
  AN2P U532 ( .A(n239), .B(n63), .Z(\ab[2][29] ) );
  AN2P U533 ( .A(n141), .B(n231), .Z(\ab[1][30] ) );
  AN2P U534 ( .A(n188), .B(n61), .Z(\ab[2][28] ) );
  AN2P U535 ( .A(n56), .B(n260), .Z(\ab[2][27] ) );
  AN2P U536 ( .A(n188), .B(n258), .Z(\ab[2][26] ) );
  AN2P U537 ( .A(n56), .B(n256), .Z(\ab[2][25] ) );
  AN2P U538 ( .A(n239), .B(B[24]), .Z(\ab[2][24] ) );
  AN2P U539 ( .A(n239), .B(B[23]), .Z(\ab[2][23] ) );
  AN2P U540 ( .A(n239), .B(B[22]), .Z(\ab[2][22] ) );
  AN2P U541 ( .A(n56), .B(B[21]), .Z(\ab[2][21] ) );
  AN2P U542 ( .A(n239), .B(B[20]), .Z(\ab[2][20] ) );
  AN2P U543 ( .A(n239), .B(B[19]), .Z(\ab[2][19] ) );
  AN2P U544 ( .A(n56), .B(B[18]), .Z(\ab[2][18] ) );
  AN2P U545 ( .A(n56), .B(B[17]), .Z(\ab[2][17] ) );
  AN2P U546 ( .A(n56), .B(B[16]), .Z(\ab[2][16] ) );
  AN2P U547 ( .A(n188), .B(B[15]), .Z(\ab[2][15] ) );
  AN2P U548 ( .A(n188), .B(B[14]), .Z(\ab[2][14] ) );
  AN2P U549 ( .A(n56), .B(B[13]), .Z(\ab[2][13] ) );
  AN2P U550 ( .A(n239), .B(B[12]), .Z(\ab[2][12] ) );
  AN2P U551 ( .A(n56), .B(B[11]), .Z(\ab[2][11] ) );
  AN2P U552 ( .A(n188), .B(B[10]), .Z(\ab[2][10] ) );
  AN2P U553 ( .A(n56), .B(B[9]), .Z(\ab[2][9] ) );
  AN2P U554 ( .A(n56), .B(B[8]), .Z(\ab[2][8] ) );
  AN2P U555 ( .A(n239), .B(B[7]), .Z(\ab[2][7] ) );
  AN2P U556 ( .A(n188), .B(B[6]), .Z(\ab[2][6] ) );
  AN2P U557 ( .A(n56), .B(B[5]), .Z(\ab[2][5] ) );
  AN2P U558 ( .A(n188), .B(B[4]), .Z(\ab[2][4] ) );
  AN2P U559 ( .A(n188), .B(B[3]), .Z(\ab[2][3] ) );
  AN2P U560 ( .A(n239), .B(B[2]), .Z(\ab[2][2] ) );
  AN2P U561 ( .A(n56), .B(B[1]), .Z(\ab[2][1] ) );
  AN2P U562 ( .A(n56), .B(B[0]), .Z(\ab[2][0] ) );
  AN3 U563 ( .A(n233), .B(B[0]), .C(n216), .Z(\CARRYB[1][0] ) );
  AN2P U564 ( .A(n215), .B(n63), .Z(\ab[3][29] ) );
  AN2P U565 ( .A(n56), .B(n231), .Z(\ab[2][30] ) );
  AN2P U566 ( .A(A[3]), .B(n61), .Z(\ab[3][28] ) );
  AN2P U567 ( .A(A[3]), .B(n260), .Z(\ab[3][27] ) );
  AN2P U568 ( .A(n215), .B(n258), .Z(\ab[3][26] ) );
  AN2P U569 ( .A(n215), .B(n256), .Z(\ab[3][25] ) );
  AN2P U570 ( .A(n215), .B(B[24]), .Z(\ab[3][24] ) );
  AN2P U571 ( .A(n215), .B(B[23]), .Z(\ab[3][23] ) );
  AN2P U572 ( .A(n215), .B(B[22]), .Z(\ab[3][22] ) );
  AN2P U573 ( .A(n215), .B(B[21]), .Z(\ab[3][21] ) );
  AN2P U574 ( .A(n215), .B(B[20]), .Z(\ab[3][20] ) );
  AN2P U575 ( .A(A[3]), .B(B[19]), .Z(\ab[3][19] ) );
  AN2P U576 ( .A(n215), .B(B[18]), .Z(\ab[3][18] ) );
  AN2P U577 ( .A(n215), .B(B[17]), .Z(\ab[3][17] ) );
  AN2P U578 ( .A(n215), .B(B[16]), .Z(\ab[3][16] ) );
  AN2P U579 ( .A(A[3]), .B(B[15]), .Z(\ab[3][15] ) );
  AN2P U580 ( .A(A[3]), .B(B[14]), .Z(\ab[3][14] ) );
  AN2P U581 ( .A(n215), .B(B[13]), .Z(\ab[3][13] ) );
  AN2P U582 ( .A(A[3]), .B(B[12]), .Z(\ab[3][12] ) );
  AN2P U583 ( .A(A[3]), .B(B[11]), .Z(\ab[3][11] ) );
  AN2P U584 ( .A(n215), .B(B[10]), .Z(\ab[3][10] ) );
  AN2P U585 ( .A(n215), .B(B[9]), .Z(\ab[3][9] ) );
  AN2P U586 ( .A(n215), .B(B[7]), .Z(\ab[3][7] ) );
  AN2P U587 ( .A(n215), .B(B[6]), .Z(\ab[3][6] ) );
  AN2P U588 ( .A(n215), .B(B[5]), .Z(\ab[3][5] ) );
  AN2P U589 ( .A(n215), .B(B[4]), .Z(\ab[3][4] ) );
  AN2P U590 ( .A(n215), .B(B[3]), .Z(\ab[3][3] ) );
  AN2P U591 ( .A(n215), .B(B[2]), .Z(\ab[3][2] ) );
  AN2P U592 ( .A(n215), .B(B[1]), .Z(\ab[3][1] ) );
  AN2P U593 ( .A(n215), .B(B[0]), .Z(\ab[3][0] ) );
  AN2P U594 ( .A(A[4]), .B(n63), .Z(\ab[4][29] ) );
  AN2P U595 ( .A(n215), .B(n231), .Z(\ab[3][30] ) );
  AN2P U596 ( .A(A[4]), .B(n61), .Z(\ab[4][28] ) );
  AN2P U597 ( .A(A[4]), .B(n260), .Z(\ab[4][27] ) );
  AN2P U598 ( .A(A[4]), .B(n258), .Z(\ab[4][26] ) );
  AN2P U599 ( .A(n59), .B(n256), .Z(\ab[4][25] ) );
  AN2P U600 ( .A(A[4]), .B(B[24]), .Z(\ab[4][24] ) );
  AN2P U601 ( .A(A[4]), .B(B[23]), .Z(\ab[4][23] ) );
  AN2P U602 ( .A(n59), .B(B[22]), .Z(\ab[4][22] ) );
  AN2P U603 ( .A(n59), .B(B[21]), .Z(\ab[4][21] ) );
  AN2P U604 ( .A(n59), .B(B[20]), .Z(\ab[4][20] ) );
  AN2P U605 ( .A(n59), .B(B[19]), .Z(\ab[4][19] ) );
  AN2P U606 ( .A(n59), .B(B[18]), .Z(\ab[4][18] ) );
  AN2P U607 ( .A(n59), .B(B[17]), .Z(\ab[4][17] ) );
  AN2P U608 ( .A(n59), .B(B[16]), .Z(\ab[4][16] ) );
  AN2P U609 ( .A(n59), .B(B[15]), .Z(\ab[4][15] ) );
  AN2P U610 ( .A(n59), .B(B[14]), .Z(\ab[4][14] ) );
  AN2P U611 ( .A(n59), .B(B[13]), .Z(\ab[4][13] ) );
  AN2P U612 ( .A(n59), .B(B[12]), .Z(\ab[4][12] ) );
  AN2P U613 ( .A(n59), .B(B[11]), .Z(\ab[4][11] ) );
  AN2P U614 ( .A(n59), .B(B[10]), .Z(\ab[4][10] ) );
  AN2P U615 ( .A(A[4]), .B(B[9]), .Z(\ab[4][9] ) );
  AN2P U616 ( .A(n59), .B(B[8]), .Z(\ab[4][8] ) );
  AN2P U617 ( .A(n59), .B(B[7]), .Z(\ab[4][7] ) );
  AN2P U618 ( .A(n59), .B(B[6]), .Z(\ab[4][6] ) );
  AN2P U619 ( .A(n59), .B(B[5]), .Z(\ab[4][5] ) );
  AN2P U620 ( .A(A[4]), .B(B[4]), .Z(\ab[4][4] ) );
  AN2P U621 ( .A(A[4]), .B(B[3]), .Z(\ab[4][3] ) );
  AN2P U622 ( .A(A[4]), .B(B[2]), .Z(\ab[4][2] ) );
  AN2P U623 ( .A(A[4]), .B(B[1]), .Z(\ab[4][1] ) );
  AN2P U624 ( .A(n59), .B(B[0]), .Z(\ab[4][0] ) );
  AN2P U625 ( .A(n242), .B(n63), .Z(\ab[5][29] ) );
  AN2P U626 ( .A(A[4]), .B(n231), .Z(\ab[4][30] ) );
  AN2P U627 ( .A(n242), .B(n61), .Z(\ab[5][28] ) );
  AN2P U628 ( .A(n242), .B(n260), .Z(\ab[5][27] ) );
  AN2P U629 ( .A(n242), .B(n258), .Z(\ab[5][26] ) );
  AN2P U630 ( .A(n242), .B(n256), .Z(\ab[5][25] ) );
  AN2P U631 ( .A(n242), .B(B[24]), .Z(\ab[5][24] ) );
  AN2P U632 ( .A(n242), .B(B[23]), .Z(\ab[5][23] ) );
  AN2P U633 ( .A(n241), .B(B[22]), .Z(\ab[5][22] ) );
  AN2P U634 ( .A(n241), .B(B[21]), .Z(\ab[5][21] ) );
  AN2P U635 ( .A(n241), .B(B[20]), .Z(\ab[5][20] ) );
  AN2P U636 ( .A(n241), .B(B[19]), .Z(\ab[5][19] ) );
  AN2P U637 ( .A(n241), .B(B[18]), .Z(\ab[5][18] ) );
  AN2P U638 ( .A(n241), .B(B[17]), .Z(\ab[5][17] ) );
  AN2P U639 ( .A(n241), .B(B[16]), .Z(\ab[5][16] ) );
  AN2P U640 ( .A(n241), .B(B[15]), .Z(\ab[5][15] ) );
  AN2P U641 ( .A(n241), .B(B[14]), .Z(\ab[5][14] ) );
  AN2P U642 ( .A(n241), .B(B[13]), .Z(\ab[5][13] ) );
  AN2P U643 ( .A(n241), .B(B[12]), .Z(\ab[5][12] ) );
  AN2P U644 ( .A(n241), .B(B[11]), .Z(\ab[5][11] ) );
  AN2P U645 ( .A(n240), .B(B[10]), .Z(\ab[5][10] ) );
  AN2P U646 ( .A(n240), .B(B[9]), .Z(\ab[5][9] ) );
  AN2P U647 ( .A(n240), .B(B[8]), .Z(\ab[5][8] ) );
  AN2P U648 ( .A(n240), .B(B[7]), .Z(\ab[5][7] ) );
  AN2P U649 ( .A(n240), .B(B[6]), .Z(\ab[5][6] ) );
  AN2P U650 ( .A(n240), .B(B[5]), .Z(\ab[5][5] ) );
  AN2P U651 ( .A(n240), .B(B[4]), .Z(\ab[5][4] ) );
  AN2P U652 ( .A(n240), .B(B[3]), .Z(\ab[5][3] ) );
  AN2P U653 ( .A(n240), .B(B[2]), .Z(\ab[5][2] ) );
  AN2P U654 ( .A(n240), .B(B[1]), .Z(\ab[5][1] ) );
  AN2P U655 ( .A(n240), .B(B[0]), .Z(\ab[5][0] ) );
  AN2P U656 ( .A(n246), .B(n63), .Z(\ab[6][29] ) );
  AN2P U657 ( .A(n240), .B(n231), .Z(\ab[5][30] ) );
  AN2P U658 ( .A(n246), .B(n61), .Z(\ab[6][28] ) );
  AN2P U659 ( .A(n246), .B(n260), .Z(\ab[6][27] ) );
  AN2P U660 ( .A(n246), .B(n258), .Z(\ab[6][26] ) );
  AN2P U661 ( .A(n246), .B(n256), .Z(\ab[6][25] ) );
  AN2P U662 ( .A(n246), .B(B[24]), .Z(\ab[6][24] ) );
  AN2P U663 ( .A(n246), .B(B[23]), .Z(\ab[6][23] ) );
  AN2P U664 ( .A(n245), .B(B[22]), .Z(\ab[6][22] ) );
  AN2P U665 ( .A(n245), .B(B[21]), .Z(\ab[6][21] ) );
  AN2P U666 ( .A(n245), .B(B[20]), .Z(\ab[6][20] ) );
  AN2P U667 ( .A(n245), .B(B[19]), .Z(\ab[6][19] ) );
  AN2P U668 ( .A(n245), .B(B[18]), .Z(\ab[6][18] ) );
  AN2P U669 ( .A(n245), .B(B[17]), .Z(\ab[6][17] ) );
  AN2P U670 ( .A(n245), .B(B[16]), .Z(\ab[6][16] ) );
  AN2P U671 ( .A(n245), .B(B[15]), .Z(\ab[6][15] ) );
  AN2P U672 ( .A(n245), .B(B[14]), .Z(\ab[6][14] ) );
  AN2P U673 ( .A(n245), .B(B[13]), .Z(\ab[6][13] ) );
  AN2P U674 ( .A(n245), .B(B[12]), .Z(\ab[6][12] ) );
  AN2P U675 ( .A(n245), .B(B[11]), .Z(\ab[6][11] ) );
  AN2P U676 ( .A(n244), .B(B[10]), .Z(\ab[6][10] ) );
  AN2P U677 ( .A(n244), .B(B[9]), .Z(\ab[6][9] ) );
  AN2P U678 ( .A(n244), .B(B[8]), .Z(\ab[6][8] ) );
  AN2P U679 ( .A(n244), .B(B[7]), .Z(\ab[6][7] ) );
  AN2P U680 ( .A(n244), .B(B[6]), .Z(\ab[6][6] ) );
  AN2P U681 ( .A(n244), .B(B[5]), .Z(\ab[6][5] ) );
  AN2P U682 ( .A(n244), .B(B[4]), .Z(\ab[6][4] ) );
  AN2P U683 ( .A(n244), .B(B[3]), .Z(\ab[6][3] ) );
  AN2P U684 ( .A(n244), .B(B[2]), .Z(\ab[6][2] ) );
  AN2P U685 ( .A(n244), .B(B[1]), .Z(\ab[6][1] ) );
  AN2P U686 ( .A(n244), .B(B[0]), .Z(\ab[6][0] ) );
  AN2P U687 ( .A(n250), .B(n63), .Z(\ab[7][29] ) );
  AN2P U688 ( .A(n244), .B(n231), .Z(\ab[6][30] ) );
  AN2P U689 ( .A(n250), .B(n61), .Z(\ab[7][28] ) );
  AN2P U690 ( .A(n250), .B(n260), .Z(\ab[7][27] ) );
  AN2P U691 ( .A(n250), .B(n258), .Z(\ab[7][26] ) );
  AN2P U692 ( .A(n250), .B(n256), .Z(\ab[7][25] ) );
  AN2P U693 ( .A(n250), .B(B[24]), .Z(\ab[7][24] ) );
  AN2P U694 ( .A(n250), .B(B[23]), .Z(\ab[7][23] ) );
  AN2P U695 ( .A(n249), .B(B[22]), .Z(\ab[7][22] ) );
  AN2P U696 ( .A(n249), .B(B[21]), .Z(\ab[7][21] ) );
  AN2P U697 ( .A(n249), .B(B[20]), .Z(\ab[7][20] ) );
  AN2P U698 ( .A(n249), .B(B[19]), .Z(\ab[7][19] ) );
  AN2P U699 ( .A(n249), .B(B[18]), .Z(\ab[7][18] ) );
  AN2P U700 ( .A(n249), .B(B[17]), .Z(\ab[7][17] ) );
  AN2P U701 ( .A(n249), .B(B[16]), .Z(\ab[7][16] ) );
  AN2P U702 ( .A(n249), .B(B[15]), .Z(\ab[7][15] ) );
  AN2P U703 ( .A(n249), .B(B[14]), .Z(\ab[7][14] ) );
  AN2P U704 ( .A(n249), .B(B[13]), .Z(\ab[7][13] ) );
  AN2P U705 ( .A(n249), .B(B[12]), .Z(\ab[7][12] ) );
  AN2P U706 ( .A(n249), .B(B[11]), .Z(\ab[7][11] ) );
  AN2P U707 ( .A(n248), .B(B[10]), .Z(\ab[7][10] ) );
  AN2P U708 ( .A(n248), .B(B[9]), .Z(\ab[7][9] ) );
  AN2P U709 ( .A(n248), .B(B[8]), .Z(\ab[7][8] ) );
  AN2P U710 ( .A(n248), .B(B[7]), .Z(\ab[7][7] ) );
  AN2P U711 ( .A(n248), .B(B[6]), .Z(\ab[7][6] ) );
  AN2P U712 ( .A(n248), .B(B[5]), .Z(\ab[7][5] ) );
  AN2P U713 ( .A(n248), .B(B[4]), .Z(\ab[7][4] ) );
  AN2P U714 ( .A(n248), .B(B[3]), .Z(\ab[7][3] ) );
  AN2P U715 ( .A(n248), .B(B[2]), .Z(\ab[7][2] ) );
  AN2P U716 ( .A(n248), .B(B[1]), .Z(\ab[7][1] ) );
  AN2P U717 ( .A(n248), .B(B[0]), .Z(\ab[7][0] ) );
  AN2P U718 ( .A(n254), .B(n63), .Z(\ab[8][29] ) );
  AN2P U719 ( .A(n248), .B(n231), .Z(\ab[7][30] ) );
  AN2P U720 ( .A(n254), .B(n61), .Z(\ab[8][28] ) );
  AN2P U721 ( .A(n254), .B(n260), .Z(\ab[8][27] ) );
  AN2P U722 ( .A(n254), .B(n258), .Z(\ab[8][26] ) );
  AN2P U723 ( .A(n254), .B(n256), .Z(\ab[8][25] ) );
  AN2P U724 ( .A(n254), .B(B[24]), .Z(\ab[8][24] ) );
  AN2P U725 ( .A(n254), .B(B[23]), .Z(\ab[8][23] ) );
  AN2P U726 ( .A(n253), .B(B[22]), .Z(\ab[8][22] ) );
  AN2P U727 ( .A(n253), .B(B[21]), .Z(\ab[8][21] ) );
  AN2P U728 ( .A(n253), .B(B[20]), .Z(\ab[8][20] ) );
  AN2P U729 ( .A(n253), .B(B[19]), .Z(\ab[8][19] ) );
  AN2P U730 ( .A(n253), .B(B[18]), .Z(\ab[8][18] ) );
  AN2P U731 ( .A(n253), .B(B[17]), .Z(\ab[8][17] ) );
  AN2P U732 ( .A(n253), .B(B[16]), .Z(\ab[8][16] ) );
  AN2P U733 ( .A(n253), .B(B[15]), .Z(\ab[8][15] ) );
  AN2P U734 ( .A(n253), .B(B[14]), .Z(\ab[8][14] ) );
  AN2P U735 ( .A(n253), .B(B[13]), .Z(\ab[8][13] ) );
  AN2P U736 ( .A(n253), .B(B[12]), .Z(\ab[8][12] ) );
  AN2P U737 ( .A(n253), .B(B[11]), .Z(\ab[8][11] ) );
  AN2P U738 ( .A(n252), .B(B[10]), .Z(\ab[8][10] ) );
  AN2P U739 ( .A(n252), .B(B[9]), .Z(\ab[8][9] ) );
  AN2P U740 ( .A(n252), .B(B[8]), .Z(\ab[8][8] ) );
  AN2P U741 ( .A(n252), .B(B[7]), .Z(\ab[8][7] ) );
  AN2P U742 ( .A(n252), .B(B[6]), .Z(\ab[8][6] ) );
  AN2P U743 ( .A(n252), .B(B[5]), .Z(\ab[8][5] ) );
  AN2P U744 ( .A(n252), .B(B[4]), .Z(\ab[8][4] ) );
  AN2P U745 ( .A(n252), .B(B[3]), .Z(\ab[8][3] ) );
  AN2P U746 ( .A(n252), .B(B[2]), .Z(\ab[8][2] ) );
  AN2P U747 ( .A(n252), .B(B[1]), .Z(\ab[8][1] ) );
  AN2P U748 ( .A(n252), .B(B[0]), .Z(\ab[8][0] ) );
  AN2P U749 ( .A(n252), .B(n231), .Z(\ab[8][30] ) );
  IVA U750 ( .A(n265), .Z(n262) );
  AN2P U751 ( .A(B[24]), .B(n221), .Z(\ab[9][24] ) );
  AN2P U752 ( .A(B[23]), .B(n220), .Z(\ab[9][23] ) );
  AN2P U753 ( .A(B[22]), .B(n220), .Z(\ab[9][22] ) );
  AN2P U754 ( .A(B[21]), .B(n220), .Z(\ab[9][21] ) );
  AN2P U755 ( .A(B[20]), .B(n220), .Z(\ab[9][20] ) );
  AN2P U756 ( .A(B[19]), .B(n220), .Z(\ab[9][19] ) );
  AN2P U757 ( .A(B[18]), .B(n220), .Z(\ab[9][18] ) );
  AN2P U758 ( .A(B[17]), .B(n220), .Z(\ab[9][17] ) );
  AN2P U759 ( .A(B[16]), .B(n220), .Z(\ab[9][16] ) );
  AN2P U760 ( .A(B[15]), .B(n220), .Z(\ab[9][15] ) );
  AN2P U761 ( .A(B[14]), .B(n220), .Z(\ab[9][14] ) );
  AN2P U762 ( .A(B[13]), .B(n220), .Z(\ab[9][13] ) );
  AN2P U763 ( .A(B[12]), .B(n220), .Z(\ab[9][12] ) );
  AN2P U764 ( .A(B[11]), .B(n219), .Z(\ab[9][11] ) );
  AN2P U765 ( .A(B[10]), .B(n219), .Z(\ab[9][10] ) );
  AN2P U766 ( .A(B[9]), .B(n219), .Z(\ab[9][9] ) );
  AN2P U767 ( .A(B[8]), .B(n219), .Z(\ab[9][8] ) );
  AN2P U768 ( .A(B[7]), .B(n219), .Z(\ab[9][7] ) );
  AN2P U769 ( .A(B[6]), .B(n219), .Z(\ab[9][6] ) );
  AN2P U770 ( .A(B[5]), .B(n219), .Z(\ab[9][5] ) );
  AN2P U771 ( .A(B[4]), .B(n219), .Z(\ab[9][4] ) );
  AN2P U772 ( .A(B[3]), .B(n219), .Z(\ab[9][3] ) );
  AN2P U773 ( .A(B[2]), .B(n219), .Z(\ab[9][2] ) );
  AN2P U774 ( .A(B[1]), .B(n219), .Z(\ab[9][1] ) );
  AN2P U775 ( .A(B[0]), .B(n219), .Z(\ab[9][0] ) );
  IVA U776 ( .A(n266), .Z(n263) );
  AN2P U777 ( .A(B[24]), .B(n225), .Z(\ab[10][24] ) );
  AN2P U778 ( .A(B[23]), .B(n224), .Z(\ab[10][23] ) );
  AN2P U779 ( .A(B[22]), .B(n224), .Z(\ab[10][22] ) );
  AN2P U780 ( .A(B[21]), .B(n224), .Z(\ab[10][21] ) );
  AN2P U781 ( .A(B[20]), .B(n224), .Z(\ab[10][20] ) );
  AN2P U782 ( .A(B[19]), .B(n224), .Z(\ab[10][19] ) );
  AN2P U783 ( .A(B[18]), .B(n224), .Z(\ab[10][18] ) );
  AN2P U784 ( .A(B[17]), .B(n224), .Z(\ab[10][17] ) );
  AN2P U785 ( .A(B[16]), .B(n224), .Z(\ab[10][16] ) );
  AN2P U786 ( .A(B[15]), .B(n224), .Z(\ab[10][15] ) );
  AN2P U787 ( .A(B[14]), .B(n224), .Z(\ab[10][14] ) );
  AN2P U788 ( .A(B[13]), .B(n224), .Z(\ab[10][13] ) );
  AN2P U789 ( .A(B[12]), .B(n224), .Z(\ab[10][12] ) );
  AN2P U790 ( .A(B[11]), .B(n223), .Z(\ab[10][11] ) );
  AN2P U791 ( .A(B[10]), .B(n223), .Z(\ab[10][10] ) );
  AN2P U792 ( .A(B[9]), .B(n223), .Z(\ab[10][9] ) );
  AN2P U793 ( .A(B[8]), .B(n223), .Z(\ab[10][8] ) );
  AN2P U794 ( .A(B[7]), .B(n223), .Z(\ab[10][7] ) );
  AN2P U795 ( .A(B[6]), .B(n223), .Z(\ab[10][6] ) );
  AN2P U796 ( .A(B[5]), .B(n223), .Z(\ab[10][5] ) );
  AN2P U797 ( .A(B[4]), .B(n223), .Z(\ab[10][4] ) );
  AN2P U798 ( .A(B[3]), .B(n223), .Z(\ab[10][3] ) );
  AN2P U799 ( .A(B[2]), .B(n223), .Z(\ab[10][2] ) );
  AN2P U800 ( .A(B[1]), .B(n223), .Z(\ab[10][1] ) );
  AN2P U801 ( .A(B[0]), .B(n223), .Z(\ab[10][0] ) );
  IVA U802 ( .A(n267), .Z(n264) );
  AN2P U803 ( .A(B[24]), .B(n229), .Z(\ab[11][24] ) );
  AN2P U804 ( .A(B[23]), .B(n228), .Z(\ab[11][23] ) );
  AN2P U805 ( .A(B[22]), .B(n228), .Z(\ab[11][22] ) );
  AN2P U806 ( .A(B[21]), .B(n228), .Z(\ab[11][21] ) );
  AN2P U807 ( .A(B[20]), .B(n228), .Z(\ab[11][20] ) );
  AN2P U808 ( .A(B[19]), .B(n228), .Z(\ab[11][19] ) );
  AN2P U809 ( .A(B[18]), .B(n228), .Z(\ab[11][18] ) );
  AN2P U810 ( .A(B[17]), .B(n228), .Z(\ab[11][17] ) );
  AN2P U811 ( .A(B[16]), .B(n228), .Z(\ab[11][16] ) );
  AN2P U812 ( .A(B[15]), .B(n228), .Z(\ab[11][15] ) );
  AN2P U813 ( .A(B[14]), .B(n228), .Z(\ab[11][14] ) );
  AN2P U814 ( .A(B[13]), .B(n228), .Z(\ab[11][13] ) );
  AN2P U815 ( .A(B[12]), .B(n228), .Z(\ab[11][12] ) );
  AN2P U816 ( .A(B[11]), .B(n227), .Z(\ab[11][11] ) );
  AN2P U817 ( .A(B[10]), .B(n227), .Z(\ab[11][10] ) );
  AN2P U818 ( .A(B[9]), .B(n227), .Z(\ab[11][9] ) );
  AN2P U819 ( .A(B[8]), .B(n227), .Z(\ab[11][8] ) );
  AN2P U820 ( .A(B[7]), .B(n227), .Z(\ab[11][7] ) );
  AN2P U821 ( .A(B[6]), .B(n227), .Z(\ab[11][6] ) );
  AN2P U822 ( .A(B[5]), .B(n227), .Z(\ab[11][5] ) );
  AN2P U823 ( .A(B[4]), .B(n227), .Z(\ab[11][4] ) );
  AN2P U824 ( .A(B[3]), .B(n227), .Z(\ab[11][3] ) );
  AN2P U825 ( .A(B[2]), .B(n227), .Z(\ab[11][2] ) );
  AN2P U826 ( .A(B[1]), .B(n227), .Z(\ab[11][1] ) );
  AN2P U827 ( .A(B[0]), .B(n227), .Z(\ab[11][0] ) );
  NR2 U829 ( .A(n265), .B(n232), .Z(\ab[9][30] ) );
  NR2 U830 ( .A(n265), .B(n62), .Z(\ab[9][29] ) );
  NR2 U831 ( .A(n265), .B(n60), .Z(\ab[9][28] ) );
  NR2 U832 ( .A(n265), .B(n261), .Z(\ab[9][27] ) );
  NR2 U833 ( .A(n265), .B(n259), .Z(\ab[9][26] ) );
  NR2 U834 ( .A(n265), .B(n257), .Z(\ab[9][25] ) );
  NR2 U835 ( .A(n232), .B(n267), .Z(\ab[11][30] ) );
  NR2 U836 ( .A(n62), .B(n267), .Z(\ab[11][29] ) );
  NR2 U837 ( .A(n60), .B(n267), .Z(\ab[11][28] ) );
  NR2 U838 ( .A(n261), .B(n267), .Z(\ab[11][27] ) );
  NR2 U839 ( .A(n259), .B(n267), .Z(\ab[11][26] ) );
  NR2 U840 ( .A(n257), .B(n267), .Z(\ab[11][25] ) );
  NR2 U841 ( .A(n232), .B(n266), .Z(\ab[10][30] ) );
  NR2 U842 ( .A(n62), .B(n266), .Z(\ab[10][29] ) );
  NR2 U843 ( .A(n60), .B(n266), .Z(\ab[10][28] ) );
  NR2 U844 ( .A(n261), .B(n266), .Z(\ab[10][27] ) );
  NR2 U845 ( .A(n259), .B(n266), .Z(\ab[10][26] ) );
  NR2 U846 ( .A(n257), .B(n266), .Z(\ab[10][25] ) );
endmodule


module SQRT_POLY ( clk, reset, RootIn, RootOut );
  input [30:0] RootIn;
  output [16:0] RootOut;
  input clk, reset;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N70, N71, N72, N73, n90, n91, n92, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415;
  wire   [39:23] Term1;
  wire   [19:4] Term2;
  wire   [13:0] FractionBit;
  wire   [39:36] Term11;
  wire   [19:17] Term21;
  wire   [3:0] IntegerBits;
  wire   [12:0] Root;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25;
  assign N36 = RootIn[30];

  AN2P U1886 ( .A(Term11[37]), .B(n97), .Z(n96) );
  SQRT_POLY_DW01_add_0 add_39 ( .A({1'b0, Term1[35:23]}), .B({1'b0, 
        Term2[16:4]}), .CI(1'b0), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, 
        N57, N56, N55, N54, N53, N52}) );
  SQRT_POLY_DW02_mult_0 mult_34 ( .A({N7, N8, N9, N10, N11, N12, N13, N14, N15, 
        N16, N17, N18}), .B({n156, n177, RootIn[28:0]}), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25}) );
  FD1 \Term1_reg[39]  ( .D(n145), .CP(clk), .Q(Term1[39]) );
  FD1 \Term1_reg[36]  ( .D(n143), .CP(clk), .Q(Term1[36]) );
  FD1 \Term1_reg[35]  ( .D(n141), .CP(clk), .Q(Term1[35]) );
  FD1 \Term1_reg[38]  ( .D(n139), .CP(clk), .Q(Term1[38]) );
  FDS2L \Term1_reg[33]  ( .CR(1'b1), .D(N29), .LD(n153), .CP(clk), .Q(
        Term1[33]) );
  FDS2L \Term11_reg[39]  ( .CR(1'b1), .D(Term1[39]), .LD(n150), .CP(clk), .Q(
        Term11[39]) );
  FDS2L \Term2_reg[16]  ( .CR(1'b1), .D(N39), .LD(n152), .CP(clk), .Q(
        Term2[16]) );
  FDS2L \Term21_reg[19]  ( .CR(1'b1), .D(Term2[19]), .LD(n150), .CP(clk), .Q(
        Term21[19]) );
  FDS2L \Term11_reg[38]  ( .CR(1'b1), .D(Term1[38]), .LD(n150), .CP(clk), .Q(
        Term11[38]) );
  FDS2L \Term1_reg[34]  ( .CR(1'b1), .D(N30), .LD(n153), .CP(clk), .Q(
        Term1[34]) );
  FDS2L \Term2_reg[15]  ( .CR(1'b1), .D(N40), .LD(n152), .CP(clk), .Q(
        Term2[15]) );
  FDS2L \Term2_reg[14]  ( .CR(1'b1), .D(N41), .LD(n152), .CP(clk), .Q(
        Term2[14]) );
  FDS2L \Term21_reg[18]  ( .CR(1'b1), .D(Term2[18]), .LD(n149), .CP(clk), .Q(
        Term21[18]) );
  FDS2L \Term1_reg[32]  ( .CR(1'b1), .D(N28), .LD(n153), .CP(clk), .Q(
        Term1[32]) );
  FDS2L \Term2_reg[13]  ( .CR(1'b1), .D(N42), .LD(n152), .CP(clk), .Q(
        Term2[13]) );
  FDS2L \Term11_reg[37]  ( .CR(1'b1), .D(Term1[37]), .LD(n150), .CP(clk), .Q(
        Term11[37]) );
  FDS2L \Term21_reg[17]  ( .CR(1'b1), .D(Term2[17]), .LD(n149), .CP(clk), .Q(
        Term21[17]), .QN(n92) );
  FDS2L \FractionBit_reg[13]  ( .CR(1'b1), .D(N65), .LD(n151), .CP(clk), .Q(
        FractionBit[13]), .QN(n90) );
  FDS2L \Term11_reg[36]  ( .CR(1'b1), .D(Term1[36]), .LD(n150), .CP(clk), .Q(
        Term11[36]), .QN(n91) );
  FDS2L \Term1_reg[31]  ( .CR(1'b1), .D(N27), .LD(n153), .CP(clk), .Q(
        Term1[31]) );
  FDS2L \Term2_reg[12]  ( .CR(1'b1), .D(N43), .LD(n152), .CP(clk), .Q(
        Term2[12]) );
  FDS2L \Term1_reg[30]  ( .CR(1'b1), .D(N26), .LD(n153), .CP(clk), .Q(
        Term1[30]) );
  FDS2L \Term2_reg[11]  ( .CR(1'b1), .D(N44), .LD(n152), .CP(clk), .Q(
        Term2[11]) );
  FDS2L \Term1_reg[29]  ( .CR(1'b1), .D(N25), .LD(n153), .CP(clk), .Q(
        Term1[29]) );
  FDS2L \Term2_reg[10]  ( .CR(1'b1), .D(N45), .LD(n152), .CP(clk), .Q(
        Term2[10]) );
  FDS2L \Term1_reg[28]  ( .CR(1'b1), .D(N24), .LD(n153), .CP(clk), .Q(
        Term1[28]) );
  FDS2L \Term2_reg[9]  ( .CR(1'b1), .D(n135), .LD(n152), .CP(clk), .Q(Term2[9]) );
  FDS2L \Term1_reg[27]  ( .CR(1'b1), .D(N23), .LD(n153), .CP(clk), .Q(
        Term1[27]) );
  FDS2L \Term2_reg[8]  ( .CR(1'b1), .D(N47), .LD(n151), .CP(clk), .Q(Term2[8])
         );
  FDS2L \Term1_reg[26]  ( .CR(1'b1), .D(N22), .LD(n153), .CP(clk), .Q(
        Term1[26]) );
  FDS2L \Term2_reg[7]  ( .CR(1'b1), .D(N48), .LD(n151), .CP(clk), .Q(Term2[7])
         );
  FDS2L \Term1_reg[25]  ( .CR(1'b1), .D(N21), .LD(n153), .CP(clk), .Q(
        Term1[25]) );
  FDS2L \Term2_reg[6]  ( .CR(1'b1), .D(N49), .LD(n151), .CP(clk), .Q(Term2[6])
         );
  FDS2L \Term1_reg[24]  ( .CR(1'b1), .D(N20), .LD(n153), .CP(clk), .Q(
        Term1[24]) );
  FDS2L \Term1_reg[23]  ( .CR(1'b1), .D(N19), .LD(n152), .CP(clk), .Q(
        Term1[23]) );
  FDS2L \Term2_reg[5]  ( .CR(1'b1), .D(N50), .LD(n151), .CP(clk), .Q(Term2[5])
         );
  FDS2L \Term2_reg[4]  ( .CR(1'b1), .D(N51), .LD(n151), .CP(clk), .Q(Term2[4])
         );
  FDS2L \FractionBit_reg[12]  ( .CR(1'b1), .D(N64), .LD(n151), .CP(clk), .Q(
        FractionBit[12]) );
  FDS2L \FractionBit_reg[11]  ( .CR(1'b1), .D(N63), .LD(n151), .CP(clk), .Q(
        FractionBit[11]) );
  FDS2L \FractionBit_reg[10]  ( .CR(1'b1), .D(N62), .LD(n151), .CP(clk), .Q(
        FractionBit[10]) );
  FDS2L \FractionBit_reg[9]  ( .CR(1'b1), .D(N61), .LD(n151), .CP(clk), .Q(
        FractionBit[9]) );
  FDS2L \FractionBit_reg[8]  ( .CR(1'b1), .D(N60), .LD(n151), .CP(clk), .Q(
        FractionBit[8]) );
  FDS2L \FractionBit_reg[7]  ( .CR(1'b1), .D(N59), .LD(n151), .CP(clk), .Q(
        FractionBit[7]) );
  FDS2L \FractionBit_reg[6]  ( .CR(1'b1), .D(N58), .LD(n150), .CP(clk), .Q(
        FractionBit[6]) );
  FDS2L \FractionBit_reg[5]  ( .CR(1'b1), .D(N57), .LD(n150), .CP(clk), .Q(
        FractionBit[5]) );
  FDS2L \FractionBit_reg[4]  ( .CR(1'b1), .D(N56), .LD(n150), .CP(clk), .Q(
        FractionBit[4]) );
  FDS2L \FractionBit_reg[3]  ( .CR(1'b1), .D(N55), .LD(n150), .CP(clk), .Q(
        FractionBit[3]) );
  FDS2L \FractionBit_reg[2]  ( .CR(1'b1), .D(N54), .LD(n150), .CP(clk), .Q(
        FractionBit[2]) );
  FDS2L \FractionBit_reg[1]  ( .CR(1'b1), .D(N53), .LD(n150), .CP(clk), .Q(
        FractionBit[1]) );
  FDS2L \FractionBit_reg[0]  ( .CR(1'b1), .D(N52), .LD(n150), .CP(clk), .Q(
        FractionBit[0]) );
  FDS2L \IntegerBits_reg[3]  ( .CR(1'b1), .D(N73), .LD(n149), .CP(clk), .Q(
        IntegerBits[3]) );
  FDS2L \IntegerBits_reg[2]  ( .CR(1'b1), .D(N72), .LD(n149), .CP(clk), .Q(
        IntegerBits[2]) );
  FDS2L \IntegerBits_reg[1]  ( .CR(1'b1), .D(N71), .LD(n149), .CP(clk), .Q(
        IntegerBits[1]) );
  FDS2L \IntegerBits_reg[0]  ( .CR(1'b1), .D(N70), .LD(n149), .CP(clk), .Q(
        IntegerBits[0]) );
  FDS2L \RootOut_reg[16]  ( .CR(1'b1), .D(IntegerBits[3]), .LD(n148), .CP(clk), 
        .Q(RootOut[16]) );
  FDS2L \RootOut_reg[15]  ( .CR(1'b1), .D(IntegerBits[2]), .LD(n148), .CP(clk), 
        .Q(RootOut[15]) );
  FDS2L \RootOut_reg[14]  ( .CR(1'b1), .D(IntegerBits[1]), .LD(n148), .CP(clk), 
        .Q(RootOut[14]) );
  FDS2L \RootOut_reg[13]  ( .CR(1'b1), .D(IntegerBits[0]), .LD(n148), .CP(clk), 
        .Q(RootOut[13]) );
  FDS2L \RootOut_reg[12]  ( .CR(1'b1), .D(Root[12]), .LD(n148), .CP(clk), .Q(
        RootOut[12]) );
  FDS2L \RootOut_reg[11]  ( .CR(1'b1), .D(Root[11]), .LD(n147), .CP(clk), .Q(
        RootOut[11]) );
  FDS2L \RootOut_reg[10]  ( .CR(1'b1), .D(Root[10]), .LD(n147), .CP(clk), .Q(
        RootOut[10]) );
  FDS2L \RootOut_reg[9]  ( .CR(1'b1), .D(Root[9]), .LD(n147), .CP(clk), .Q(
        RootOut[9]) );
  FDS2L \RootOut_reg[8]  ( .CR(1'b1), .D(Root[8]), .LD(n147), .CP(clk), .Q(
        RootOut[8]) );
  FDS2L \RootOut_reg[7]  ( .CR(1'b1), .D(Root[7]), .LD(n147), .CP(clk), .Q(
        RootOut[7]) );
  FDS2L \RootOut_reg[6]  ( .CR(1'b1), .D(Root[6]), .LD(n147), .CP(clk), .Q(
        RootOut[6]) );
  FDS2L \RootOut_reg[5]  ( .CR(1'b1), .D(Root[5]), .LD(n147), .CP(clk), .Q(
        RootOut[5]) );
  FDS2L \RootOut_reg[4]  ( .CR(1'b1), .D(Root[4]), .LD(n147), .CP(clk), .Q(
        RootOut[4]) );
  FDS2L \RootOut_reg[3]  ( .CR(1'b1), .D(Root[3]), .LD(n147), .CP(clk), .Q(
        RootOut[3]) );
  FDS2L \RootOut_reg[2]  ( .CR(1'b1), .D(Root[2]), .LD(n147), .CP(clk), .Q(
        RootOut[2]) );
  FDS2L \RootOut_reg[1]  ( .CR(1'b1), .D(Root[1]), .LD(n147), .CP(clk), .Q(
        RootOut[1]) );
  FDS2L \RootOut_reg[0]  ( .CR(1'b1), .D(Root[0]), .LD(n147), .CP(clk), .Q(
        RootOut[0]) );
  FDS2L \Term2_reg[19]  ( .CR(1'b1), .D(n128), .LD(n152), .CP(clk), .Q(
        Term2[19]) );
  FDS2L \Term2_reg[18]  ( .CR(1'b1), .D(N37), .LD(n152), .CP(clk), .Q(
        Term2[18]) );
  FDS2L \Term2_reg[17]  ( .CR(1'b1), .D(N38), .LD(n152), .CP(clk), .Q(
        Term2[17]) );
  FDS2L \Root_reg[12]  ( .CR(1'b1), .D(FractionBit[12]), .LD(n149), .CP(clk), 
        .Q(Root[12]) );
  FDS2L \Root_reg[11]  ( .CR(1'b1), .D(FractionBit[11]), .LD(n149), .CP(clk), 
        .Q(Root[11]) );
  FDS2L \Root_reg[10]  ( .CR(1'b1), .D(FractionBit[10]), .LD(n149), .CP(clk), 
        .Q(Root[10]) );
  FDS2L \Root_reg[9]  ( .CR(1'b1), .D(FractionBit[9]), .LD(n149), .CP(clk), 
        .Q(Root[9]) );
  FDS2L \Root_reg[8]  ( .CR(1'b1), .D(FractionBit[8]), .LD(n149), .CP(clk), 
        .Q(Root[8]) );
  FDS2L \Root_reg[7]  ( .CR(1'b1), .D(FractionBit[7]), .LD(n149), .CP(clk), 
        .Q(Root[7]) );
  FDS2L \Root_reg[6]  ( .CR(1'b1), .D(FractionBit[6]), .LD(n148), .CP(clk), 
        .Q(Root[6]) );
  FDS2L \Root_reg[5]  ( .CR(1'b1), .D(FractionBit[5]), .LD(n148), .CP(clk), 
        .Q(Root[5]) );
  FDS2L \Root_reg[4]  ( .CR(1'b1), .D(FractionBit[4]), .LD(n148), .CP(clk), 
        .Q(Root[4]) );
  FDS2L \Root_reg[3]  ( .CR(1'b1), .D(FractionBit[3]), .LD(n148), .CP(clk), 
        .Q(Root[3]) );
  FDS2L \Root_reg[2]  ( .CR(1'b1), .D(FractionBit[2]), .LD(n148), .CP(clk), 
        .Q(Root[2]) );
  FDS2L \Root_reg[1]  ( .CR(1'b1), .D(FractionBit[1]), .LD(n148), .CP(clk), 
        .Q(Root[1]) );
  FDS2L \Root_reg[0]  ( .CR(1'b1), .D(FractionBit[0]), .LD(n148), .CP(clk), 
        .Q(Root[0]) );
  FDS2L \Term1_reg[37]  ( .CR(1'b1), .D(N33), .LD(n154), .CP(clk), .Q(
        Term1[37]) );
  B5I U1901 ( .A(n138), .Z(n139) );
  IVP U1902 ( .A(RootIn[27]), .Z(n105) );
  IVP U1903 ( .A(RootIn[27]), .Z(n106) );
  ND2P U1904 ( .A(RootIn[26]), .B(n173), .Z(n217) );
  IVP U1905 ( .A(n125), .Z(n386) );
  IVP U1906 ( .A(RootIn[25]), .Z(n120) );
  ND3 U1907 ( .A(RootIn[29]), .B(RootIn[28]), .C(N36), .Z(n184) );
  EO U1908 ( .A(RootIn[25]), .B(RootIn[26]), .Z(n181) );
  AO3 U1909 ( .A(n173), .B(n188), .C(n187), .D(n186), .Z(n195) );
  ND2 U1910 ( .A(n178), .B(n181), .Z(n188) );
  AO7 U1911 ( .A(RootIn[28]), .B(n185), .C(n184), .Z(n186) );
  ND2 U1912 ( .A(n183), .B(n182), .Z(n187) );
  IVP U1913 ( .A(RootIn[25]), .Z(n164) );
  IVP U1914 ( .A(n387), .Z(n339) );
  IVP U1915 ( .A(n123), .Z(n163) );
  ND2 U1916 ( .A(n174), .B(n160), .Z(n304) );
  MUX41 U1917 ( .D0(n345), .D1(n344), .D2(n343), .D3(n342), .A(n177), .B(n128), 
        .Z(n346) );
  IVP U1918 ( .A(n140), .Z(n141) );
  IVP U1919 ( .A(n142), .Z(n143) );
  IVP U1920 ( .A(n144), .Z(n145) );
  MUX51HP U1921 ( .D0(n354), .D1(n280), .D2(n350), .D3(n130), .D4(n234), .A(
        n156), .B(n176), .C(RootIn[28]), .Z(N14) );
  AN2P U1922 ( .A(RootIn[26]), .B(n164), .Z(n107) );
  IVP U1923 ( .A(RootIn[28]), .Z(n175) );
  IVDAP U1924 ( .A(RootIn[25]), .Y(n108), .Z(n109) );
  IVAP U1925 ( .A(RootIn[26]), .Z(n167) );
  IVP U1926 ( .A(n217), .Z(n192) );
  IVP U1927 ( .A(RootIn[27]), .Z(n170) );
  AN2P U1928 ( .A(n170), .B(n167), .Z(n110) );
  IVP U1929 ( .A(RootIn[28]), .Z(n174) );
  IVP U1930 ( .A(RootIn[25]), .Z(n122) );
  IVDAP U1931 ( .A(n110), .Y(n111), .Z(n112) );
  IVP U1932 ( .A(N36), .Z(n161) );
  MUX21H U1933 ( .A(n362), .B(RootIn[25]), .S(RootIn[26]), .Z(n113) );
  B5IP U1934 ( .A(RootIn[29]), .Z(n179) );
  AN2P U1935 ( .A(n389), .B(RootIn[25]), .Z(n114) );
  B4I U1936 ( .A(n179), .Z(n177) );
  AN2P U1937 ( .A(n291), .B(n161), .Z(n115) );
  AN2P U1938 ( .A(n179), .B(n174), .Z(n116) );
  MUX21H U1939 ( .A(n161), .B(n246), .S(RootIn[28]), .Z(n117) );
  AN2P U1940 ( .A(n341), .B(n340), .Z(n118) );
  IVP U1941 ( .A(RootIn[26]), .Z(n166) );
  EO U1943 ( .A(RootIn[26]), .B(n169), .Z(n201) );
  MUX21L U1944 ( .A(n203), .B(n202), .S(RootIn[26]), .Z(n204) );
  MUX21L U1945 ( .A(n201), .B(n200), .S(n157), .Z(n215) );
  ND3 U1946 ( .A(n190), .B(n189), .C(n177), .Z(n194) );
  IV U1947 ( .A(n295), .Z(n369) );
  AO6 U1948 ( .A(n157), .B(RootIn[25]), .C(n204), .Z(n214) );
  IVP U1949 ( .A(RootIn[27]), .Z(n172) );
  ND2P U1950 ( .A(RootIn[27]), .B(RootIn[25]), .Z(n202) );
  B4I U1951 ( .A(RootIn[27]), .Z(n173) );
  EOP U1952 ( .A(n172), .B(n109), .Z(n295) );
  IVAP U1953 ( .A(RootIn[27]), .Z(n121) );
  IVP U1954 ( .A(n173), .Z(n169) );
  ND2P U1955 ( .A(RootIn[26]), .B(n121), .Z(n205) );
  ND2P U1956 ( .A(n163), .B(n167), .Z(n247) );
  ND2P U1957 ( .A(n295), .B(n111), .Z(n345) );
  MUX21LP U1958 ( .A(Term1[39]), .B(N35), .S(n154), .Z(n144) );
  MUX21LP U1959 ( .A(Term1[35]), .B(N31), .S(n153), .Z(n140) );
  MUX21LP U1960 ( .A(Term1[36]), .B(N32), .S(n154), .Z(n142) );
  MUX21LP U1961 ( .A(Term1[38]), .B(N34), .S(n154), .Z(n138) );
  B4IP U1962 ( .A(RootIn[25]), .Z(n123) );
  IVA U1963 ( .A(RootIn[25]), .Z(n165) );
  ND2 U1964 ( .A(n170), .B(n164), .Z(n124) );
  ND6P U1965 ( .A(n198), .B(n197), .C(n196), .D(n195), .E(n194), .F(n193), .Z(
        N18) );
  NR2P U1966 ( .A(n170), .B(RootIn[26]), .Z(n125) );
  B4IP U1967 ( .A(RootIn[27]), .Z(n126) );
  AN2P U1968 ( .A(n172), .B(n165), .Z(n127) );
  B4IP U1969 ( .A(RootIn[27]), .Z(n171) );
  IVA U1970 ( .A(N36), .Z(n159) );
  IVDA U1971 ( .A(n159), .Y(n128) );
  B3I U1972 ( .A(n360), .Z1(n130), .Z2(n129) );
  ND2 U1973 ( .A(n127), .B(n166), .Z(n360) );
  EO U1974 ( .A(RootIn[26]), .B(n120), .Z(n182) );
  MUX41 U1975 ( .D0(n224), .D1(n108), .D2(n223), .D3(n222), .A(n176), .B(n156), 
        .Z(n232) );
  MUX21L U1976 ( .A(n232), .B(n231), .S(RootIn[28]), .Z(N15) );
  OR2P U1977 ( .A(n132), .B(n192), .Z(n297) );
  ND2 U1978 ( .A(n126), .B(n123), .Z(n206) );
  IV U1979 ( .A(n304), .Z(n189) );
  ND2 U1980 ( .A(n131), .B(n386), .Z(n394) );
  MUX21L U1981 ( .A(RootIn[25]), .B(n127), .S(RootIn[26]), .Z(n131) );
  IVP U1982 ( .A(n346), .Z(n136) );
  IVDA U1983 ( .A(n400), .Y(n362) );
  IVDA U1984 ( .A(n280), .Y(n281) );
  IVP U1985 ( .A(N36), .Z(n160) );
  MUX21L U1986 ( .A(n390), .B(RootIn[27]), .S(RootIn[26]), .Z(n305) );
  MUX41 U1987 ( .D0(n284), .D1(n283), .D2(n282), .D3(n281), .A(n176), .B(n128), 
        .Z(n285) );
  MUX31L U1988 ( .D0(n277), .D1(RootIn[27]), .D2(n276), .A(n128), .B(n176), 
        .Z(n286) );
  B4I U1989 ( .A(n179), .Z(n176) );
  IVP U1990 ( .A(n160), .Z(n157) );
  IVP U1991 ( .A(n159), .Z(n158) );
  IVP U1992 ( .A(n161), .Z(n156) );
  ND2 U1993 ( .A(n167), .B(n122), .Z(n387) );
  MUX31L U1994 ( .D0(n114), .D1(n112), .D2(n233), .A(n156), .B(n177), .Z(n234)
         );
  MUX21H U1995 ( .A(n125), .B(n106), .S(RootIn[25]), .Z(n132) );
  ND3 U1996 ( .A(n117), .B(n253), .C(n252), .Z(N12) );
  AO6 U1997 ( .A(n251), .B(n156), .C(n250), .Z(n252) );
  MUX21L U1998 ( .A(n248), .B(n133), .S(n177), .Z(n253) );
  ND2 U1999 ( .A(n329), .B(n179), .Z(n246) );
  AN2P U2000 ( .A(n280), .B(n175), .Z(n133) );
  NR3 U2001 ( .A(n170), .B(n247), .C(RootIn[28]), .Z(n248) );
  MUX21L U2002 ( .A(n339), .B(n107), .S(n173), .Z(n255) );
  AN3 U2003 ( .A(n179), .B(n161), .C(n175), .Z(n134) );
  AO3 U2004 ( .A(n318), .B(n317), .C(n316), .D(n315), .Z(N43) );
  ND2 U2005 ( .A(n176), .B(n174), .Z(n318) );
  AO7 U2006 ( .A(n362), .B(n167), .C(n128), .Z(n317) );
  NR2 U2007 ( .A(n314), .B(n313), .Z(n315) );
  MUX31L U2008 ( .D0(n137), .D1(n118), .D2(n136), .A(n176), .B(RootIn[28]), 
        .Z(n135) );
  MUX21H U2009 ( .A(n127), .B(n114), .S(n128), .Z(n137) );
  MUX21L U2010 ( .A(n308), .B(n307), .S(n176), .Z(n316) );
  NR3 U2011 ( .A(n413), .B(n387), .C(RootIn[27]), .Z(n307) );
  AO6 U2012 ( .A(n306), .B(n305), .C(n304), .Z(n308) );
  NR2 U2013 ( .A(n176), .B(n372), .Z(n373) );
  AO3 U2014 ( .A(n179), .B(n272), .C(n271), .D(n270), .Z(N39) );
  ND2 U2015 ( .A(n175), .B(n110), .Z(n272) );
  NR2 U2016 ( .A(n269), .B(n268), .Z(n270) );
  MUX21L U2017 ( .A(n265), .B(n264), .S(n177), .Z(n271) );
  NR2 U2018 ( .A(n267), .B(n266), .Z(n268) );
  ND2 U2019 ( .A(n128), .B(RootIn[28]), .Z(n267) );
  ND2 U2020 ( .A(n129), .B(n179), .Z(n266) );
  MUX41 U2021 ( .D0(n338), .D1(n337), .D2(n336), .D3(n335), .A(RootIn[28]), 
        .B(n176), .Z(N45) );
  NR2 U2022 ( .A(n130), .B(n263), .Z(n264) );
  ND2 U2023 ( .A(n161), .B(RootIn[28]), .Z(n263) );
  MUX21L U2024 ( .A(n310), .B(n309), .S(n177), .Z(n314) );
  ND3 U2025 ( .A(n394), .B(n128), .C(RootIn[28]), .Z(n309) );
  ND3 U2026 ( .A(n161), .B(RootIn[28]), .C(n371), .Z(n310) );
  MUX21L U2027 ( .A(n312), .B(n311), .S(RootIn[28]), .Z(n313) );
  AO3 U2028 ( .A(n359), .B(n105), .C(n179), .D(n128), .Z(n311) );
  ND2 U2029 ( .A(n115), .B(n176), .Z(n312) );
  AO6 U2030 ( .A(n320), .B(n202), .C(n174), .Z(n269) );
  IVP U2031 ( .A(n155), .Z(n153) );
  IVP U2032 ( .A(n155), .Z(n147) );
  IVP U2033 ( .A(n155), .Z(n148) );
  IVP U2034 ( .A(n155), .Z(n149) );
  IVP U2035 ( .A(n155), .Z(n150) );
  IVP U2036 ( .A(n155), .Z(n151) );
  IVP U2037 ( .A(n155), .Z(n152) );
  IVA U2038 ( .A(N36), .Z(n162) );
  IVP U2039 ( .A(RootIn[26]), .Z(n168) );
  MUX21L U2040 ( .A(RootIn[25]), .B(n167), .S(RootIn[27]), .Z(n190) );
  IVP U2041 ( .A(RootIn[29]), .Z(n178) );
  ND2 U2042 ( .A(n169), .B(n108), .Z(n400) );
  NR2 U2043 ( .A(n387), .B(RootIn[27]), .Z(n251) );
  AO5 U2044 ( .A(n91), .B(n90), .C(n92), .Z(n97) );
  EN U2045 ( .A(Term11[39]), .B(n94), .Z(N73) );
  AO5 U2046 ( .A(n415), .B(Term11[38]), .C(Term21[19]), .Z(n94) );
  IVP U2047 ( .A(n95), .Z(n415) );
  AO4 U2048 ( .A(n96), .B(Term21[18]), .C(n97), .D(Term11[37]), .Z(n95) );
  NR2 U2049 ( .A(n262), .B(n304), .Z(n265) );
  MUX21L U2050 ( .A(RootIn[25]), .B(RootIn[27]), .S(RootIn[26]), .Z(n262) );
  MUX41 U2051 ( .D0(n301), .D1(n300), .D2(n299), .D3(n298), .A(n177), .B(n128), 
        .Z(n302) );
  MUX31L U2052 ( .D0(n297), .D1(RootIn[25]), .D2(n296), .A(n128), .B(n177), 
        .Z(n303) );
  ND2 U2053 ( .A(Term11[36]), .B(FractionBit[13]), .Z(n101) );
  EN U2054 ( .A(n97), .B(n102), .Z(N71) );
  EN U2055 ( .A(Term11[37]), .B(Term21[18]), .Z(n102) );
  EO U2056 ( .A(n98), .B(n99), .Z(N72) );
  EN U2057 ( .A(Term11[38]), .B(Term21[19]), .Z(n99) );
  AO5 U2058 ( .A(Term11[37]), .B(n100), .C(Term21[18]), .Z(n98) );
  AO2 U2059 ( .A(n101), .B(n92), .C(n90), .D(n91), .Z(n100) );
  EO U2060 ( .A(FractionBit[13]), .B(n103), .Z(N70) );
  EO U2061 ( .A(Term21[17]), .B(Term11[36]), .Z(n103) );
  IVP U2062 ( .A(n414), .Z(n155) );
  IVP U2063 ( .A(reset), .Z(n414) );
  OR3 U2064 ( .A(n212), .B(n211), .C(n210), .Z(n213) );
  ND2 U2065 ( .A(n126), .B(n168), .Z(n408) );
  EON1 U2066 ( .A(n209), .B(n249), .C(n208), .D(n207), .Z(n210) );
  ND2 U2067 ( .A(RootIn[26]), .B(n105), .Z(n146) );
  MUX21L U2068 ( .A(n205), .B(n106), .S(RootIn[25]), .Z(n209) );
  IVP U2069 ( .A(n249), .Z(n250) );
  OR2P U2070 ( .A(n162), .B(RootIn[29]), .Z(n249) );
  AN2 U2071 ( .A(n115), .B(RootIn[28]), .Z(n236) );
  ND4 U2072 ( .A(RootIn[28]), .B(n161), .C(n176), .D(n180), .Z(n197) );
  AO1 U2073 ( .A(n156), .B(n129), .C(n192), .D(n390), .Z(n233) );
  ND4 U2074 ( .A(n247), .B(n161), .C(n172), .D(n179), .Z(n198) );
  ND5 U2075 ( .A(n166), .B(n124), .C(RootIn[28]), .D(n178), .E(n158), .Z(n196)
         );
  AN2 U2076 ( .A(n158), .B(n178), .Z(n191) );
  ND2 U2077 ( .A(n178), .B(n159), .Z(n185) );
  AO7 U2078 ( .A(n109), .B(n169), .C(RootIn[26]), .Z(n180) );
  IV U2079 ( .A(n155), .Z(n154) );
  AN2P U2080 ( .A(n408), .B(RootIn[29]), .Z(n183) );
  AO3P U2081 ( .A(n192), .B(n107), .C(n175), .D(n191), .Z(n193) );
  ND2 U2082 ( .A(RootIn[26]), .B(n109), .Z(n199) );
  ND2 U2083 ( .A(n169), .B(n199), .Z(n200) );
  ND2 U2084 ( .A(RootIn[25]), .B(n105), .Z(n203) );
  AN3 U2085 ( .A(n247), .B(n170), .C(RootIn[29]), .Z(n212) );
  NR5 U2086 ( .A(n178), .B(n160), .C(n172), .D(RootIn[26]), .E(n122), .Z(n211)
         );
  AO1P U2087 ( .A(RootIn[26]), .B(n171), .C(N36), .D(RootIn[29]), .Z(n208) );
  ND2 U2088 ( .A(n206), .B(n167), .Z(n207) );
  MUX31LP U2089 ( .D0(n215), .D1(n214), .D2(n213), .A(n177), .B(RootIn[28]), 
        .Z(N17) );
  ND2 U2090 ( .A(RootIn[25]), .B(n106), .Z(n348) );
  MUX21L U2091 ( .A(n348), .B(RootIn[25]), .S(RootIn[26]), .Z(n220) );
  ND2 U2092 ( .A(n172), .B(n123), .Z(n388) );
  IVA U2093 ( .A(n202), .Z(n216) );
  MUX21L U2094 ( .A(n216), .B(n122), .S(RootIn[26]), .Z(n218) );
  ND3 U2095 ( .A(n218), .B(n217), .C(n388), .Z(n219) );
  EO U2096 ( .A(n166), .B(RootIn[25]), .Z(n352) );
  IVA U2097 ( .A(n352), .Z(n350) );
  ND2 U2098 ( .A(n348), .B(n166), .Z(n405) );
  MUX81P U2099 ( .D0(n192), .D1(n220), .D2(n130), .D3(n345), .D4(n295), .D5(
        n219), .D6(n350), .D7(n405), .A(RootIn[28]), .B(n177), .C(n156), .Z(
        N16) );
  MUX21L U2100 ( .A(n173), .B(RootIn[26]), .S(RootIn[25]), .Z(n240) );
  IVA U2101 ( .A(n240), .Z(n224) );
  ND2 U2102 ( .A(RootIn[26]), .B(n122), .Z(n349) );
  MUX21L U2103 ( .A(n166), .B(n107), .S(RootIn[27]), .Z(n221) );
  ND2 U2104 ( .A(n221), .B(n247), .Z(n290) );
  IVA U2105 ( .A(n290), .Z(n223) );
  IVA U2106 ( .A(n297), .Z(n222) );
  MUX21L U2107 ( .A(RootIn[26]), .B(n339), .S(RootIn[27]), .Z(n332) );
  EO U2108 ( .A(n105), .B(RootIn[26]), .Z(n329) );
  ND2 U2109 ( .A(n329), .B(n400), .Z(n225) );
  ND2 U2110 ( .A(n225), .B(n160), .Z(n226) );
  ND2 U2111 ( .A(n332), .B(n226), .Z(n230) );
  IVA U2112 ( .A(n394), .Z(n228) );
  IVA U2113 ( .A(n329), .Z(n389) );
  ND2 U2114 ( .A(n156), .B(n389), .Z(n227) );
  ND2 U2115 ( .A(n228), .B(n227), .Z(n229) );
  MUX21L U2116 ( .A(n230), .B(n229), .S(n177), .Z(n231) );
  MUX21L U2117 ( .A(RootIn[25]), .B(n167), .S(RootIn[27]), .Z(n354) );
  ND2 U2118 ( .A(RootIn[27]), .B(n387), .Z(n280) );
  IVA U2119 ( .A(n348), .Z(n390) );
  ND2 U2120 ( .A(n388), .B(n166), .Z(n291) );
  AN3 U2121 ( .A(n156), .B(n129), .C(RootIn[28]), .Z(n235) );
  MUX21L U2122 ( .A(n236), .B(n235), .S(n176), .Z(n245) );
  MUX21L U2123 ( .A(n112), .B(RootIn[27]), .S(RootIn[25]), .Z(n237) );
  ND2 U2124 ( .A(RootIn[27]), .B(RootIn[26]), .Z(n320) );
  ND2 U2125 ( .A(n237), .B(n320), .Z(n279) );
  AN3 U2126 ( .A(n279), .B(n174), .C(n176), .Z(n239) );
  AN3 U2127 ( .A(n167), .B(n179), .C(n105), .Z(n238) );
  MUX21L U2128 ( .A(n239), .B(n238), .S(n156), .Z(n244) );
  ND3 U2129 ( .A(n240), .B(n174), .C(n179), .Z(n243) );
  AN3 U2130 ( .A(n177), .B(n106), .C(n339), .Z(n241) );
  MUX21L U2131 ( .A(n241), .B(n116), .S(n156), .Z(n242) );
  ND4 U2132 ( .A(n245), .B(n244), .C(n243), .D(n242), .Z(N13) );
  ND2 U2133 ( .A(RootIn[25]), .B(n166), .Z(n347) );
  IVA U2134 ( .A(n347), .Z(n254) );
  ND2 U2135 ( .A(n254), .B(n172), .Z(n399) );
  ND3 U2136 ( .A(n255), .B(n399), .C(n174), .Z(n256) );
  ND3 U2137 ( .A(n320), .B(n179), .C(n256), .Z(n257) );
  ND2 U2138 ( .A(n161), .B(n257), .Z(N11) );
  ND2 U2139 ( .A(n388), .B(n146), .Z(n260) );
  ND2 U2140 ( .A(n176), .B(n161), .Z(n412) );
  IVA U2141 ( .A(n412), .Z(n259) );
  ND2 U2142 ( .A(RootIn[28]), .B(n161), .Z(n413) );
  IVA U2143 ( .A(n413), .Z(n258) );
  AO1P U2144 ( .A(n260), .B(n161), .C(n259), .D(n258), .Z(n261) );
  IVA U2145 ( .A(n261), .Z(N10) );
  AN3 U2146 ( .A(n111), .B(n161), .C(n116), .Z(N9) );
  AN3 U2147 ( .A(n110), .B(RootIn[25]), .C(n134), .Z(N8) );
  AN2P U2148 ( .A(n134), .B(n130), .Z(N7) );
  ND2 U2149 ( .A(n295), .B(n389), .Z(n277) );
  MUX21L U2150 ( .A(RootIn[27]), .B(n202), .S(RootIn[26]), .Z(n374) );
  IVA U2151 ( .A(n374), .Z(n275) );
  ND2 U2152 ( .A(n202), .B(n389), .Z(n273) );
  ND2 U2153 ( .A(n273), .B(n161), .Z(n274) );
  ND2 U2154 ( .A(n275), .B(n274), .Z(n276) );
  MUX21L U2155 ( .A(n362), .B(n173), .S(RootIn[26]), .Z(n278) );
  ND2 U2156 ( .A(RootIn[26]), .B(RootIn[25]), .Z(n401) );
  ND2 U2157 ( .A(n278), .B(n401), .Z(n289) );
  IVA U2158 ( .A(n289), .Z(n284) );
  ND2 U2159 ( .A(n387), .B(n106), .Z(n404) );
  IVA U2160 ( .A(n404), .Z(n283) );
  IVA U2161 ( .A(n279), .Z(n282) );
  MUX21L U2162 ( .A(n286), .B(n285), .S(RootIn[28]), .Z(N40) );
  MUX21L U2163 ( .A(RootIn[26]), .B(n105), .S(RootIn[25]), .Z(n293) );
  IVA U2164 ( .A(n320), .Z(n287) );
  MUX21L U2165 ( .A(n125), .B(n287), .S(RootIn[25]), .Z(n288) );
  ND2 U2166 ( .A(n288), .B(n399), .Z(n292) );
  MUX21L U2167 ( .A(RootIn[26]), .B(n146), .S(RootIn[25]), .Z(n395) );
  MUX81P U2168 ( .D0(n293), .D1(n369), .D2(n292), .D3(n291), .D4(RootIn[26]), 
        .D5(n395), .D6(n290), .D7(n289), .A(RootIn[28]), .B(n176), .C(n128), 
        .Z(N41) );
  ND2 U2169 ( .A(n345), .B(n161), .Z(n294) );
  ND2 U2170 ( .A(n295), .B(n294), .Z(n296) );
  ND2 U2171 ( .A(n386), .B(n400), .Z(n342) );
  IVA U2172 ( .A(n342), .Z(n301) );
  ND2 U2173 ( .A(n111), .B(n108), .Z(n322) );
  IVA U2174 ( .A(n322), .Z(n300) );
  AN2P U2175 ( .A(RootIn[25]), .B(n320), .Z(n299) );
  IVA U2176 ( .A(n345), .Z(n298) );
  MUX21L U2177 ( .A(n303), .B(n302), .S(RootIn[28]), .Z(N42) );
  AN2P U2178 ( .A(n400), .B(n349), .Z(n306) );
  ND2 U2179 ( .A(n369), .B(RootIn[26]), .Z(n371) );
  ND2 U2180 ( .A(n349), .B(n170), .Z(n324) );
  MUX21L U2181 ( .A(RootIn[26]), .B(RootIn[27]), .S(RootIn[25]), .Z(n323) );
  ND2 U2182 ( .A(n350), .B(n172), .Z(n321) );
  ND2 U2183 ( .A(n369), .B(n386), .Z(n319) );
  MUX81P U2184 ( .D0(n324), .D1(n323), .D2(n322), .D3(n321), .D4(n320), .D5(
        n371), .D6(n319), .D7(n369), .A(RootIn[28]), .B(n177), .C(n128), .Z(
        N44) );
  ND2 U2185 ( .A(n202), .B(n386), .Z(n326) );
  ND2 U2186 ( .A(RootIn[27]), .B(n349), .Z(n325) );
  MUX21H U2187 ( .A(n326), .B(n325), .S(n128), .Z(n338) );
  ND2 U2188 ( .A(n388), .B(n387), .Z(n328) );
  ND2 U2189 ( .A(n389), .B(n400), .Z(n327) );
  MUX21H U2190 ( .A(n328), .B(n327), .S(n128), .Z(n337) );
  ND2 U2191 ( .A(n329), .B(RootIn[25]), .Z(n330) );
  ND2 U2192 ( .A(n330), .B(n161), .Z(n331) );
  ND2 U2193 ( .A(n332), .B(n331), .Z(n336) );
  ND2 U2194 ( .A(n192), .B(RootIn[25]), .Z(n333) );
  ND2 U2195 ( .A(n333), .B(n161), .Z(n334) );
  ND2 U2196 ( .A(n106), .B(n334), .Z(n335) );
  MUX21L U2197 ( .A(RootIn[25]), .B(n339), .S(RootIn[27]), .Z(n341) );
  ND2 U2198 ( .A(n349), .B(n161), .Z(n340) );
  ND2 U2199 ( .A(n369), .B(n167), .Z(n344) );
  ND2 U2200 ( .A(n350), .B(n386), .Z(n343) );
  ND2 U2201 ( .A(n348), .B(n347), .Z(n357) );
  ND2 U2202 ( .A(n386), .B(n108), .Z(n356) );
  ND2 U2203 ( .A(n349), .B(n400), .Z(n355) );
  ND2 U2204 ( .A(n350), .B(n111), .Z(n353) );
  IVA U2205 ( .A(n401), .Z(n359) );
  MUX21L U2206 ( .A(n166), .B(n359), .S(RootIn[27]), .Z(n351) );
  ND2 U2207 ( .A(n351), .B(n387), .Z(n379) );
  ND2 U2208 ( .A(RootIn[26]), .B(n388), .Z(n397) );
  MUX81P U2209 ( .D0(n357), .D1(n356), .D2(n355), .D3(n354), .D4(n353), .D5(
        n352), .D6(n379), .D7(n397), .A(RootIn[28]), .B(n177), .C(n128), .Z(
        N47) );
  MUX21L U2210 ( .A(n217), .B(n173), .S(RootIn[25]), .Z(n368) );
  MUX21L U2211 ( .A(RootIn[25]), .B(RootIn[26]), .S(RootIn[27]), .Z(n367) );
  ND2 U2212 ( .A(n202), .B(n401), .Z(n366) );
  MUX21L U2213 ( .A(n108), .B(n359), .S(RootIn[27]), .Z(n358) );
  ND2 U2214 ( .A(n358), .B(n387), .Z(n365) );
  MUX21L U2215 ( .A(n111), .B(n386), .S(RootIn[25]), .Z(n364) );
  MUX21L U2216 ( .A(n359), .B(n107), .S(RootIn[27]), .Z(n361) );
  ND2 U2217 ( .A(n361), .B(n129), .Z(n363) );
  MUX81P U2218 ( .D0(n368), .D1(n367), .D2(n366), .D3(n365), .D4(n364), .D5(
        n363), .D6(n107), .D7(n113), .A(RootIn[28]), .B(n176), .C(n128), .Z(
        N48) );
  ND2 U2219 ( .A(n369), .B(n389), .Z(n370) );
  MUX21L U2220 ( .A(n371), .B(n370), .S(n128), .Z(n372) );
  AO1P U2221 ( .A(n374), .B(n161), .C(n373), .D(n130), .Z(n385) );
  MUX21L U2222 ( .A(n112), .B(n192), .S(RootIn[25]), .Z(n377) );
  MUX21L U2223 ( .A(n108), .B(n400), .S(RootIn[26]), .Z(n375) );
  ND2 U2224 ( .A(n375), .B(n161), .Z(n376) );
  ND2 U2225 ( .A(n377), .B(n376), .Z(n383) );
  MUX21L U2226 ( .A(n127), .B(RootIn[27]), .S(RootIn[26]), .Z(n378) );
  AN3 U2227 ( .A(n378), .B(n202), .C(n401), .Z(n381) );
  IVA U2228 ( .A(n379), .Z(n380) );
  MUX21L U2229 ( .A(n381), .B(n380), .S(n128), .Z(n382) );
  MUX21L U2230 ( .A(n383), .B(n382), .S(n177), .Z(n384) );
  MUX21L U2231 ( .A(n385), .B(n384), .S(RootIn[28]), .Z(N49) );
  ND3 U2232 ( .A(n400), .B(n387), .C(n386), .Z(n398) );
  MUX21L U2233 ( .A(n388), .B(n126), .S(RootIn[26]), .Z(n396) );
  ND2 U2234 ( .A(n389), .B(n388), .Z(n393) );
  MUX21L U2235 ( .A(n390), .B(n108), .S(RootIn[26]), .Z(n391) );
  ND2 U2236 ( .A(n391), .B(n400), .Z(n392) );
  MUX81P U2237 ( .D0(n398), .D1(n397), .D2(n396), .D3(n395), .D4(n394), .D5(
        n393), .D6(n392), .D7(RootIn[27]), .A(RootIn[28]), .B(n176), .C(n128), 
        .Z(N50) );
  MUX21L U2238 ( .A(n108), .B(RootIn[26]), .S(RootIn[27]), .Z(n407) );
  IVA U2239 ( .A(n399), .Z(n406) );
  MUX21L U2240 ( .A(RootIn[27]), .B(n400), .S(RootIn[26]), .Z(n403) );
  ND2 U2241 ( .A(n401), .B(n217), .Z(n402) );
  MUX81P U2242 ( .D0(n407), .D1(RootIn[26]), .D2(n406), .D3(n405), .D4(n404), 
        .D5(n403), .D6(n402), .D7(n113), .A(RootIn[28]), .B(n177), .C(n128), 
        .Z(N51) );
  ND2 U2243 ( .A(n177), .B(n111), .Z(n411) );
  AN2P U2244 ( .A(n111), .B(n161), .Z(n409) );
  MUX21L U2245 ( .A(n409), .B(n177), .S(RootIn[28]), .Z(n410) );
  ND2 U2246 ( .A(n411), .B(n410), .Z(N38) );
  ND2 U2247 ( .A(n413), .B(n412), .Z(N37) );
endmodule

