
module LOG_POLY_DW01_add_4 ( A, B, CI, SUM, CO );
  input [67:0] A;
  input [67:0] B;
  output [67:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230;

  IVP U2 ( .A(n55), .Z(n2) );
  IVP U3 ( .A(n160), .Z(n24) );
  IVP U4 ( .A(n59), .Z(n3) );
  IVP U5 ( .A(n100), .Z(n11) );
  IVP U6 ( .A(n64), .Z(n5) );
  IVP U7 ( .A(n54), .Z(n1) );
  IVP U8 ( .A(n113), .Z(n16) );
  IVP U9 ( .A(n106), .Z(n13) );
  IVP U10 ( .A(n109), .Z(n15) );
  IVP U11 ( .A(n121), .Z(n21) );
  IVP U12 ( .A(n125), .Z(n18) );
  IVP U13 ( .A(n180), .Z(n31) );
  IVP U14 ( .A(n171), .Z(n28) );
  IVP U15 ( .A(n143), .Z(n25) );
  IVP U16 ( .A(n122), .Z(n23) );
  IVP U17 ( .A(n176), .Z(n30) );
  IVP U18 ( .A(n148), .Z(n27) );
  IVP U19 ( .A(n194), .Z(n36) );
  IVP U20 ( .A(n201), .Z(n35) );
  IVP U21 ( .A(n195), .Z(n33) );
  IVP U22 ( .A(n191), .Z(n34) );
  IVP U23 ( .A(n203), .Z(n37) );
  IVP U24 ( .A(n179), .Z(n29) );
  IVP U25 ( .A(n166), .Z(n26) );
  IVP U26 ( .A(n130), .Z(n19) );
  IVP U27 ( .A(n123), .Z(n20) );
  IVP U28 ( .A(n112), .Z(n14) );
  IVP U29 ( .A(n85), .Z(n7) );
  IVP U30 ( .A(n97), .Z(n9) );
  IVP U31 ( .A(n91), .Z(n10) );
  IVP U32 ( .A(n101), .Z(n12) );
  IVP U33 ( .A(n86), .Z(n8) );
  IVP U34 ( .A(n82), .Z(n6) );
  IVP U35 ( .A(n177), .Z(n32) );
  IVP U36 ( .A(n110), .Z(n17) );
  IVP U37 ( .A(n77), .Z(n4) );
  IVP U38 ( .A(n132), .Z(n22) );
  IVP U39 ( .A(n225), .Z(n48) );
  IVP U40 ( .A(n222), .Z(n45) );
  IVP U41 ( .A(n224), .Z(n46) );
  IVP U42 ( .A(n216), .Z(n43) );
  IVP U43 ( .A(A[22]), .Z(n49) );
  IVP U44 ( .A(n205), .Z(n38) );
  IVP U45 ( .A(n154), .Z(n39) );
  IVP U46 ( .A(n211), .Z(n40) );
  IVP U47 ( .A(A[32]), .Z(n41) );
  IVP U48 ( .A(n219), .Z(n44) );
  IVP U49 ( .A(A[24]), .Z(n47) );
  IVP U50 ( .A(n229), .Z(n50) );
  IVP U51 ( .A(A[29]), .Z(n42) );
  ND2 U52 ( .A(A[21]), .B(B[21]), .Z(n229) );
  EO U53 ( .A(n51), .B(n52), .Z(SUM[65]) );
  EO U54 ( .A(B[65]), .B(A[65]), .Z(n52) );
  AO7 U55 ( .A(n53), .B(n2), .C(n54), .Z(n51) );
  EO U56 ( .A(n55), .B(n56), .Z(SUM[64]) );
  NR2 U57 ( .A(n1), .B(n53), .Z(n56) );
  NR2 U58 ( .A(B[64]), .B(A[64]), .Z(n53) );
  ND2 U59 ( .A(B[64]), .B(A[64]), .Z(n54) );
  AO7 U60 ( .A(n57), .B(n58), .C(n59), .Z(n55) );
  AO6 U61 ( .A(n60), .B(n61), .C(n4), .Z(n58) );
  AO7 U62 ( .A(n62), .B(n63), .C(n64), .Z(n60) );
  AO6 U63 ( .A(n65), .B(n6), .C(n66), .Z(n63) );
  AO7 U64 ( .A(n67), .B(n68), .C(n7), .Z(n65) );
  AO1 U65 ( .A(n69), .B(n70), .C(n71), .D(n72), .Z(n67) );
  AN2 U66 ( .A(n73), .B(n70), .Z(n72) );
  EN U67 ( .A(n74), .B(n75), .Z(SUM[63]) );
  NR2 U68 ( .A(n3), .B(n57), .Z(n75) );
  NR2 U69 ( .A(B[63]), .B(A[63]), .Z(n57) );
  ND2 U70 ( .A(B[63]), .B(A[63]), .Z(n59) );
  AO6 U71 ( .A(n61), .B(n76), .C(n4), .Z(n74) );
  EN U72 ( .A(n78), .B(n76), .Z(SUM[62]) );
  AO7 U73 ( .A(n62), .B(n79), .C(n64), .Z(n76) );
  ND2 U74 ( .A(n61), .B(n77), .Z(n78) );
  ND2 U75 ( .A(B[62]), .B(A[62]), .Z(n77) );
  OR2 U76 ( .A(B[62]), .B(A[62]), .Z(n61) );
  EN U77 ( .A(n79), .B(n80), .Z(SUM[61]) );
  NR2 U78 ( .A(n5), .B(n62), .Z(n80) );
  NR2 U79 ( .A(B[61]), .B(A[61]), .Z(n62) );
  ND2 U80 ( .A(B[61]), .B(A[61]), .Z(n64) );
  AO6 U81 ( .A(n6), .B(n81), .C(n66), .Z(n79) );
  EO U82 ( .A(n81), .B(n83), .Z(SUM[60]) );
  NR2 U83 ( .A(n66), .B(n82), .Z(n83) );
  NR2 U84 ( .A(B[60]), .B(A[60]), .Z(n82) );
  AN2 U85 ( .A(B[60]), .B(A[60]), .Z(n66) );
  AO7 U86 ( .A(n84), .B(n68), .C(n7), .Z(n81) );
  AO7 U87 ( .A(n86), .B(n87), .C(n88), .Z(n85) );
  AO6 U88 ( .A(n89), .B(n9), .C(n90), .Z(n87) );
  AO7 U89 ( .A(n91), .B(n92), .C(n93), .Z(n89) );
  ND4 U90 ( .A(n8), .B(n9), .C(n10), .D(n12), .Z(n68) );
  EO U91 ( .A(n94), .B(n95), .Z(SUM[59]) );
  AO6 U92 ( .A(n96), .B(n9), .C(n90), .Z(n95) );
  ND2 U93 ( .A(n8), .B(n88), .Z(n94) );
  ND2 U94 ( .A(B[59]), .B(A[59]), .Z(n88) );
  NR2 U95 ( .A(B[59]), .B(A[59]), .Z(n86) );
  EO U96 ( .A(n96), .B(n98), .Z(SUM[58]) );
  NR2 U97 ( .A(n90), .B(n97), .Z(n98) );
  NR2 U98 ( .A(B[58]), .B(A[58]), .Z(n97) );
  AN2 U99 ( .A(B[58]), .B(A[58]), .Z(n90) );
  AO7 U100 ( .A(n91), .B(n11), .C(n93), .Z(n96) );
  EO U101 ( .A(n11), .B(n99), .Z(SUM[57]) );
  ND2 U102 ( .A(n93), .B(n10), .Z(n99) );
  NR2 U103 ( .A(B[57]), .B(A[57]), .Z(n91) );
  ND2 U104 ( .A(B[57]), .B(A[57]), .Z(n93) );
  AO7 U105 ( .A(n101), .B(n84), .C(n92), .Z(n100) );
  EO U106 ( .A(n102), .B(n84), .Z(SUM[56]) );
  AO6 U107 ( .A(n103), .B(n70), .C(n71), .Z(n84) );
  AO7 U108 ( .A(n104), .B(n105), .C(n106), .Z(n71) );
  AO6 U109 ( .A(n107), .B(n14), .C(n108), .Z(n105) );
  AO7 U110 ( .A(n109), .B(n110), .C(n111), .Z(n107) );
  NR4 U111 ( .A(n104), .B(n112), .C(n109), .D(n113), .Z(n70) );
  ND2 U112 ( .A(n12), .B(n92), .Z(n102) );
  ND2 U113 ( .A(B[56]), .B(A[56]), .Z(n92) );
  NR2 U114 ( .A(B[56]), .B(A[56]), .Z(n101) );
  EN U115 ( .A(n114), .B(n115), .Z(SUM[55]) );
  NR2 U116 ( .A(n13), .B(n104), .Z(n115) );
  NR2 U117 ( .A(B[55]), .B(A[55]), .Z(n104) );
  ND2 U118 ( .A(B[55]), .B(A[55]), .Z(n106) );
  AO6 U119 ( .A(n14), .B(n116), .C(n108), .Z(n114) );
  EO U120 ( .A(n116), .B(n117), .Z(SUM[54]) );
  NR2 U121 ( .A(n108), .B(n112), .Z(n117) );
  NR2 U122 ( .A(B[54]), .B(A[54]), .Z(n112) );
  AN2 U123 ( .A(B[54]), .B(A[54]), .Z(n108) );
  AO7 U124 ( .A(n109), .B(n118), .C(n111), .Z(n116) );
  EO U125 ( .A(n119), .B(n118), .Z(SUM[53]) );
  AO6 U126 ( .A(n16), .B(n103), .C(n17), .Z(n118) );
  ND2 U127 ( .A(n15), .B(n111), .Z(n119) );
  ND2 U128 ( .A(B[53]), .B(A[53]), .Z(n111) );
  NR2 U129 ( .A(B[53]), .B(A[53]), .Z(n109) );
  EO U130 ( .A(n103), .B(n120), .Z(SUM[52]) );
  NR2 U131 ( .A(n17), .B(n113), .Z(n120) );
  NR2 U132 ( .A(B[52]), .B(A[52]), .Z(n113) );
  ND2 U133 ( .A(B[52]), .B(A[52]), .Z(n110) );
  OR2 U134 ( .A(n73), .B(n69), .Z(n103) );
  NR4 U135 ( .A(n121), .B(n122), .C(n123), .D(n124), .Z(n69) );
  OR2 U136 ( .A(n125), .B(n126), .Z(n124) );
  AO7 U137 ( .A(n125), .B(n127), .C(n128), .Z(n73) );
  AO6 U138 ( .A(n129), .B(n20), .C(n19), .Z(n127) );
  AO7 U139 ( .A(n121), .B(n131), .C(n132), .Z(n129) );
  EN U140 ( .A(n133), .B(n134), .Z(SUM[51]) );
  ND2 U141 ( .A(n128), .B(n18), .Z(n134) );
  NR2 U142 ( .A(B[51]), .B(A[51]), .Z(n125) );
  ND2 U143 ( .A(B[51]), .B(A[51]), .Z(n128) );
  AO7 U144 ( .A(n123), .B(n135), .C(n130), .Z(n133) );
  EO U145 ( .A(n136), .B(n135), .Z(SUM[50]) );
  AO6 U146 ( .A(n21), .B(n137), .C(n22), .Z(n135) );
  ND2 U147 ( .A(n20), .B(n130), .Z(n136) );
  ND2 U148 ( .A(B[50]), .B(A[50]), .Z(n130) );
  NR2 U149 ( .A(B[50]), .B(A[50]), .Z(n123) );
  EO U150 ( .A(n137), .B(n138), .Z(SUM[49]) );
  NR2 U151 ( .A(n22), .B(n121), .Z(n138) );
  NR2 U152 ( .A(B[49]), .B(A[49]), .Z(n121) );
  ND2 U153 ( .A(B[49]), .B(A[49]), .Z(n132) );
  AO7 U154 ( .A(n122), .B(n126), .C(n131), .Z(n137) );
  EO U155 ( .A(n139), .B(n126), .Z(SUM[48]) );
  AO6 U156 ( .A(n24), .B(n140), .C(n141), .Z(n126) );
  AO7 U157 ( .A(n142), .B(n143), .C(n144), .Z(n140) );
  AO6 U158 ( .A(n26), .B(n145), .C(n146), .Z(n142) );
  AO3 U159 ( .A(n147), .B(n148), .C(n149), .D(n150), .Z(n145) );
  OR4 U160 ( .A(n151), .B(n152), .C(n153), .D(n148), .Z(n149) );
  ND2 U161 ( .A(n154), .B(n155), .Z(n151) );
  AO6 U162 ( .A(n156), .B(n155), .C(n157), .Z(n147) );
  AO7 U163 ( .A(n152), .B(n158), .C(n159), .Z(n156) );
  ND2 U164 ( .A(n23), .B(n131), .Z(n139) );
  ND2 U165 ( .A(B[48]), .B(A[48]), .Z(n131) );
  NR2 U166 ( .A(B[48]), .B(A[48]), .Z(n122) );
  EO U167 ( .A(n161), .B(n162), .Z(SUM[47]) );
  NR2 U168 ( .A(n141), .B(n160), .Z(n162) );
  NR2 U169 ( .A(B[47]), .B(A[47]), .Z(n160) );
  AN2 U170 ( .A(B[47]), .B(A[47]), .Z(n141) );
  AO7 U171 ( .A(n143), .B(n163), .C(n144), .Z(n161) );
  EO U172 ( .A(n164), .B(n163), .Z(SUM[46]) );
  AO6 U173 ( .A(n26), .B(n165), .C(n146), .Z(n163) );
  ND2 U174 ( .A(n25), .B(n144), .Z(n164) );
  ND2 U175 ( .A(B[46]), .B(A[46]), .Z(n144) );
  NR2 U176 ( .A(B[46]), .B(A[46]), .Z(n143) );
  EO U177 ( .A(n165), .B(n167), .Z(SUM[45]) );
  NR2 U178 ( .A(n146), .B(n166), .Z(n167) );
  NR2 U179 ( .A(B[45]), .B(A[45]), .Z(n166) );
  AN2 U180 ( .A(B[45]), .B(A[45]), .Z(n146) );
  AO7 U181 ( .A(n148), .B(n168), .C(n150), .Z(n165) );
  EO U182 ( .A(n169), .B(n168), .Z(SUM[44]) );
  AO6 U183 ( .A(n170), .B(n155), .C(n157), .Z(n168) );
  AO7 U184 ( .A(n171), .B(n172), .C(n173), .Z(n157) );
  AO6 U185 ( .A(n174), .B(n29), .C(n175), .Z(n172) );
  AO7 U186 ( .A(n176), .B(n177), .C(n178), .Z(n174) );
  NR4 U187 ( .A(n171), .B(n179), .C(n176), .D(n180), .Z(n155) );
  ND2 U188 ( .A(n27), .B(n150), .Z(n169) );
  ND2 U189 ( .A(B[44]), .B(A[44]), .Z(n150) );
  NR2 U190 ( .A(B[44]), .B(A[44]), .Z(n148) );
  EO U191 ( .A(n181), .B(n182), .Z(SUM[43]) );
  AO6 U192 ( .A(n183), .B(n29), .C(n175), .Z(n182) );
  ND2 U193 ( .A(n28), .B(n173), .Z(n181) );
  ND2 U194 ( .A(B[43]), .B(A[43]), .Z(n173) );
  NR2 U195 ( .A(B[43]), .B(A[43]), .Z(n171) );
  EO U196 ( .A(n183), .B(n184), .Z(SUM[42]) );
  NR2 U197 ( .A(n175), .B(n179), .Z(n184) );
  NR2 U198 ( .A(B[42]), .B(A[42]), .Z(n179) );
  AN2 U199 ( .A(B[42]), .B(A[42]), .Z(n175) );
  AO7 U200 ( .A(n176), .B(n185), .C(n178), .Z(n183) );
  EO U201 ( .A(n186), .B(n185), .Z(SUM[41]) );
  AO6 U202 ( .A(n31), .B(n170), .C(n32), .Z(n185) );
  ND2 U203 ( .A(n30), .B(n178), .Z(n186) );
  ND2 U204 ( .A(B[41]), .B(A[41]), .Z(n178) );
  NR2 U205 ( .A(B[41]), .B(A[41]), .Z(n176) );
  EO U206 ( .A(n170), .B(n187), .Z(SUM[40]) );
  NR2 U207 ( .A(n32), .B(n180), .Z(n187) );
  NR2 U208 ( .A(B[40]), .B(A[40]), .Z(n180) );
  ND2 U209 ( .A(B[40]), .B(A[40]), .Z(n177) );
  AO7 U210 ( .A(n38), .B(n152), .C(n159), .Z(n170) );
  AO6 U211 ( .A(n33), .B(n188), .C(n189), .Z(n159) );
  AO7 U212 ( .A(n190), .B(n191), .C(n192), .Z(n188) );
  AO6 U213 ( .A(n35), .B(n36), .C(n193), .Z(n190) );
  ND4 U214 ( .A(n33), .B(n34), .C(n35), .D(n37), .Z(n152) );
  EO U215 ( .A(n196), .B(n197), .Z(SUM[39]) );
  NR2 U216 ( .A(n189), .B(n195), .Z(n197) );
  NR2 U217 ( .A(B[39]), .B(A[39]), .Z(n195) );
  AN2 U218 ( .A(B[39]), .B(A[39]), .Z(n189) );
  AO7 U219 ( .A(n191), .B(n198), .C(n192), .Z(n196) );
  EO U220 ( .A(n199), .B(n198), .Z(SUM[38]) );
  AO6 U221 ( .A(n35), .B(n200), .C(n193), .Z(n198) );
  ND2 U222 ( .A(n34), .B(n192), .Z(n199) );
  ND2 U223 ( .A(B[38]), .B(A[38]), .Z(n192) );
  NR2 U224 ( .A(B[38]), .B(A[38]), .Z(n191) );
  EO U225 ( .A(n200), .B(n202), .Z(SUM[37]) );
  NR2 U226 ( .A(n193), .B(n201), .Z(n202) );
  NR2 U227 ( .A(B[37]), .B(A[37]), .Z(n201) );
  AN2 U228 ( .A(B[37]), .B(A[37]), .Z(n193) );
  AO7 U229 ( .A(n203), .B(n38), .C(n194), .Z(n200) );
  EO U230 ( .A(n204), .B(n38), .Z(SUM[36]) );
  AO7 U231 ( .A(n153), .B(n39), .C(n158), .Z(n205) );
  AO2 U232 ( .A(A[35]), .B(B[35]), .C(n40), .D(n206), .Z(n158) );
  EON1 U233 ( .A(n207), .B(n208), .C(B[34]), .D(A[34]), .Z(n206) );
  AO2 U234 ( .A(A[33]), .B(B[33]), .C(B[32]), .D(n209), .Z(n207) );
  NR2 U235 ( .A(n41), .B(n210), .Z(n209) );
  NR4 U236 ( .A(n212), .B(n211), .C(n208), .D(n210), .Z(n154) );
  NR2 U237 ( .A(B[33]), .B(A[33]), .Z(n210) );
  NR2 U238 ( .A(B[34]), .B(A[34]), .Z(n208) );
  NR2 U239 ( .A(B[35]), .B(A[35]), .Z(n211) );
  NR2 U240 ( .A(B[32]), .B(A[32]), .Z(n212) );
  EO1 U241 ( .A(A[31]), .B(B[31]), .C(n213), .D(n214), .Z(n153) );
  AO5 U242 ( .A(A[30]), .B(B[30]), .C(n215), .Z(n214) );
  AO7 U243 ( .A(n216), .B(n42), .C(n217), .Z(n215) );
  AO7 U244 ( .A(A[29]), .B(n43), .C(B[29]), .Z(n217) );
  AO6 U245 ( .A(n218), .B(A[28]), .C(n44), .Z(n216) );
  AO7 U246 ( .A(A[28]), .B(n218), .C(B[28]), .Z(n219) );
  EON1 U247 ( .A(n220), .B(n221), .C(A[27]), .D(B[27]), .Z(n218) );
  AO5 U248 ( .A(A[26]), .B(B[26]), .C(n45), .Z(n221) );
  AO6 U249 ( .A(n223), .B(A[25]), .C(n46), .Z(n222) );
  AO7 U250 ( .A(A[25]), .B(n223), .C(B[25]), .Z(n224) );
  AO7 U251 ( .A(n225), .B(n47), .C(n226), .Z(n223) );
  AO7 U252 ( .A(A[24]), .B(n48), .C(B[24]), .Z(n226) );
  AO2 U253 ( .A(n227), .B(A[23]), .C(B[23]), .D(n228), .Z(n225) );
  OR2 U254 ( .A(n227), .B(A[23]), .Z(n228) );
  AO7 U255 ( .A(n229), .B(n49), .C(n230), .Z(n227) );
  AO7 U256 ( .A(A[22]), .B(n50), .C(B[22]), .Z(n230) );
  NR2 U257 ( .A(A[27]), .B(B[27]), .Z(n220) );
  NR2 U258 ( .A(A[31]), .B(B[31]), .Z(n213) );
  ND2 U259 ( .A(n37), .B(n194), .Z(n204) );
  ND2 U260 ( .A(B[36]), .B(A[36]), .Z(n194) );
  NR2 U261 ( .A(B[36]), .B(A[36]), .Z(n203) );
endmodule


module LOG_POLY_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [21:0] A;
  input [47:0] B;
  output [69:0] PRODUCT;
  input TC;
  wire   \ab[21][47] , \ab[21][46] , \ab[21][45] , \ab[21][44] , \ab[21][43] ,
         \ab[21][42] , \ab[21][41] , \ab[21][40] , \ab[21][39] , \ab[21][38] ,
         \ab[21][37] , \ab[21][36] , \ab[21][35] , \ab[21][34] , \ab[21][33] ,
         \ab[21][32] , \ab[21][31] , \ab[21][30] , \ab[21][29] , \ab[21][28] ,
         \ab[21][27] , \ab[21][26] , \ab[21][25] , \ab[21][24] , \ab[21][23] ,
         \ab[21][22] , \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] ,
         \ab[21][17] , \ab[21][16] , \ab[21][15] , \ab[21][14] , \ab[21][13] ,
         \ab[21][12] , \ab[21][11] , \ab[21][10] , \ab[21][9] , \ab[21][8] ,
         \ab[21][7] , \ab[21][6] , \ab[21][5] , \ab[21][4] , \ab[21][3] ,
         \ab[21][2] , \ab[21][1] , \ab[21][0] , \ab[20][47] , \ab[20][46] ,
         \ab[20][45] , \ab[20][44] , \ab[20][43] , \ab[20][42] , \ab[20][41] ,
         \ab[20][40] , \ab[20][39] , \ab[20][38] , \ab[20][37] , \ab[20][36] ,
         \ab[20][35] , \ab[20][34] , \ab[20][33] , \ab[20][32] , \ab[20][31] ,
         \ab[20][30] , \ab[20][29] , \ab[20][28] , \ab[20][27] , \ab[20][26] ,
         \ab[20][25] , \ab[20][24] , \ab[20][23] , \ab[20][22] , \ab[20][21] ,
         \ab[20][20] , \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] ,
         \ab[20][15] , \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] ,
         \ab[20][10] , \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] ,
         \ab[20][5] , \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] ,
         \ab[20][0] , \ab[19][47] , \ab[19][46] , \ab[19][45] , \ab[19][44] ,
         \ab[19][43] , \ab[19][42] , \ab[19][41] , \ab[19][40] , \ab[19][39] ,
         \ab[19][38] , \ab[19][37] , \ab[19][36] , \ab[19][35] , \ab[19][34] ,
         \ab[19][33] , \ab[19][32] , \ab[19][31] , \ab[19][30] , \ab[19][29] ,
         \ab[19][28] , \ab[19][27] , \ab[19][26] , \ab[19][25] , \ab[19][24] ,
         \ab[19][23] , \ab[19][22] , \ab[19][21] , \ab[19][20] , \ab[19][19] ,
         \ab[19][18] , \ab[19][17] , \ab[19][16] , \ab[19][15] , \ab[19][14] ,
         \ab[19][13] , \ab[19][12] , \ab[19][11] , \ab[19][10] , \ab[19][9] ,
         \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] , \ab[19][4] ,
         \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] , \ab[18][47] ,
         \ab[18][46] , \ab[18][45] , \ab[18][44] , \ab[18][43] , \ab[18][42] ,
         \ab[18][41] , \ab[18][40] , \ab[18][39] , \ab[18][38] , \ab[18][37] ,
         \ab[18][36] , \ab[18][35] , \ab[18][34] , \ab[18][33] , \ab[18][32] ,
         \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] , \ab[18][27] ,
         \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] , \ab[18][22] ,
         \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] , \ab[18][17] ,
         \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] , \ab[18][12] ,
         \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] , \ab[18][7] ,
         \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] , \ab[18][2] ,
         \ab[18][1] , \ab[18][0] , \ab[17][47] , \ab[17][46] , \ab[17][45] ,
         \ab[17][44] , \ab[17][43] , \ab[17][42] , \ab[17][41] , \ab[17][40] ,
         \ab[17][39] , \ab[17][38] , \ab[17][37] , \ab[17][36] , \ab[17][35] ,
         \ab[17][34] , \ab[17][33] , \ab[17][32] , \ab[17][31] , \ab[17][30] ,
         \ab[17][29] , \ab[17][28] , \ab[17][27] , \ab[17][26] , \ab[17][25] ,
         \ab[17][24] , \ab[17][23] , \ab[17][22] , \ab[17][21] , \ab[17][20] ,
         \ab[17][19] , \ab[17][18] , \ab[17][17] , \ab[17][16] , \ab[17][15] ,
         \ab[17][14] , \ab[17][13] , \ab[17][12] , \ab[17][11] , \ab[17][10] ,
         \ab[17][9] , \ab[17][8] , \ab[17][7] , \ab[17][6] , \ab[17][5] ,
         \ab[17][4] , \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] ,
         \ab[16][47] , \ab[16][46] , \ab[16][45] , \ab[16][44] , \ab[16][43] ,
         \ab[16][42] , \ab[16][41] , \ab[16][40] , \ab[16][39] , \ab[16][38] ,
         \ab[16][37] , \ab[16][36] , \ab[16][35] , \ab[16][34] , \ab[16][33] ,
         \ab[16][32] , \ab[16][31] , \ab[16][30] , \ab[16][29] , \ab[16][28] ,
         \ab[16][27] , \ab[16][26] , \ab[16][25] , \ab[16][24] , \ab[16][23] ,
         \ab[16][22] , \ab[16][21] , \ab[16][20] , \ab[16][19] , \ab[16][18] ,
         \ab[16][17] , \ab[16][16] , \ab[16][15] , \ab[16][14] , \ab[16][13] ,
         \ab[16][12] , \ab[16][11] , \ab[16][10] , \ab[16][9] , \ab[16][8] ,
         \ab[16][7] , \ab[16][6] , \ab[16][5] , \ab[16][4] , \ab[16][3] ,
         \ab[16][2] , \ab[16][1] , \ab[16][0] , \ab[15][47] , \ab[15][46] ,
         \ab[15][45] , \ab[15][44] , \ab[15][43] , \ab[15][42] , \ab[15][41] ,
         \ab[15][40] , \ab[15][39] , \ab[15][38] , \ab[15][37] , \ab[15][36] ,
         \ab[15][35] , \ab[15][34] , \ab[15][33] , \ab[15][32] , \ab[15][31] ,
         \ab[15][30] , \ab[15][29] , \ab[15][28] , \ab[15][27] , \ab[15][26] ,
         \ab[15][25] , \ab[15][24] , \ab[15][23] , \ab[15][22] , \ab[15][21] ,
         \ab[15][20] , \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] ,
         \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][47] , \ab[14][46] , \ab[14][45] , \ab[14][44] ,
         \ab[14][43] , \ab[14][42] , \ab[14][41] , \ab[14][40] , \ab[14][39] ,
         \ab[14][38] , \ab[14][37] , \ab[14][36] , \ab[14][35] , \ab[14][34] ,
         \ab[14][33] , \ab[14][32] , \ab[14][31] , \ab[14][30] , \ab[14][29] ,
         \ab[14][28] , \ab[14][27] , \ab[14][26] , \ab[14][25] , \ab[14][24] ,
         \ab[14][23] , \ab[14][22] , \ab[14][21] , \ab[14][20] , \ab[14][19] ,
         \ab[14][18] , \ab[14][17] , \ab[14][16] , \ab[14][15] , \ab[14][14] ,
         \ab[14][13] , \ab[14][12] , \ab[14][11] , \ab[14][10] , \ab[14][9] ,
         \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] ,
         \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][47] ,
         \ab[13][46] , \ab[13][45] , \ab[13][44] , \ab[13][43] , \ab[13][42] ,
         \ab[13][41] , \ab[13][40] , \ab[13][39] , \ab[13][38] , \ab[13][37] ,
         \ab[13][36] , \ab[13][35] , \ab[13][34] , \ab[13][33] , \ab[13][32] ,
         \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] , \ab[13][27] ,
         \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] , \ab[13][22] ,
         \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] , \ab[13][17] ,
         \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] , \ab[13][12] ,
         \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] , \ab[13][7] ,
         \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] , \ab[13][2] ,
         \ab[13][1] , \ab[13][0] , \ab[12][47] , \ab[12][46] , \ab[12][45] ,
         \ab[12][44] , \ab[12][43] , \ab[12][42] , \ab[12][41] , \ab[12][40] ,
         \ab[12][39] , \ab[12][38] , \ab[12][37] , \ab[12][36] , \ab[12][35] ,
         \ab[12][34] , \ab[12][33] , \ab[12][32] , \ab[12][31] , \ab[12][30] ,
         \ab[12][29] , \ab[12][28] , \ab[12][27] , \ab[12][26] , \ab[12][25] ,
         \ab[12][24] , \ab[12][23] , \ab[12][22] , \ab[12][21] , \ab[12][20] ,
         \ab[12][19] , \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][47] , \ab[11][46] , \ab[11][45] , \ab[11][44] , \ab[11][43] ,
         \ab[11][42] , \ab[11][41] , \ab[11][40] , \ab[11][39] , \ab[11][38] ,
         \ab[11][37] , \ab[11][36] , \ab[11][35] , \ab[11][34] , \ab[11][33] ,
         \ab[11][32] , \ab[11][31] , \ab[11][30] , \ab[11][29] , \ab[11][28] ,
         \ab[11][27] , \ab[11][26] , \ab[11][25] , \ab[11][24] , \ab[11][23] ,
         \ab[11][22] , \ab[11][21] , \ab[11][20] , \ab[11][19] , \ab[11][18] ,
         \ab[11][17] , \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] ,
         \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] ,
         \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] ,
         \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][47] , \ab[10][46] ,
         \ab[10][45] , \ab[10][44] , \ab[10][43] , \ab[10][42] , \ab[10][41] ,
         \ab[10][40] , \ab[10][39] , \ab[10][38] , \ab[10][37] , \ab[10][36] ,
         \ab[10][35] , \ab[10][34] , \ab[10][33] , \ab[10][32] , \ab[10][31] ,
         \ab[10][30] , \ab[10][29] , \ab[10][28] , \ab[10][27] , \ab[10][26] ,
         \ab[10][25] , \ab[10][24] , \ab[10][23] , \ab[10][22] , \ab[10][21] ,
         \ab[10][20] , \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][47] , \ab[9][46] , \ab[9][45] , \ab[9][44] ,
         \ab[9][43] , \ab[9][42] , \ab[9][41] , \ab[9][40] , \ab[9][39] ,
         \ab[9][38] , \ab[9][37] , \ab[9][36] , \ab[9][35] , \ab[9][34] ,
         \ab[9][33] , \ab[9][32] , \ab[9][31] , \ab[9][30] , \ab[9][29] ,
         \ab[9][28] , \ab[9][27] , \ab[9][26] , \ab[9][25] , \ab[9][24] ,
         \ab[9][23] , \ab[9][22] , \ab[9][21] , \ab[9][20] , \ab[9][19] ,
         \ab[9][18] , \ab[9][17] , \ab[9][16] , \ab[9][15] , \ab[9][14] ,
         \ab[9][13] , \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] ,
         \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] ,
         \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][47] ,
         \ab[8][46] , \ab[8][45] , \ab[8][44] , \ab[8][43] , \ab[8][42] ,
         \ab[8][41] , \ab[8][40] , \ab[8][39] , \ab[8][38] , \ab[8][37] ,
         \ab[8][36] , \ab[8][35] , \ab[8][34] , \ab[8][33] , \ab[8][32] ,
         \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] , \ab[8][27] ,
         \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] , \ab[8][22] ,
         \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] , \ab[8][17] ,
         \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] , \ab[8][12] ,
         \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] ,
         \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] ,
         \ab[8][1] , \ab[8][0] , \ab[7][47] , \ab[7][46] , \ab[7][45] ,
         \ab[7][44] , \ab[7][43] , \ab[7][42] , \ab[7][41] , \ab[7][40] ,
         \ab[7][39] , \ab[7][38] , \ab[7][37] , \ab[7][36] , \ab[7][35] ,
         \ab[7][34] , \ab[7][33] , \ab[7][32] , \ab[7][31] , \ab[7][30] ,
         \ab[7][29] , \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][47] , \ab[6][46] , \ab[6][45] , \ab[6][44] , \ab[6][43] ,
         \ab[6][42] , \ab[6][41] , \ab[6][40] , \ab[6][39] , \ab[6][38] ,
         \ab[6][37] , \ab[6][36] , \ab[6][35] , \ab[6][34] , \ab[6][33] ,
         \ab[6][32] , \ab[6][31] , \ab[6][30] , \ab[6][29] , \ab[6][28] ,
         \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] , \ab[6][23] ,
         \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] , \ab[6][18] ,
         \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] ,
         \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] ,
         \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] ,
         \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][47] , \ab[5][46] ,
         \ab[5][45] , \ab[5][44] , \ab[5][43] , \ab[5][42] , \ab[5][41] ,
         \ab[5][40] , \ab[5][39] , \ab[5][38] , \ab[5][37] , \ab[5][36] ,
         \ab[5][35] , \ab[5][34] , \ab[5][33] , \ab[5][32] , \ab[5][31] ,
         \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] ,
         \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][47] , \ab[4][46] , \ab[4][45] , \ab[4][44] ,
         \ab[4][43] , \ab[4][42] , \ab[4][41] , \ab[4][40] , \ab[4][39] ,
         \ab[4][38] , \ab[4][37] , \ab[4][36] , \ab[4][35] , \ab[4][34] ,
         \ab[4][33] , \ab[4][32] , \ab[4][31] , \ab[4][30] , \ab[4][29] ,
         \ab[4][28] , \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] ,
         \ab[4][23] , \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] ,
         \ab[4][18] , \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] ,
         \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] ,
         \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] ,
         \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][47] ,
         \ab[3][46] , \ab[3][45] , \ab[3][44] , \ab[3][43] , \ab[3][42] ,
         \ab[3][41] , \ab[3][40] , \ab[3][39] , \ab[3][38] , \ab[3][37] ,
         \ab[3][36] , \ab[3][35] , \ab[3][34] , \ab[3][33] , \ab[3][32] ,
         \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] , \ab[3][27] ,
         \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] , \ab[3][22] ,
         \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] , \ab[3][17] ,
         \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] , \ab[3][12] ,
         \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] ,
         \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] ,
         \ab[3][1] , \ab[3][0] , \ab[2][47] , \ab[2][46] , \ab[2][45] ,
         \ab[2][44] , \ab[2][43] , \ab[2][42] , \ab[2][41] , \ab[2][40] ,
         \ab[2][39] , \ab[2][38] , \ab[2][37] , \ab[2][36] , \ab[2][35] ,
         \ab[2][34] , \ab[2][33] , \ab[2][32] , \ab[2][31] , \ab[2][30] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][47] , \ab[1][46] , \ab[1][45] , \ab[1][44] , \ab[1][43] ,
         \ab[1][42] , \ab[1][41] , \ab[1][40] , \ab[1][39] , \ab[1][38] ,
         \ab[1][37] , \ab[1][36] , \ab[1][35] , \ab[1][34] , \ab[1][33] ,
         \ab[1][32] , \ab[1][31] , \ab[1][30] , \ab[1][29] , \ab[1][28] ,
         \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] , \ab[1][23] ,
         \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] ,
         \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[0][47] , \ab[0][46] , \ab[0][45] ,
         \ab[0][44] , \ab[0][43] , \ab[0][42] , \ab[0][41] , \ab[0][40] ,
         \ab[0][39] , \ab[0][38] , \ab[0][37] , \ab[0][36] , \ab[0][35] ,
         \ab[0][34] , \ab[0][33] , \ab[0][32] , \ab[0][31] , \ab[0][30] ,
         \ab[0][29] , \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] ,
         \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] ,
         \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] ,
         \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \CARRYB[11][15] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][46] , \CARRYB[10][45] , \CARRYB[10][44] ,
         \CARRYB[10][43] , \CARRYB[10][42] , \CARRYB[10][41] ,
         \CARRYB[10][40] , \CARRYB[10][39] , \CARRYB[10][38] ,
         \CARRYB[10][37] , \CARRYB[10][36] , \CARRYB[10][35] ,
         \CARRYB[10][34] , \CARRYB[10][33] , \CARRYB[10][32] ,
         \CARRYB[10][31] , \CARRYB[10][30] , \CARRYB[10][29] ,
         \CARRYB[10][28] , \CARRYB[10][27] , \CARRYB[10][26] ,
         \CARRYB[10][25] , \CARRYB[10][24] , \CARRYB[10][23] ,
         \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][46] ,
         \CARRYB[9][45] , \CARRYB[9][44] , \CARRYB[9][43] , \CARRYB[9][42] ,
         \CARRYB[9][41] , \CARRYB[9][40] , \CARRYB[9][39] , \CARRYB[9][38] ,
         \CARRYB[9][37] , \CARRYB[9][36] , \CARRYB[9][35] , \CARRYB[9][34] ,
         \CARRYB[9][33] , \CARRYB[9][32] , \CARRYB[9][31] , \CARRYB[9][30] ,
         \CARRYB[9][29] , \CARRYB[9][28] , \CARRYB[9][27] , \CARRYB[9][26] ,
         \CARRYB[9][25] , \CARRYB[9][24] , \CARRYB[9][23] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][46] , \CARRYB[8][45] ,
         \CARRYB[8][44] , \CARRYB[8][43] , \CARRYB[8][42] , \CARRYB[8][41] ,
         \CARRYB[8][40] , \CARRYB[8][39] , \CARRYB[8][38] , \CARRYB[8][37] ,
         \CARRYB[8][36] , \CARRYB[8][35] , \CARRYB[8][34] , \CARRYB[8][33] ,
         \CARRYB[8][32] , \CARRYB[8][31] , \CARRYB[8][30] , \CARRYB[8][29] ,
         \CARRYB[8][28] , \CARRYB[8][27] , \CARRYB[8][26] , \CARRYB[8][25] ,
         \CARRYB[8][24] , \CARRYB[8][23] , \CARRYB[8][22] , \CARRYB[8][21] ,
         \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] ,
         \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][46] , \CARRYB[7][45] , \CARRYB[7][44] ,
         \CARRYB[7][43] , \CARRYB[7][42] , \CARRYB[7][41] , \CARRYB[7][40] ,
         \CARRYB[7][39] , \CARRYB[7][38] , \CARRYB[7][37] , \CARRYB[7][36] ,
         \CARRYB[7][35] , \CARRYB[7][34] , \CARRYB[7][33] , \CARRYB[7][32] ,
         \CARRYB[7][31] , \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] ,
         \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] ,
         \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][46] , \CARRYB[6][45] , \CARRYB[6][44] , \CARRYB[6][43] ,
         \CARRYB[6][42] , \CARRYB[6][41] , \CARRYB[6][40] , \CARRYB[6][39] ,
         \CARRYB[6][38] , \CARRYB[6][37] , \CARRYB[6][36] , \CARRYB[6][35] ,
         \CARRYB[6][34] , \CARRYB[6][33] , \CARRYB[6][32] , \CARRYB[6][31] ,
         \CARRYB[6][30] , \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] ,
         \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][46] ,
         \CARRYB[5][45] , \CARRYB[5][44] , \CARRYB[5][43] , \CARRYB[5][42] ,
         \CARRYB[5][41] , \CARRYB[5][40] , \CARRYB[5][39] , \CARRYB[5][38] ,
         \CARRYB[5][37] , \CARRYB[5][36] , \CARRYB[5][35] , \CARRYB[5][34] ,
         \CARRYB[5][33] , \CARRYB[5][32] , \CARRYB[5][31] , \CARRYB[5][30] ,
         \CARRYB[5][29] , \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][46] , \CARRYB[4][45] ,
         \CARRYB[4][44] , \CARRYB[4][43] , \CARRYB[4][42] , \CARRYB[4][41] ,
         \CARRYB[4][40] , \CARRYB[4][39] , \CARRYB[4][38] , \CARRYB[4][37] ,
         \CARRYB[4][36] , \CARRYB[4][35] , \CARRYB[4][34] , \CARRYB[4][33] ,
         \CARRYB[4][32] , \CARRYB[4][31] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][46] , \CARRYB[3][45] , \CARRYB[3][44] ,
         \CARRYB[3][43] , \CARRYB[3][42] , \CARRYB[3][41] , \CARRYB[3][40] ,
         \CARRYB[3][39] , \CARRYB[3][38] , \CARRYB[3][37] , \CARRYB[3][36] ,
         \CARRYB[3][35] , \CARRYB[3][34] , \CARRYB[3][33] , \CARRYB[3][32] ,
         \CARRYB[3][31] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][46] , \CARRYB[2][45] , \CARRYB[2][44] , \CARRYB[2][43] ,
         \CARRYB[2][42] , \CARRYB[2][41] , \CARRYB[2][40] , \CARRYB[2][39] ,
         \CARRYB[2][38] , \CARRYB[2][37] , \CARRYB[2][36] , \CARRYB[2][35] ,
         \CARRYB[2][34] , \CARRYB[2][33] , \CARRYB[2][32] , \CARRYB[2][31] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][46] ,
         \CARRYB[1][45] , \CARRYB[1][44] , \CARRYB[1][43] , \CARRYB[1][42] ,
         \CARRYB[1][41] , \CARRYB[1][40] , \CARRYB[1][39] , \CARRYB[1][38] ,
         \CARRYB[1][37] , \CARRYB[1][36] , \CARRYB[1][35] , \CARRYB[1][34] ,
         \CARRYB[1][33] , \CARRYB[1][32] , \CARRYB[1][31] , \CARRYB[1][30] ,
         \CARRYB[1][29] , \CARRYB[1][28] , \CARRYB[1][27] , \CARRYB[1][26] ,
         \CARRYB[1][25] , \CARRYB[1][24] , \CARRYB[1][23] , \CARRYB[1][22] ,
         \CARRYB[1][21] , \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] ,
         \CARRYB[1][17] , \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] ,
         \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] ,
         \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] ,
         \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] ,
         \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[11][15] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][46] , \SUMB[10][45] , \SUMB[10][44] ,
         \SUMB[10][43] , \SUMB[10][42] , \SUMB[10][41] , \SUMB[10][40] ,
         \SUMB[10][39] , \SUMB[10][38] , \SUMB[10][37] , \SUMB[10][36] ,
         \SUMB[10][35] , \SUMB[10][34] , \SUMB[10][33] , \SUMB[10][32] ,
         \SUMB[10][31] , \SUMB[10][30] , \SUMB[10][29] , \SUMB[10][28] ,
         \SUMB[10][27] , \SUMB[10][26] , \SUMB[10][25] , \SUMB[10][24] ,
         \SUMB[10][23] , \SUMB[10][22] , \SUMB[10][21] , \SUMB[10][20] ,
         \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] , \SUMB[10][16] ,
         \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] , \SUMB[10][12] ,
         \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] , \SUMB[10][8] ,
         \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] ,
         \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][46] ,
         \SUMB[9][45] , \SUMB[9][44] , \SUMB[9][43] , \SUMB[9][42] ,
         \SUMB[9][41] , \SUMB[9][40] , \SUMB[9][39] , \SUMB[9][38] ,
         \SUMB[9][37] , \SUMB[9][36] , \SUMB[9][35] , \SUMB[9][34] ,
         \SUMB[9][33] , \SUMB[9][32] , \SUMB[9][31] , \SUMB[9][30] ,
         \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] , \SUMB[9][26] ,
         \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] , \SUMB[9][22] ,
         \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] ,
         \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][46] ,
         \SUMB[8][45] , \SUMB[8][44] , \SUMB[8][43] , \SUMB[8][42] ,
         \SUMB[8][41] , \SUMB[8][40] , \SUMB[8][39] , \SUMB[8][38] ,
         \SUMB[8][37] , \SUMB[8][36] , \SUMB[8][35] , \SUMB[8][34] ,
         \SUMB[8][33] , \SUMB[8][32] , \SUMB[8][31] , \SUMB[8][30] ,
         \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] , \SUMB[8][26] ,
         \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] , \SUMB[8][22] ,
         \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] ,
         \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][46] ,
         \SUMB[7][45] , \SUMB[7][44] , \SUMB[7][43] , \SUMB[7][42] ,
         \SUMB[7][41] , \SUMB[7][40] , \SUMB[7][39] , \SUMB[7][38] ,
         \SUMB[7][37] , \SUMB[7][36] , \SUMB[7][35] , \SUMB[7][34] ,
         \SUMB[7][33] , \SUMB[7][32] , \SUMB[7][31] , \SUMB[7][30] ,
         \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] ,
         \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][46] ,
         \SUMB[6][45] , \SUMB[6][44] , \SUMB[6][43] , \SUMB[6][42] ,
         \SUMB[6][41] , \SUMB[6][40] , \SUMB[6][39] , \SUMB[6][38] ,
         \SUMB[6][37] , \SUMB[6][36] , \SUMB[6][35] , \SUMB[6][34] ,
         \SUMB[6][33] , \SUMB[6][32] , \SUMB[6][31] , \SUMB[6][30] ,
         \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][46] ,
         \SUMB[5][45] , \SUMB[5][44] , \SUMB[5][43] , \SUMB[5][42] ,
         \SUMB[5][41] , \SUMB[5][40] , \SUMB[5][39] , \SUMB[5][38] ,
         \SUMB[5][37] , \SUMB[5][36] , \SUMB[5][35] , \SUMB[5][34] ,
         \SUMB[5][33] , \SUMB[5][32] , \SUMB[5][31] , \SUMB[5][30] ,
         \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] ,
         \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][46] ,
         \SUMB[4][45] , \SUMB[4][44] , \SUMB[4][43] , \SUMB[4][42] ,
         \SUMB[4][41] , \SUMB[4][40] , \SUMB[4][39] , \SUMB[4][38] ,
         \SUMB[4][37] , \SUMB[4][36] , \SUMB[4][35] , \SUMB[4][34] ,
         \SUMB[4][33] , \SUMB[4][32] , \SUMB[4][31] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][46] ,
         \SUMB[3][45] , \SUMB[3][44] , \SUMB[3][43] , \SUMB[3][42] ,
         \SUMB[3][41] , \SUMB[3][40] , \SUMB[3][39] , \SUMB[3][38] ,
         \SUMB[3][37] , \SUMB[3][36] , \SUMB[3][35] , \SUMB[3][34] ,
         \SUMB[3][33] , \SUMB[3][32] , \SUMB[3][31] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][46] ,
         \SUMB[2][45] , \SUMB[2][44] , \SUMB[2][43] , \SUMB[2][42] ,
         \SUMB[2][41] , \SUMB[2][40] , \SUMB[2][39] , \SUMB[2][38] ,
         \SUMB[2][37] , \SUMB[2][36] , \SUMB[2][35] , \SUMB[2][34] ,
         \SUMB[2][33] , \SUMB[2][32] , \SUMB[2][31] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][46] ,
         \SUMB[1][45] , \SUMB[1][44] , \SUMB[1][43] , \SUMB[1][42] ,
         \SUMB[1][41] , \SUMB[1][40] , \SUMB[1][39] , \SUMB[1][38] ,
         \SUMB[1][37] , \SUMB[1][36] , \SUMB[1][35] , \SUMB[1][34] ,
         \SUMB[1][33] , \SUMB[1][32] , \SUMB[1][31] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[21][46] , \CARRYB[21][45] , \CARRYB[21][44] ,
         \CARRYB[21][43] , \CARRYB[21][42] , \CARRYB[21][41] ,
         \CARRYB[21][40] , \CARRYB[21][39] , \CARRYB[21][38] ,
         \CARRYB[21][37] , \CARRYB[21][36] , \CARRYB[21][35] ,
         \CARRYB[21][34] , \CARRYB[21][33] , \CARRYB[21][32] ,
         \CARRYB[21][31] , \CARRYB[21][30] , \CARRYB[21][29] ,
         \CARRYB[21][28] , \CARRYB[21][27] , \CARRYB[21][26] ,
         \CARRYB[21][25] , \CARRYB[21][24] , \CARRYB[21][23] ,
         \CARRYB[21][22] , \CARRYB[21][21] , \CARRYB[21][20] ,
         \CARRYB[21][19] , \CARRYB[21][18] , \CARRYB[21][17] ,
         \CARRYB[21][16] , \CARRYB[21][15] , \CARRYB[21][14] ,
         \CARRYB[21][13] , \CARRYB[21][12] , \CARRYB[21][11] ,
         \CARRYB[21][10] , \CARRYB[21][9] , \CARRYB[21][8] , \CARRYB[21][7] ,
         \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] , \CARRYB[21][3] ,
         \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] , \CARRYB[20][46] ,
         \CARRYB[20][45] , \CARRYB[20][44] , \CARRYB[20][43] ,
         \CARRYB[20][42] , \CARRYB[20][41] , \CARRYB[20][40] ,
         \CARRYB[20][39] , \CARRYB[20][38] , \CARRYB[20][37] ,
         \CARRYB[20][36] , \CARRYB[20][35] , \CARRYB[20][34] ,
         \CARRYB[20][33] , \CARRYB[20][32] , \CARRYB[20][31] ,
         \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][46] , \CARRYB[19][45] , \CARRYB[19][44] ,
         \CARRYB[19][43] , \CARRYB[19][42] , \CARRYB[19][41] ,
         \CARRYB[19][40] , \CARRYB[19][39] , \CARRYB[19][38] ,
         \CARRYB[19][37] , \CARRYB[19][36] , \CARRYB[19][35] ,
         \CARRYB[19][34] , \CARRYB[19][33] , \CARRYB[19][32] ,
         \CARRYB[19][31] , \CARRYB[19][30] , \CARRYB[19][29] ,
         \CARRYB[19][28] , \CARRYB[19][27] , \CARRYB[19][26] ,
         \CARRYB[19][25] , \CARRYB[19][24] , \CARRYB[19][23] ,
         \CARRYB[19][22] , \CARRYB[19][21] , \CARRYB[19][20] ,
         \CARRYB[19][19] , \CARRYB[19][18] , \CARRYB[19][17] ,
         \CARRYB[19][16] , \CARRYB[19][15] , \CARRYB[19][14] ,
         \CARRYB[19][13] , \CARRYB[19][12] , \CARRYB[19][11] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][46] ,
         \CARRYB[18][45] , \CARRYB[18][44] , \CARRYB[18][43] ,
         \CARRYB[18][42] , \CARRYB[18][41] , \CARRYB[18][40] ,
         \CARRYB[18][39] , \CARRYB[18][38] , \CARRYB[18][37] ,
         \CARRYB[18][36] , \CARRYB[18][35] , \CARRYB[18][34] ,
         \CARRYB[18][33] , \CARRYB[18][32] , \CARRYB[18][31] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][46] , \CARRYB[17][45] , \CARRYB[17][44] ,
         \CARRYB[17][43] , \CARRYB[17][42] , \CARRYB[17][41] ,
         \CARRYB[17][40] , \CARRYB[17][39] , \CARRYB[17][38] ,
         \CARRYB[17][37] , \CARRYB[17][36] , \CARRYB[17][35] ,
         \CARRYB[17][34] , \CARRYB[17][33] , \CARRYB[17][32] ,
         \CARRYB[17][31] , \CARRYB[17][30] , \CARRYB[17][29] ,
         \CARRYB[17][28] , \CARRYB[17][27] , \CARRYB[17][26] ,
         \CARRYB[17][25] , \CARRYB[17][24] , \CARRYB[17][23] ,
         \CARRYB[17][22] , \CARRYB[17][21] , \CARRYB[17][20] ,
         \CARRYB[17][19] , \CARRYB[17][18] , \CARRYB[17][17] ,
         \CARRYB[17][16] , \CARRYB[17][15] , \CARRYB[17][14] ,
         \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][46] ,
         \CARRYB[16][45] , \CARRYB[16][44] , \CARRYB[16][43] ,
         \CARRYB[16][42] , \CARRYB[16][41] , \CARRYB[16][40] ,
         \CARRYB[16][39] , \CARRYB[16][38] , \CARRYB[16][37] ,
         \CARRYB[16][36] , \CARRYB[16][35] , \CARRYB[16][34] ,
         \CARRYB[16][33] , \CARRYB[16][32] , \CARRYB[16][31] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \CARRYB[15][46] , \CARRYB[15][45] , \CARRYB[15][44] ,
         \CARRYB[15][43] , \CARRYB[15][42] , \CARRYB[15][41] ,
         \CARRYB[15][40] , \CARRYB[15][39] , \CARRYB[15][38] ,
         \CARRYB[15][37] , \CARRYB[15][36] , \CARRYB[15][35] ,
         \CARRYB[15][34] , \CARRYB[15][33] , \CARRYB[15][32] ,
         \CARRYB[15][31] , \CARRYB[15][30] , \CARRYB[15][29] ,
         \CARRYB[15][28] , \CARRYB[15][27] , \CARRYB[15][26] ,
         \CARRYB[15][25] , \CARRYB[15][24] , \CARRYB[15][23] ,
         \CARRYB[15][22] , \CARRYB[15][21] , \CARRYB[15][20] ,
         \CARRYB[15][19] , \CARRYB[15][18] , \CARRYB[15][17] ,
         \CARRYB[15][16] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][46] ,
         \CARRYB[14][45] , \CARRYB[14][44] , \CARRYB[14][43] ,
         \CARRYB[14][42] , \CARRYB[14][41] , \CARRYB[14][40] ,
         \CARRYB[14][39] , \CARRYB[14][38] , \CARRYB[14][37] ,
         \CARRYB[14][36] , \CARRYB[14][35] , \CARRYB[14][34] ,
         \CARRYB[14][33] , \CARRYB[14][32] , \CARRYB[14][31] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][46] , \CARRYB[13][45] , \CARRYB[13][44] ,
         \CARRYB[13][43] , \CARRYB[13][42] , \CARRYB[13][41] ,
         \CARRYB[13][40] , \CARRYB[13][39] , \CARRYB[13][38] ,
         \CARRYB[13][37] , \CARRYB[13][36] , \CARRYB[13][35] ,
         \CARRYB[13][34] , \CARRYB[13][33] , \CARRYB[13][32] ,
         \CARRYB[13][31] , \CARRYB[13][30] , \CARRYB[13][29] ,
         \CARRYB[13][28] , \CARRYB[13][27] , \CARRYB[13][26] ,
         \CARRYB[13][25] , \CARRYB[13][24] , \CARRYB[13][23] ,
         \CARRYB[13][22] , \CARRYB[13][21] , \CARRYB[13][20] ,
         \CARRYB[13][19] , \CARRYB[13][18] , \CARRYB[13][17] ,
         \CARRYB[13][16] , \CARRYB[13][15] , \CARRYB[13][14] ,
         \CARRYB[13][13] , \CARRYB[13][12] , \CARRYB[13][11] ,
         \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] , \CARRYB[13][7] ,
         \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] , \CARRYB[13][3] ,
         \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] , \CARRYB[12][46] ,
         \CARRYB[12][45] , \CARRYB[12][44] , \CARRYB[12][43] ,
         \CARRYB[12][42] , \CARRYB[12][41] , \CARRYB[12][40] ,
         \CARRYB[12][39] , \CARRYB[12][38] , \CARRYB[12][37] ,
         \CARRYB[12][36] , \CARRYB[12][35] , \CARRYB[12][34] ,
         \CARRYB[12][33] , \CARRYB[12][32] , \CARRYB[12][31] ,
         \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][46] , \CARRYB[11][45] , \CARRYB[11][44] ,
         \CARRYB[11][43] , \CARRYB[11][42] , \CARRYB[11][41] ,
         \CARRYB[11][40] , \CARRYB[11][39] , \CARRYB[11][38] ,
         \CARRYB[11][37] , \CARRYB[11][36] , \CARRYB[11][35] ,
         \CARRYB[11][34] , \CARRYB[11][33] , \CARRYB[11][32] ,
         \CARRYB[11][31] , \CARRYB[11][30] , \CARRYB[11][29] ,
         \CARRYB[11][28] , \CARRYB[11][27] , \CARRYB[11][26] ,
         \CARRYB[11][25] , \CARRYB[11][24] , \CARRYB[11][23] ,
         \CARRYB[11][22] , \CARRYB[11][21] , \CARRYB[11][20] ,
         \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \SUMB[21][46] , \SUMB[21][45] , \SUMB[21][44] ,
         \SUMB[21][43] , \SUMB[21][42] , \SUMB[21][41] , \SUMB[21][40] ,
         \SUMB[21][39] , \SUMB[21][38] , \SUMB[21][37] , \SUMB[21][36] ,
         \SUMB[21][35] , \SUMB[21][34] , \SUMB[21][33] , \SUMB[21][32] ,
         \SUMB[21][31] , \SUMB[21][30] , \SUMB[21][29] , \SUMB[21][28] ,
         \SUMB[21][27] , \SUMB[21][26] , \SUMB[21][25] , \SUMB[21][24] ,
         \SUMB[21][23] , \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] ,
         \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] ,
         \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] ,
         \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] ,
         \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] ,
         \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] , \SUMB[21][0] ,
         \SUMB[20][46] , \SUMB[20][45] , \SUMB[20][44] , \SUMB[20][43] ,
         \SUMB[20][42] , \SUMB[20][41] , \SUMB[20][40] , \SUMB[20][39] ,
         \SUMB[20][38] , \SUMB[20][37] , \SUMB[20][36] , \SUMB[20][35] ,
         \SUMB[20][34] , \SUMB[20][33] , \SUMB[20][32] , \SUMB[20][31] ,
         \SUMB[20][30] , \SUMB[20][29] , \SUMB[20][28] , \SUMB[20][27] ,
         \SUMB[20][26] , \SUMB[20][25] , \SUMB[20][24] , \SUMB[20][23] ,
         \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] , \SUMB[20][19] ,
         \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] , \SUMB[20][15] ,
         \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] ,
         \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] ,
         \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] ,
         \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][46] , \SUMB[19][45] ,
         \SUMB[19][44] , \SUMB[19][43] , \SUMB[19][42] , \SUMB[19][41] ,
         \SUMB[19][40] , \SUMB[19][39] , \SUMB[19][38] , \SUMB[19][37] ,
         \SUMB[19][36] , \SUMB[19][35] , \SUMB[19][34] , \SUMB[19][33] ,
         \SUMB[19][32] , \SUMB[19][31] , \SUMB[19][30] , \SUMB[19][29] ,
         \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] , \SUMB[19][25] ,
         \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] , \SUMB[19][21] ,
         \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] ,
         \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] ,
         \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] ,
         \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] ,
         \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] ,
         \SUMB[18][46] , \SUMB[18][45] , \SUMB[18][44] , \SUMB[18][43] ,
         \SUMB[18][42] , \SUMB[18][41] , \SUMB[18][40] , \SUMB[18][39] ,
         \SUMB[18][38] , \SUMB[18][37] , \SUMB[18][36] , \SUMB[18][35] ,
         \SUMB[18][34] , \SUMB[18][33] , \SUMB[18][32] , \SUMB[18][31] ,
         \SUMB[18][30] , \SUMB[18][29] , \SUMB[18][28] , \SUMB[18][27] ,
         \SUMB[18][26] , \SUMB[18][25] , \SUMB[18][24] , \SUMB[18][23] ,
         \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] ,
         \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] ,
         \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] ,
         \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] ,
         \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][46] , \SUMB[17][45] ,
         \SUMB[17][44] , \SUMB[17][43] , \SUMB[17][42] , \SUMB[17][41] ,
         \SUMB[17][40] , \SUMB[17][39] , \SUMB[17][38] , \SUMB[17][37] ,
         \SUMB[17][36] , \SUMB[17][35] , \SUMB[17][34] , \SUMB[17][33] ,
         \SUMB[17][32] , \SUMB[17][31] , \SUMB[17][30] , \SUMB[17][29] ,
         \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] , \SUMB[17][25] ,
         \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] , \SUMB[17][21] ,
         \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] ,
         \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][46] , \SUMB[16][45] , \SUMB[16][44] , \SUMB[16][43] ,
         \SUMB[16][42] , \SUMB[16][41] , \SUMB[16][40] , \SUMB[16][39] ,
         \SUMB[16][38] , \SUMB[16][37] , \SUMB[16][36] , \SUMB[16][35] ,
         \SUMB[16][34] , \SUMB[16][33] , \SUMB[16][32] , \SUMB[16][31] ,
         \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] , \SUMB[16][27] ,
         \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] , \SUMB[16][23] ,
         \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][19] ,
         \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] , \SUMB[16][15] ,
         \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] ,
         \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] ,
         \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] ,
         \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][46] , \SUMB[15][45] ,
         \SUMB[15][44] , \SUMB[15][43] , \SUMB[15][42] , \SUMB[15][41] ,
         \SUMB[15][40] , \SUMB[15][39] , \SUMB[15][38] , \SUMB[15][37] ,
         \SUMB[15][36] , \SUMB[15][35] , \SUMB[15][34] , \SUMB[15][33] ,
         \SUMB[15][32] , \SUMB[15][31] , \SUMB[15][30] , \SUMB[15][29] ,
         \SUMB[15][28] , \SUMB[15][27] , \SUMB[15][26] , \SUMB[15][25] ,
         \SUMB[15][24] , \SUMB[15][23] , \SUMB[15][22] , \SUMB[15][21] ,
         \SUMB[15][20] , \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] ,
         \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][46] , \SUMB[14][45] , \SUMB[14][44] , \SUMB[14][43] ,
         \SUMB[14][42] , \SUMB[14][41] , \SUMB[14][40] , \SUMB[14][39] ,
         \SUMB[14][38] , \SUMB[14][37] , \SUMB[14][36] , \SUMB[14][35] ,
         \SUMB[14][34] , \SUMB[14][33] , \SUMB[14][32] , \SUMB[14][31] ,
         \SUMB[14][30] , \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] ,
         \SUMB[14][26] , \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] ,
         \SUMB[14][22] , \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] ,
         \SUMB[14][18] , \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] ,
         \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] ,
         \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] ,
         \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] ,
         \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][46] , \SUMB[13][45] ,
         \SUMB[13][44] , \SUMB[13][43] , \SUMB[13][42] , \SUMB[13][41] ,
         \SUMB[13][40] , \SUMB[13][39] , \SUMB[13][38] , \SUMB[13][37] ,
         \SUMB[13][36] , \SUMB[13][35] , \SUMB[13][34] , \SUMB[13][33] ,
         \SUMB[13][32] , \SUMB[13][31] , \SUMB[13][30] , \SUMB[13][29] ,
         \SUMB[13][28] , \SUMB[13][27] , \SUMB[13][26] , \SUMB[13][25] ,
         \SUMB[13][24] , \SUMB[13][23] , \SUMB[13][22] , \SUMB[13][21] ,
         \SUMB[13][20] , \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] ,
         \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][46] , \SUMB[12][45] , \SUMB[12][44] , \SUMB[12][43] ,
         \SUMB[12][42] , \SUMB[12][41] , \SUMB[12][40] , \SUMB[12][39] ,
         \SUMB[12][38] , \SUMB[12][37] , \SUMB[12][36] , \SUMB[12][35] ,
         \SUMB[12][34] , \SUMB[12][33] , \SUMB[12][32] , \SUMB[12][31] ,
         \SUMB[12][30] , \SUMB[12][29] , \SUMB[12][28] , \SUMB[12][27] ,
         \SUMB[12][26] , \SUMB[12][25] , \SUMB[12][24] , \SUMB[12][23] ,
         \SUMB[12][22] , \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] ,
         \SUMB[12][18] , \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] ,
         \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] ,
         \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] ,
         \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] ,
         \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][46] , \SUMB[11][45] ,
         \SUMB[11][44] , \SUMB[11][43] , \SUMB[11][42] , \SUMB[11][41] ,
         \SUMB[11][40] , \SUMB[11][39] , \SUMB[11][38] , \SUMB[11][37] ,
         \SUMB[11][36] , \SUMB[11][35] , \SUMB[11][34] , \SUMB[11][33] ,
         \SUMB[11][32] , \SUMB[11][31] , \SUMB[11][30] , \SUMB[11][29] ,
         \SUMB[11][28] , \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] ,
         \SUMB[11][24] , \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] ,
         \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] ,
         \SUMB[11][16] , \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] ,
         \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] ,
         \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] ,
         \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] ,
         \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] ,
         \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] ,
         \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] ,
         \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[67] , \A2[66] ,
         \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] ,
         \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] ,
         \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] ,
         \A2[23] , \A2[22] , \A2[21] , n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37;

  LOG_POLY_DW01_add_4 FS_1 ( .A({1'b0, \A1[66] , \A1[65] , \A1[64] , \A1[63] , 
        \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , 
        \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , 
        \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , 
        \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , 
        \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , 
        \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , 
        \A1[20] , \SUMB[21][0] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , 
        \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[67] , \A2[66] , \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , 
        \A2[60] , \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , 
        \A2[53] , \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , 
        \A2[46] , \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , 
        \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , 
        \A2[32] , \A2[31] , \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , 
        \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, PRODUCT[67:38], 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37}) );
  FA1A S3_20_46 ( .A(\ab[20][46] ), .B(\CARRYB[19][46] ), .CI(\ab[19][47] ), 
        .CO(\CARRYB[20][46] ), .S(\SUMB[20][46] ) );
  FA1A S3_19_46 ( .A(\ab[19][46] ), .B(\CARRYB[18][46] ), .CI(\ab[18][47] ), 
        .CO(\CARRYB[19][46] ), .S(\SUMB[19][46] ) );
  FA1A S3_18_46 ( .A(\ab[18][46] ), .B(\CARRYB[17][46] ), .CI(\ab[17][47] ), 
        .CO(\CARRYB[18][46] ), .S(\SUMB[18][46] ) );
  FA1A S3_17_46 ( .A(\ab[17][46] ), .B(\CARRYB[16][46] ), .CI(\ab[16][47] ), 
        .CO(\CARRYB[17][46] ), .S(\SUMB[17][46] ) );
  FA1A S3_16_46 ( .A(\ab[16][46] ), .B(\CARRYB[15][46] ), .CI(\ab[15][47] ), 
        .CO(\CARRYB[16][46] ), .S(\SUMB[16][46] ) );
  FA1A S3_15_46 ( .A(\ab[15][46] ), .B(\CARRYB[14][46] ), .CI(\ab[14][47] ), 
        .CO(\CARRYB[15][46] ), .S(\SUMB[15][46] ) );
  FA1A S3_14_46 ( .A(\ab[14][46] ), .B(\CARRYB[13][46] ), .CI(\ab[13][47] ), 
        .CO(\CARRYB[14][46] ), .S(\SUMB[14][46] ) );
  FA1A S3_13_46 ( .A(\ab[13][46] ), .B(\CARRYB[12][46] ), .CI(\ab[12][47] ), 
        .CO(\CARRYB[13][46] ), .S(\SUMB[13][46] ) );
  FA1A S3_12_46 ( .A(\ab[12][46] ), .B(\CARRYB[11][46] ), .CI(\ab[11][47] ), 
        .CO(\CARRYB[12][46] ), .S(\SUMB[12][46] ) );
  FA1A S3_11_46 ( .A(\ab[11][46] ), .B(\CARRYB[10][46] ), .CI(\ab[10][47] ), 
        .CO(\CARRYB[11][46] ), .S(\SUMB[11][46] ) );
  FA1A S3_10_46 ( .A(\ab[10][46] ), .B(\CARRYB[9][46] ), .CI(\ab[9][47] ), 
        .CO(\CARRYB[10][46] ), .S(\SUMB[10][46] ) );
  FA1A S3_9_46 ( .A(\ab[9][46] ), .B(\CARRYB[8][46] ), .CI(\ab[8][47] ), .CO(
        \CARRYB[9][46] ), .S(\SUMB[9][46] ) );
  FA1A S3_8_46 ( .A(\ab[8][46] ), .B(\CARRYB[7][46] ), .CI(\ab[7][47] ), .CO(
        \CARRYB[8][46] ), .S(\SUMB[8][46] ) );
  FA1A S3_7_46 ( .A(\ab[7][46] ), .B(\CARRYB[6][46] ), .CI(\ab[6][47] ), .CO(
        \CARRYB[7][46] ), .S(\SUMB[7][46] ) );
  FA1A S3_6_46 ( .A(\ab[6][46] ), .B(\CARRYB[5][46] ), .CI(\ab[5][47] ), .CO(
        \CARRYB[6][46] ), .S(\SUMB[6][46] ) );
  FA1A S3_5_46 ( .A(\ab[5][46] ), .B(\CARRYB[4][46] ), .CI(\ab[4][47] ), .CO(
        \CARRYB[5][46] ), .S(\SUMB[5][46] ) );
  FA1A S3_4_46 ( .A(\ab[4][46] ), .B(\CARRYB[3][46] ), .CI(\ab[3][47] ), .CO(
        \CARRYB[4][46] ), .S(\SUMB[4][46] ) );
  FA1A S3_3_46 ( .A(\ab[3][46] ), .B(\CARRYB[2][46] ), .CI(\ab[2][47] ), .CO(
        \CARRYB[3][46] ), .S(\SUMB[3][46] ) );
  FA1A S5_46 ( .A(\ab[21][46] ), .B(\CARRYB[20][46] ), .CI(\ab[20][47] ), .CO(
        \CARRYB[21][46] ), .S(\SUMB[21][46] ) );
  FA1A S2_20_45 ( .A(\ab[20][45] ), .B(\CARRYB[19][45] ), .CI(\SUMB[19][46] ), 
        .CO(\CARRYB[20][45] ), .S(\SUMB[20][45] ) );
  FA1A S2_19_45 ( .A(\ab[19][45] ), .B(\CARRYB[18][45] ), .CI(\SUMB[18][46] ), 
        .CO(\CARRYB[19][45] ), .S(\SUMB[19][45] ) );
  FA1A S2_18_45 ( .A(\ab[18][45] ), .B(\CARRYB[17][45] ), .CI(\SUMB[17][46] ), 
        .CO(\CARRYB[18][45] ), .S(\SUMB[18][45] ) );
  FA1A S2_17_45 ( .A(\ab[17][45] ), .B(\CARRYB[16][45] ), .CI(\SUMB[16][46] ), 
        .CO(\CARRYB[17][45] ), .S(\SUMB[17][45] ) );
  FA1A S2_16_45 ( .A(\ab[16][45] ), .B(\CARRYB[15][45] ), .CI(\SUMB[15][46] ), 
        .CO(\CARRYB[16][45] ), .S(\SUMB[16][45] ) );
  FA1A S2_15_45 ( .A(\ab[15][45] ), .B(\CARRYB[14][45] ), .CI(\SUMB[14][46] ), 
        .CO(\CARRYB[15][45] ), .S(\SUMB[15][45] ) );
  FA1A S2_14_45 ( .A(\ab[14][45] ), .B(\CARRYB[13][45] ), .CI(\SUMB[13][46] ), 
        .CO(\CARRYB[14][45] ), .S(\SUMB[14][45] ) );
  FA1A S2_13_45 ( .A(\ab[13][45] ), .B(\CARRYB[12][45] ), .CI(\SUMB[12][46] ), 
        .CO(\CARRYB[13][45] ), .S(\SUMB[13][45] ) );
  FA1A S2_12_45 ( .A(\ab[12][45] ), .B(\CARRYB[11][45] ), .CI(\SUMB[11][46] ), 
        .CO(\CARRYB[12][45] ), .S(\SUMB[12][45] ) );
  FA1A S2_11_45 ( .A(\ab[11][45] ), .B(\CARRYB[10][45] ), .CI(\SUMB[10][46] ), 
        .CO(\CARRYB[11][45] ), .S(\SUMB[11][45] ) );
  FA1A S2_10_45 ( .A(\ab[10][45] ), .B(\CARRYB[9][45] ), .CI(\SUMB[9][46] ), 
        .CO(\CARRYB[10][45] ), .S(\SUMB[10][45] ) );
  FA1A S2_9_45 ( .A(\ab[9][45] ), .B(\CARRYB[8][45] ), .CI(\SUMB[8][46] ), 
        .CO(\CARRYB[9][45] ), .S(\SUMB[9][45] ) );
  FA1A S2_8_45 ( .A(\ab[8][45] ), .B(\CARRYB[7][45] ), .CI(\SUMB[7][46] ), 
        .CO(\CARRYB[8][45] ), .S(\SUMB[8][45] ) );
  FA1A S2_7_45 ( .A(\ab[7][45] ), .B(\CARRYB[6][45] ), .CI(\SUMB[6][46] ), 
        .CO(\CARRYB[7][45] ), .S(\SUMB[7][45] ) );
  FA1A S2_6_45 ( .A(\ab[6][45] ), .B(\CARRYB[5][45] ), .CI(\SUMB[5][46] ), 
        .CO(\CARRYB[6][45] ), .S(\SUMB[6][45] ) );
  FA1A S2_5_45 ( .A(\ab[5][45] ), .B(\CARRYB[4][45] ), .CI(\SUMB[4][46] ), 
        .CO(\CARRYB[5][45] ), .S(\SUMB[5][45] ) );
  FA1A S2_4_45 ( .A(\ab[4][45] ), .B(\CARRYB[3][45] ), .CI(\SUMB[3][46] ), 
        .CO(\CARRYB[4][45] ), .S(\SUMB[4][45] ) );
  FA1A S2_3_45 ( .A(\ab[3][45] ), .B(\CARRYB[2][45] ), .CI(\SUMB[2][46] ), 
        .CO(\CARRYB[3][45] ), .S(\SUMB[3][45] ) );
  FA1A S3_2_46 ( .A(\ab[2][46] ), .B(\CARRYB[1][46] ), .CI(\ab[1][47] ), .CO(
        \CARRYB[2][46] ), .S(\SUMB[2][46] ) );
  FA1A S2_2_45 ( .A(\ab[2][45] ), .B(\CARRYB[1][45] ), .CI(\SUMB[1][46] ), 
        .CO(\CARRYB[2][45] ), .S(\SUMB[2][45] ) );
  FA1A S4_45 ( .A(\ab[21][45] ), .B(\CARRYB[20][45] ), .CI(\SUMB[20][46] ), 
        .CO(\CARRYB[21][45] ), .S(\SUMB[21][45] ) );
  FA1A S2_20_44 ( .A(\ab[20][44] ), .B(\CARRYB[19][44] ), .CI(\SUMB[19][45] ), 
        .CO(\CARRYB[20][44] ), .S(\SUMB[20][44] ) );
  FA1A S2_19_44 ( .A(\ab[19][44] ), .B(\CARRYB[18][44] ), .CI(\SUMB[18][45] ), 
        .CO(\CARRYB[19][44] ), .S(\SUMB[19][44] ) );
  FA1A S2_18_44 ( .A(\ab[18][44] ), .B(\CARRYB[17][44] ), .CI(\SUMB[17][45] ), 
        .CO(\CARRYB[18][44] ), .S(\SUMB[18][44] ) );
  FA1A S2_17_44 ( .A(\ab[17][44] ), .B(\CARRYB[16][44] ), .CI(\SUMB[16][45] ), 
        .CO(\CARRYB[17][44] ), .S(\SUMB[17][44] ) );
  FA1A S2_16_44 ( .A(\ab[16][44] ), .B(\CARRYB[15][44] ), .CI(\SUMB[15][45] ), 
        .CO(\CARRYB[16][44] ), .S(\SUMB[16][44] ) );
  FA1A S2_15_44 ( .A(\ab[15][44] ), .B(\CARRYB[14][44] ), .CI(\SUMB[14][45] ), 
        .CO(\CARRYB[15][44] ), .S(\SUMB[15][44] ) );
  FA1A S2_14_44 ( .A(\ab[14][44] ), .B(\CARRYB[13][44] ), .CI(\SUMB[13][45] ), 
        .CO(\CARRYB[14][44] ), .S(\SUMB[14][44] ) );
  FA1A S2_13_44 ( .A(\ab[13][44] ), .B(\CARRYB[12][44] ), .CI(\SUMB[12][45] ), 
        .CO(\CARRYB[13][44] ), .S(\SUMB[13][44] ) );
  FA1A S2_12_44 ( .A(\ab[12][44] ), .B(\CARRYB[11][44] ), .CI(\SUMB[11][45] ), 
        .CO(\CARRYB[12][44] ), .S(\SUMB[12][44] ) );
  FA1A S2_11_44 ( .A(\ab[11][44] ), .B(\CARRYB[10][44] ), .CI(\SUMB[10][45] ), 
        .CO(\CARRYB[11][44] ), .S(\SUMB[11][44] ) );
  FA1A S2_10_44 ( .A(\ab[10][44] ), .B(\CARRYB[9][44] ), .CI(\SUMB[9][45] ), 
        .CO(\CARRYB[10][44] ), .S(\SUMB[10][44] ) );
  FA1A S2_9_44 ( .A(\ab[9][44] ), .B(\CARRYB[8][44] ), .CI(\SUMB[8][45] ), 
        .CO(\CARRYB[9][44] ), .S(\SUMB[9][44] ) );
  FA1A S2_8_44 ( .A(\ab[8][44] ), .B(\CARRYB[7][44] ), .CI(\SUMB[7][45] ), 
        .CO(\CARRYB[8][44] ), .S(\SUMB[8][44] ) );
  FA1A S2_7_44 ( .A(\ab[7][44] ), .B(\CARRYB[6][44] ), .CI(\SUMB[6][45] ), 
        .CO(\CARRYB[7][44] ), .S(\SUMB[7][44] ) );
  FA1A S2_6_44 ( .A(\ab[6][44] ), .B(\CARRYB[5][44] ), .CI(\SUMB[5][45] ), 
        .CO(\CARRYB[6][44] ), .S(\SUMB[6][44] ) );
  FA1A S2_5_44 ( .A(\ab[5][44] ), .B(\CARRYB[4][44] ), .CI(\SUMB[4][45] ), 
        .CO(\CARRYB[5][44] ), .S(\SUMB[5][44] ) );
  FA1A S2_4_44 ( .A(\ab[4][44] ), .B(\CARRYB[3][44] ), .CI(\SUMB[3][45] ), 
        .CO(\CARRYB[4][44] ), .S(\SUMB[4][44] ) );
  FA1A S2_3_44 ( .A(\ab[3][44] ), .B(\CARRYB[2][44] ), .CI(\SUMB[2][45] ), 
        .CO(\CARRYB[3][44] ), .S(\SUMB[3][44] ) );
  FA1A S2_2_44 ( .A(\ab[2][44] ), .B(\CARRYB[1][44] ), .CI(\SUMB[1][45] ), 
        .CO(\CARRYB[2][44] ), .S(\SUMB[2][44] ) );
  FA1A S4_44 ( .A(\ab[21][44] ), .B(\CARRYB[20][44] ), .CI(\SUMB[20][45] ), 
        .CO(\CARRYB[21][44] ), .S(\SUMB[21][44] ) );
  FA1A S2_20_43 ( .A(\ab[20][43] ), .B(\CARRYB[19][43] ), .CI(\SUMB[19][44] ), 
        .CO(\CARRYB[20][43] ), .S(\SUMB[20][43] ) );
  FA1A S2_19_43 ( .A(\ab[19][43] ), .B(\CARRYB[18][43] ), .CI(\SUMB[18][44] ), 
        .CO(\CARRYB[19][43] ), .S(\SUMB[19][43] ) );
  FA1A S2_18_43 ( .A(\ab[18][43] ), .B(\CARRYB[17][43] ), .CI(\SUMB[17][44] ), 
        .CO(\CARRYB[18][43] ), .S(\SUMB[18][43] ) );
  FA1A S2_17_43 ( .A(\ab[17][43] ), .B(\CARRYB[16][43] ), .CI(\SUMB[16][44] ), 
        .CO(\CARRYB[17][43] ), .S(\SUMB[17][43] ) );
  FA1A S2_16_43 ( .A(\ab[16][43] ), .B(\CARRYB[15][43] ), .CI(\SUMB[15][44] ), 
        .CO(\CARRYB[16][43] ), .S(\SUMB[16][43] ) );
  FA1A S2_15_43 ( .A(\ab[15][43] ), .B(\CARRYB[14][43] ), .CI(\SUMB[14][44] ), 
        .CO(\CARRYB[15][43] ), .S(\SUMB[15][43] ) );
  FA1A S2_14_43 ( .A(\ab[14][43] ), .B(\CARRYB[13][43] ), .CI(\SUMB[13][44] ), 
        .CO(\CARRYB[14][43] ), .S(\SUMB[14][43] ) );
  FA1A S2_13_43 ( .A(\ab[13][43] ), .B(\CARRYB[12][43] ), .CI(\SUMB[12][44] ), 
        .CO(\CARRYB[13][43] ), .S(\SUMB[13][43] ) );
  FA1A S2_12_43 ( .A(\ab[12][43] ), .B(\CARRYB[11][43] ), .CI(\SUMB[11][44] ), 
        .CO(\CARRYB[12][43] ), .S(\SUMB[12][43] ) );
  FA1A S2_11_43 ( .A(\ab[11][43] ), .B(\CARRYB[10][43] ), .CI(\SUMB[10][44] ), 
        .CO(\CARRYB[11][43] ), .S(\SUMB[11][43] ) );
  FA1A S2_10_43 ( .A(\ab[10][43] ), .B(\CARRYB[9][43] ), .CI(\SUMB[9][44] ), 
        .CO(\CARRYB[10][43] ), .S(\SUMB[10][43] ) );
  FA1A S2_9_43 ( .A(\ab[9][43] ), .B(\CARRYB[8][43] ), .CI(\SUMB[8][44] ), 
        .CO(\CARRYB[9][43] ), .S(\SUMB[9][43] ) );
  FA1A S2_8_43 ( .A(\ab[8][43] ), .B(\CARRYB[7][43] ), .CI(\SUMB[7][44] ), 
        .CO(\CARRYB[8][43] ), .S(\SUMB[8][43] ) );
  FA1A S2_7_43 ( .A(\ab[7][43] ), .B(\CARRYB[6][43] ), .CI(\SUMB[6][44] ), 
        .CO(\CARRYB[7][43] ), .S(\SUMB[7][43] ) );
  FA1A S2_6_43 ( .A(\ab[6][43] ), .B(\CARRYB[5][43] ), .CI(\SUMB[5][44] ), 
        .CO(\CARRYB[6][43] ), .S(\SUMB[6][43] ) );
  FA1A S2_5_43 ( .A(\ab[5][43] ), .B(\CARRYB[4][43] ), .CI(\SUMB[4][44] ), 
        .CO(\CARRYB[5][43] ), .S(\SUMB[5][43] ) );
  FA1A S2_4_43 ( .A(\ab[4][43] ), .B(\CARRYB[3][43] ), .CI(\SUMB[3][44] ), 
        .CO(\CARRYB[4][43] ), .S(\SUMB[4][43] ) );
  FA1A S2_3_43 ( .A(\ab[3][43] ), .B(\CARRYB[2][43] ), .CI(\SUMB[2][44] ), 
        .CO(\CARRYB[3][43] ), .S(\SUMB[3][43] ) );
  FA1A S2_2_43 ( .A(\ab[2][43] ), .B(\CARRYB[1][43] ), .CI(\SUMB[1][44] ), 
        .CO(\CARRYB[2][43] ), .S(\SUMB[2][43] ) );
  FA1A S4_43 ( .A(\ab[21][43] ), .B(\CARRYB[20][43] ), .CI(\SUMB[20][44] ), 
        .CO(\CARRYB[21][43] ), .S(\SUMB[21][43] ) );
  FA1A S4_42 ( .A(\ab[21][42] ), .B(\CARRYB[20][42] ), .CI(\SUMB[20][43] ), 
        .CO(\CARRYB[21][42] ), .S(\SUMB[21][42] ) );
  FA1A S2_20_42 ( .A(\ab[20][42] ), .B(\CARRYB[19][42] ), .CI(\SUMB[19][43] ), 
        .CO(\CARRYB[20][42] ), .S(\SUMB[20][42] ) );
  FA1A S2_19_42 ( .A(\ab[19][42] ), .B(\CARRYB[18][42] ), .CI(\SUMB[18][43] ), 
        .CO(\CARRYB[19][42] ), .S(\SUMB[19][42] ) );
  FA1A S2_18_42 ( .A(\ab[18][42] ), .B(\CARRYB[17][42] ), .CI(\SUMB[17][43] ), 
        .CO(\CARRYB[18][42] ), .S(\SUMB[18][42] ) );
  FA1A S2_17_42 ( .A(\ab[17][42] ), .B(\CARRYB[16][42] ), .CI(\SUMB[16][43] ), 
        .CO(\CARRYB[17][42] ), .S(\SUMB[17][42] ) );
  FA1A S2_16_42 ( .A(\ab[16][42] ), .B(\CARRYB[15][42] ), .CI(\SUMB[15][43] ), 
        .CO(\CARRYB[16][42] ), .S(\SUMB[16][42] ) );
  FA1A S2_15_42 ( .A(\ab[15][42] ), .B(\CARRYB[14][42] ), .CI(\SUMB[14][43] ), 
        .CO(\CARRYB[15][42] ), .S(\SUMB[15][42] ) );
  FA1A S2_14_42 ( .A(\ab[14][42] ), .B(\CARRYB[13][42] ), .CI(\SUMB[13][43] ), 
        .CO(\CARRYB[14][42] ), .S(\SUMB[14][42] ) );
  FA1A S2_13_42 ( .A(\ab[13][42] ), .B(\CARRYB[12][42] ), .CI(\SUMB[12][43] ), 
        .CO(\CARRYB[13][42] ), .S(\SUMB[13][42] ) );
  FA1A S2_12_42 ( .A(\ab[12][42] ), .B(\CARRYB[11][42] ), .CI(\SUMB[11][43] ), 
        .CO(\CARRYB[12][42] ), .S(\SUMB[12][42] ) );
  FA1A S2_11_42 ( .A(\ab[11][42] ), .B(\CARRYB[10][42] ), .CI(\SUMB[10][43] ), 
        .CO(\CARRYB[11][42] ), .S(\SUMB[11][42] ) );
  FA1A S2_10_42 ( .A(\ab[10][42] ), .B(\CARRYB[9][42] ), .CI(\SUMB[9][43] ), 
        .CO(\CARRYB[10][42] ), .S(\SUMB[10][42] ) );
  FA1A S2_9_42 ( .A(\ab[9][42] ), .B(\CARRYB[8][42] ), .CI(\SUMB[8][43] ), 
        .CO(\CARRYB[9][42] ), .S(\SUMB[9][42] ) );
  FA1A S2_8_42 ( .A(\ab[8][42] ), .B(\CARRYB[7][42] ), .CI(\SUMB[7][43] ), 
        .CO(\CARRYB[8][42] ), .S(\SUMB[8][42] ) );
  FA1A S2_7_42 ( .A(\ab[7][42] ), .B(\CARRYB[6][42] ), .CI(\SUMB[6][43] ), 
        .CO(\CARRYB[7][42] ), .S(\SUMB[7][42] ) );
  FA1A S2_6_42 ( .A(\ab[6][42] ), .B(\CARRYB[5][42] ), .CI(\SUMB[5][43] ), 
        .CO(\CARRYB[6][42] ), .S(\SUMB[6][42] ) );
  FA1A S2_5_42 ( .A(\ab[5][42] ), .B(\CARRYB[4][42] ), .CI(\SUMB[4][43] ), 
        .CO(\CARRYB[5][42] ), .S(\SUMB[5][42] ) );
  FA1A S2_4_42 ( .A(\ab[4][42] ), .B(\CARRYB[3][42] ), .CI(\SUMB[3][43] ), 
        .CO(\CARRYB[4][42] ), .S(\SUMB[4][42] ) );
  FA1A S2_3_42 ( .A(\ab[3][42] ), .B(\CARRYB[2][42] ), .CI(\SUMB[2][43] ), 
        .CO(\CARRYB[3][42] ), .S(\SUMB[3][42] ) );
  FA1A S2_2_42 ( .A(\ab[2][42] ), .B(\CARRYB[1][42] ), .CI(\SUMB[1][43] ), 
        .CO(\CARRYB[2][42] ), .S(\SUMB[2][42] ) );
  FA1A S2_20_41 ( .A(\ab[20][41] ), .B(\CARRYB[19][41] ), .CI(\SUMB[19][42] ), 
        .CO(\CARRYB[20][41] ), .S(\SUMB[20][41] ) );
  FA1A S2_19_41 ( .A(\ab[19][41] ), .B(\CARRYB[18][41] ), .CI(\SUMB[18][42] ), 
        .CO(\CARRYB[19][41] ), .S(\SUMB[19][41] ) );
  FA1A S2_18_41 ( .A(\ab[18][41] ), .B(\CARRYB[17][41] ), .CI(\SUMB[17][42] ), 
        .CO(\CARRYB[18][41] ), .S(\SUMB[18][41] ) );
  FA1A S2_17_41 ( .A(\ab[17][41] ), .B(\CARRYB[16][41] ), .CI(\SUMB[16][42] ), 
        .CO(\CARRYB[17][41] ), .S(\SUMB[17][41] ) );
  FA1A S2_16_41 ( .A(\ab[16][41] ), .B(\CARRYB[15][41] ), .CI(\SUMB[15][42] ), 
        .CO(\CARRYB[16][41] ), .S(\SUMB[16][41] ) );
  FA1A S2_15_41 ( .A(\ab[15][41] ), .B(\CARRYB[14][41] ), .CI(\SUMB[14][42] ), 
        .CO(\CARRYB[15][41] ), .S(\SUMB[15][41] ) );
  FA1A S2_14_41 ( .A(\ab[14][41] ), .B(\CARRYB[13][41] ), .CI(\SUMB[13][42] ), 
        .CO(\CARRYB[14][41] ), .S(\SUMB[14][41] ) );
  FA1A S2_13_41 ( .A(\ab[13][41] ), .B(\CARRYB[12][41] ), .CI(\SUMB[12][42] ), 
        .CO(\CARRYB[13][41] ), .S(\SUMB[13][41] ) );
  FA1A S2_12_41 ( .A(\ab[12][41] ), .B(\CARRYB[11][41] ), .CI(\SUMB[11][42] ), 
        .CO(\CARRYB[12][41] ), .S(\SUMB[12][41] ) );
  FA1A S2_11_41 ( .A(\ab[11][41] ), .B(\CARRYB[10][41] ), .CI(\SUMB[10][42] ), 
        .CO(\CARRYB[11][41] ), .S(\SUMB[11][41] ) );
  FA1A S2_10_41 ( .A(\ab[10][41] ), .B(\CARRYB[9][41] ), .CI(\SUMB[9][42] ), 
        .CO(\CARRYB[10][41] ), .S(\SUMB[10][41] ) );
  FA1A S2_9_41 ( .A(\ab[9][41] ), .B(\CARRYB[8][41] ), .CI(\SUMB[8][42] ), 
        .CO(\CARRYB[9][41] ), .S(\SUMB[9][41] ) );
  FA1A S2_8_41 ( .A(\ab[8][41] ), .B(\CARRYB[7][41] ), .CI(\SUMB[7][42] ), 
        .CO(\CARRYB[8][41] ), .S(\SUMB[8][41] ) );
  FA1A S2_7_41 ( .A(\ab[7][41] ), .B(\CARRYB[6][41] ), .CI(\SUMB[6][42] ), 
        .CO(\CARRYB[7][41] ), .S(\SUMB[7][41] ) );
  FA1A S2_6_41 ( .A(\ab[6][41] ), .B(\CARRYB[5][41] ), .CI(\SUMB[5][42] ), 
        .CO(\CARRYB[6][41] ), .S(\SUMB[6][41] ) );
  FA1A S2_5_41 ( .A(\ab[5][41] ), .B(\CARRYB[4][41] ), .CI(\SUMB[4][42] ), 
        .CO(\CARRYB[5][41] ), .S(\SUMB[5][41] ) );
  FA1A S2_4_41 ( .A(\ab[4][41] ), .B(\CARRYB[3][41] ), .CI(\SUMB[3][42] ), 
        .CO(\CARRYB[4][41] ), .S(\SUMB[4][41] ) );
  FA1A S2_3_41 ( .A(\ab[3][41] ), .B(\CARRYB[2][41] ), .CI(\SUMB[2][42] ), 
        .CO(\CARRYB[3][41] ), .S(\SUMB[3][41] ) );
  FA1A S4_41 ( .A(\ab[21][41] ), .B(\CARRYB[20][41] ), .CI(\SUMB[20][42] ), 
        .CO(\CARRYB[21][41] ), .S(\SUMB[21][41] ) );
  FA1A S2_20_40 ( .A(\ab[20][40] ), .B(\CARRYB[19][40] ), .CI(\SUMB[19][41] ), 
        .CO(\CARRYB[20][40] ), .S(\SUMB[20][40] ) );
  FA1A S2_19_40 ( .A(\ab[19][40] ), .B(\CARRYB[18][40] ), .CI(\SUMB[18][41] ), 
        .CO(\CARRYB[19][40] ), .S(\SUMB[19][40] ) );
  FA1A S2_18_40 ( .A(\ab[18][40] ), .B(\CARRYB[17][40] ), .CI(\SUMB[17][41] ), 
        .CO(\CARRYB[18][40] ), .S(\SUMB[18][40] ) );
  FA1A S2_17_40 ( .A(\ab[17][40] ), .B(\CARRYB[16][40] ), .CI(\SUMB[16][41] ), 
        .CO(\CARRYB[17][40] ), .S(\SUMB[17][40] ) );
  FA1A S2_16_40 ( .A(\ab[16][40] ), .B(\CARRYB[15][40] ), .CI(\SUMB[15][41] ), 
        .CO(\CARRYB[16][40] ), .S(\SUMB[16][40] ) );
  FA1A S2_15_40 ( .A(\ab[15][40] ), .B(\CARRYB[14][40] ), .CI(\SUMB[14][41] ), 
        .CO(\CARRYB[15][40] ), .S(\SUMB[15][40] ) );
  FA1A S2_14_40 ( .A(\ab[14][40] ), .B(\CARRYB[13][40] ), .CI(\SUMB[13][41] ), 
        .CO(\CARRYB[14][40] ), .S(\SUMB[14][40] ) );
  FA1A S2_13_40 ( .A(\ab[13][40] ), .B(\CARRYB[12][40] ), .CI(\SUMB[12][41] ), 
        .CO(\CARRYB[13][40] ), .S(\SUMB[13][40] ) );
  FA1A S2_12_40 ( .A(\ab[12][40] ), .B(\CARRYB[11][40] ), .CI(\SUMB[11][41] ), 
        .CO(\CARRYB[12][40] ), .S(\SUMB[12][40] ) );
  FA1A S2_11_40 ( .A(\ab[11][40] ), .B(\CARRYB[10][40] ), .CI(\SUMB[10][41] ), 
        .CO(\CARRYB[11][40] ), .S(\SUMB[11][40] ) );
  FA1A S2_10_40 ( .A(\ab[10][40] ), .B(\CARRYB[9][40] ), .CI(\SUMB[9][41] ), 
        .CO(\CARRYB[10][40] ), .S(\SUMB[10][40] ) );
  FA1A S2_9_40 ( .A(\ab[9][40] ), .B(\CARRYB[8][40] ), .CI(\SUMB[8][41] ), 
        .CO(\CARRYB[9][40] ), .S(\SUMB[9][40] ) );
  FA1A S2_8_40 ( .A(\ab[8][40] ), .B(\CARRYB[7][40] ), .CI(\SUMB[7][41] ), 
        .CO(\CARRYB[8][40] ), .S(\SUMB[8][40] ) );
  FA1A S2_7_40 ( .A(\ab[7][40] ), .B(\CARRYB[6][40] ), .CI(\SUMB[6][41] ), 
        .CO(\CARRYB[7][40] ), .S(\SUMB[7][40] ) );
  FA1A S2_6_40 ( .A(\ab[6][40] ), .B(\CARRYB[5][40] ), .CI(\SUMB[5][41] ), 
        .CO(\CARRYB[6][40] ), .S(\SUMB[6][40] ) );
  FA1A S2_5_40 ( .A(\ab[5][40] ), .B(\CARRYB[4][40] ), .CI(\SUMB[4][41] ), 
        .CO(\CARRYB[5][40] ), .S(\SUMB[5][40] ) );
  FA1A S2_4_40 ( .A(\ab[4][40] ), .B(\CARRYB[3][40] ), .CI(\SUMB[3][41] ), 
        .CO(\CARRYB[4][40] ), .S(\SUMB[4][40] ) );
  FA1A S2_2_41 ( .A(\ab[2][41] ), .B(\CARRYB[1][41] ), .CI(\SUMB[1][42] ), 
        .CO(\CARRYB[2][41] ), .S(\SUMB[2][41] ) );
  FA1A S4_40 ( .A(\ab[21][40] ), .B(\CARRYB[20][40] ), .CI(\SUMB[20][41] ), 
        .CO(\CARRYB[21][40] ), .S(\SUMB[21][40] ) );
  FA1A S2_20_39 ( .A(\ab[20][39] ), .B(\CARRYB[19][39] ), .CI(\SUMB[19][40] ), 
        .CO(\CARRYB[20][39] ), .S(\SUMB[20][39] ) );
  FA1A S2_19_39 ( .A(\ab[19][39] ), .B(\CARRYB[18][39] ), .CI(\SUMB[18][40] ), 
        .CO(\CARRYB[19][39] ), .S(\SUMB[19][39] ) );
  FA1A S2_18_39 ( .A(\ab[18][39] ), .B(\CARRYB[17][39] ), .CI(\SUMB[17][40] ), 
        .CO(\CARRYB[18][39] ), .S(\SUMB[18][39] ) );
  FA1A S2_17_39 ( .A(\ab[17][39] ), .B(\CARRYB[16][39] ), .CI(\SUMB[16][40] ), 
        .CO(\CARRYB[17][39] ), .S(\SUMB[17][39] ) );
  FA1A S2_16_39 ( .A(\ab[16][39] ), .B(\CARRYB[15][39] ), .CI(\SUMB[15][40] ), 
        .CO(\CARRYB[16][39] ), .S(\SUMB[16][39] ) );
  FA1A S2_15_39 ( .A(\ab[15][39] ), .B(\CARRYB[14][39] ), .CI(\SUMB[14][40] ), 
        .CO(\CARRYB[15][39] ), .S(\SUMB[15][39] ) );
  FA1A S2_14_39 ( .A(\ab[14][39] ), .B(\CARRYB[13][39] ), .CI(\SUMB[13][40] ), 
        .CO(\CARRYB[14][39] ), .S(\SUMB[14][39] ) );
  FA1A S2_13_39 ( .A(\ab[13][39] ), .B(\CARRYB[12][39] ), .CI(\SUMB[12][40] ), 
        .CO(\CARRYB[13][39] ), .S(\SUMB[13][39] ) );
  FA1A S2_12_39 ( .A(\ab[12][39] ), .B(\CARRYB[11][39] ), .CI(\SUMB[11][40] ), 
        .CO(\CARRYB[12][39] ), .S(\SUMB[12][39] ) );
  FA1A S2_11_39 ( .A(\ab[11][39] ), .B(\CARRYB[10][39] ), .CI(\SUMB[10][40] ), 
        .CO(\CARRYB[11][39] ), .S(\SUMB[11][39] ) );
  FA1A S2_10_39 ( .A(\ab[10][39] ), .B(\CARRYB[9][39] ), .CI(\SUMB[9][40] ), 
        .CO(\CARRYB[10][39] ), .S(\SUMB[10][39] ) );
  FA1A S2_9_39 ( .A(\ab[9][39] ), .B(\CARRYB[8][39] ), .CI(\SUMB[8][40] ), 
        .CO(\CARRYB[9][39] ), .S(\SUMB[9][39] ) );
  FA1A S2_8_39 ( .A(\ab[8][39] ), .B(\CARRYB[7][39] ), .CI(\SUMB[7][40] ), 
        .CO(\CARRYB[8][39] ), .S(\SUMB[8][39] ) );
  FA1A S2_7_39 ( .A(\ab[7][39] ), .B(\CARRYB[6][39] ), .CI(\SUMB[6][40] ), 
        .CO(\CARRYB[7][39] ), .S(\SUMB[7][39] ) );
  FA1A S2_6_39 ( .A(\ab[6][39] ), .B(\CARRYB[5][39] ), .CI(\SUMB[5][40] ), 
        .CO(\CARRYB[6][39] ), .S(\SUMB[6][39] ) );
  FA1A S2_5_39 ( .A(\ab[5][39] ), .B(\CARRYB[4][39] ), .CI(\SUMB[4][40] ), 
        .CO(\CARRYB[5][39] ), .S(\SUMB[5][39] ) );
  FA1A S2_4_39 ( .A(\ab[4][39] ), .B(\CARRYB[3][39] ), .CI(\SUMB[3][40] ), 
        .CO(\CARRYB[4][39] ), .S(\SUMB[4][39] ) );
  FA1A S2_3_40 ( .A(\ab[3][40] ), .B(\CARRYB[2][40] ), .CI(\SUMB[2][41] ), 
        .CO(\CARRYB[3][40] ), .S(\SUMB[3][40] ) );
  FA1A S2_3_39 ( .A(\ab[3][39] ), .B(\CARRYB[2][39] ), .CI(\SUMB[2][40] ), 
        .CO(\CARRYB[3][39] ), .S(\SUMB[3][39] ) );
  FA1A S2_2_40 ( .A(\ab[2][40] ), .B(\CARRYB[1][40] ), .CI(\SUMB[1][41] ), 
        .CO(\CARRYB[2][40] ), .S(\SUMB[2][40] ) );
  FA1A S2_2_39 ( .A(\ab[2][39] ), .B(\CARRYB[1][39] ), .CI(\SUMB[1][40] ), 
        .CO(\CARRYB[2][39] ), .S(\SUMB[2][39] ) );
  FA1A S4_39 ( .A(\ab[21][39] ), .B(\CARRYB[20][39] ), .CI(\SUMB[20][40] ), 
        .CO(\CARRYB[21][39] ), .S(\SUMB[21][39] ) );
  FA1A S4_36 ( .A(\ab[21][36] ), .B(\CARRYB[20][36] ), .CI(\SUMB[20][37] ), 
        .CO(\CARRYB[21][36] ), .S(\SUMB[21][36] ) );
  FA1A S2_20_36 ( .A(\ab[20][36] ), .B(\CARRYB[19][36] ), .CI(\SUMB[19][37] ), 
        .CO(\CARRYB[20][36] ), .S(\SUMB[20][36] ) );
  FA1A S2_19_36 ( .A(\ab[19][36] ), .B(\CARRYB[18][36] ), .CI(\SUMB[18][37] ), 
        .CO(\CARRYB[19][36] ), .S(\SUMB[19][36] ) );
  FA1A S4_37 ( .A(\ab[21][37] ), .B(\CARRYB[20][37] ), .CI(\SUMB[20][38] ), 
        .CO(\CARRYB[21][37] ), .S(\SUMB[21][37] ) );
  FA1A S2_18_36 ( .A(\ab[18][36] ), .B(\CARRYB[17][36] ), .CI(\SUMB[17][37] ), 
        .CO(\CARRYB[18][36] ), .S(\SUMB[18][36] ) );
  FA1A S2_20_38 ( .A(\ab[20][38] ), .B(\CARRYB[19][38] ), .CI(\SUMB[19][39] ), 
        .CO(\CARRYB[20][38] ), .S(\SUMB[20][38] ) );
  FA1A S2_20_37 ( .A(\ab[20][37] ), .B(\CARRYB[19][37] ), .CI(\SUMB[19][38] ), 
        .CO(\CARRYB[20][37] ), .S(\SUMB[20][37] ) );
  FA1A S2_17_36 ( .A(\ab[17][36] ), .B(\CARRYB[16][36] ), .CI(\SUMB[16][37] ), 
        .CO(\CARRYB[17][36] ), .S(\SUMB[17][36] ) );
  FA1A S2_19_38 ( .A(\ab[19][38] ), .B(\CARRYB[18][38] ), .CI(\SUMB[18][39] ), 
        .CO(\CARRYB[19][38] ), .S(\SUMB[19][38] ) );
  FA1A S2_19_37 ( .A(\ab[19][37] ), .B(\CARRYB[18][37] ), .CI(\SUMB[18][38] ), 
        .CO(\CARRYB[19][37] ), .S(\SUMB[19][37] ) );
  FA1A S2_18_38 ( .A(\ab[18][38] ), .B(\CARRYB[17][38] ), .CI(\SUMB[17][39] ), 
        .CO(\CARRYB[18][38] ), .S(\SUMB[18][38] ) );
  FA1A S2_18_37 ( .A(\ab[18][37] ), .B(\CARRYB[17][37] ), .CI(\SUMB[17][38] ), 
        .CO(\CARRYB[18][37] ), .S(\SUMB[18][37] ) );
  FA1A S2_17_38 ( .A(\ab[17][38] ), .B(\CARRYB[16][38] ), .CI(\SUMB[16][39] ), 
        .CO(\CARRYB[17][38] ), .S(\SUMB[17][38] ) );
  FA1A S2_17_37 ( .A(\ab[17][37] ), .B(\CARRYB[16][37] ), .CI(\SUMB[16][38] ), 
        .CO(\CARRYB[17][37] ), .S(\SUMB[17][37] ) );
  FA1A S2_16_38 ( .A(\ab[16][38] ), .B(\CARRYB[15][38] ), .CI(\SUMB[15][39] ), 
        .CO(\CARRYB[16][38] ), .S(\SUMB[16][38] ) );
  FA1A S2_16_37 ( .A(\ab[16][37] ), .B(\CARRYB[15][37] ), .CI(\SUMB[15][38] ), 
        .CO(\CARRYB[16][37] ), .S(\SUMB[16][37] ) );
  FA1A S2_16_36 ( .A(\ab[16][36] ), .B(\CARRYB[15][36] ), .CI(\SUMB[15][37] ), 
        .CO(\CARRYB[16][36] ), .S(\SUMB[16][36] ) );
  FA1A S2_15_38 ( .A(\ab[15][38] ), .B(\CARRYB[14][38] ), .CI(\SUMB[14][39] ), 
        .CO(\CARRYB[15][38] ), .S(\SUMB[15][38] ) );
  FA1A S2_15_37 ( .A(\ab[15][37] ), .B(\CARRYB[14][37] ), .CI(\SUMB[14][38] ), 
        .CO(\CARRYB[15][37] ), .S(\SUMB[15][37] ) );
  FA1A S2_15_36 ( .A(\ab[15][36] ), .B(\CARRYB[14][36] ), .CI(\SUMB[14][37] ), 
        .CO(\CARRYB[15][36] ), .S(\SUMB[15][36] ) );
  FA1A S2_14_38 ( .A(\ab[14][38] ), .B(\CARRYB[13][38] ), .CI(\SUMB[13][39] ), 
        .CO(\CARRYB[14][38] ), .S(\SUMB[14][38] ) );
  FA1A S2_14_37 ( .A(\ab[14][37] ), .B(\CARRYB[13][37] ), .CI(\SUMB[13][38] ), 
        .CO(\CARRYB[14][37] ), .S(\SUMB[14][37] ) );
  FA1A S2_14_36 ( .A(\ab[14][36] ), .B(\CARRYB[13][36] ), .CI(\SUMB[13][37] ), 
        .CO(\CARRYB[14][36] ), .S(\SUMB[14][36] ) );
  FA1A S2_13_38 ( .A(\ab[13][38] ), .B(\CARRYB[12][38] ), .CI(\SUMB[12][39] ), 
        .CO(\CARRYB[13][38] ), .S(\SUMB[13][38] ) );
  FA1A S2_13_37 ( .A(\ab[13][37] ), .B(\CARRYB[12][37] ), .CI(\SUMB[12][38] ), 
        .CO(\CARRYB[13][37] ), .S(\SUMB[13][37] ) );
  FA1A S2_12_38 ( .A(\ab[12][38] ), .B(\CARRYB[11][38] ), .CI(\SUMB[11][39] ), 
        .CO(\CARRYB[12][38] ), .S(\SUMB[12][38] ) );
  FA1A S2_13_36 ( .A(\ab[13][36] ), .B(\CARRYB[12][36] ), .CI(\SUMB[12][37] ), 
        .CO(\CARRYB[13][36] ), .S(\SUMB[13][36] ) );
  FA1A S2_12_37 ( .A(\ab[12][37] ), .B(\CARRYB[11][37] ), .CI(\SUMB[11][38] ), 
        .CO(\CARRYB[12][37] ), .S(\SUMB[12][37] ) );
  FA1A S2_12_36 ( .A(\ab[12][36] ), .B(\CARRYB[11][36] ), .CI(\SUMB[11][37] ), 
        .CO(\CARRYB[12][36] ), .S(\SUMB[12][36] ) );
  FA1A S2_11_38 ( .A(\ab[11][38] ), .B(\CARRYB[10][38] ), .CI(\SUMB[10][39] ), 
        .CO(\CARRYB[11][38] ), .S(\SUMB[11][38] ) );
  FA1A S2_11_37 ( .A(\ab[11][37] ), .B(\CARRYB[10][37] ), .CI(\SUMB[10][38] ), 
        .CO(\CARRYB[11][37] ), .S(\SUMB[11][37] ) );
  FA1A S2_11_36 ( .A(\ab[11][36] ), .B(\CARRYB[10][36] ), .CI(\SUMB[10][37] ), 
        .CO(\CARRYB[11][36] ), .S(\SUMB[11][36] ) );
  FA1A S2_10_38 ( .A(\ab[10][38] ), .B(\CARRYB[9][38] ), .CI(\SUMB[9][39] ), 
        .CO(\CARRYB[10][38] ), .S(\SUMB[10][38] ) );
  FA1A S2_10_37 ( .A(\ab[10][37] ), .B(\CARRYB[9][37] ), .CI(\SUMB[9][38] ), 
        .CO(\CARRYB[10][37] ), .S(\SUMB[10][37] ) );
  FA1A S2_10_36 ( .A(\ab[10][36] ), .B(\CARRYB[9][36] ), .CI(\SUMB[9][37] ), 
        .CO(\CARRYB[10][36] ), .S(\SUMB[10][36] ) );
  FA1A S2_9_38 ( .A(\ab[9][38] ), .B(\CARRYB[8][38] ), .CI(\SUMB[8][39] ), 
        .CO(\CARRYB[9][38] ), .S(\SUMB[9][38] ) );
  FA1A S2_9_37 ( .A(\ab[9][37] ), .B(\CARRYB[8][37] ), .CI(\SUMB[8][38] ), 
        .CO(\CARRYB[9][37] ), .S(\SUMB[9][37] ) );
  FA1A S2_9_36 ( .A(\ab[9][36] ), .B(\CARRYB[8][36] ), .CI(\SUMB[8][37] ), 
        .CO(\CARRYB[9][36] ), .S(\SUMB[9][36] ) );
  FA1A S2_8_38 ( .A(\ab[8][38] ), .B(\CARRYB[7][38] ), .CI(\SUMB[7][39] ), 
        .CO(\CARRYB[8][38] ), .S(\SUMB[8][38] ) );
  FA1A S2_8_37 ( .A(\ab[8][37] ), .B(\CARRYB[7][37] ), .CI(\SUMB[7][38] ), 
        .CO(\CARRYB[8][37] ), .S(\SUMB[8][37] ) );
  FA1A S2_8_36 ( .A(\ab[8][36] ), .B(\CARRYB[7][36] ), .CI(\SUMB[7][37] ), 
        .CO(\CARRYB[8][36] ), .S(\SUMB[8][36] ) );
  FA1A S2_7_38 ( .A(\ab[7][38] ), .B(\CARRYB[6][38] ), .CI(\SUMB[6][39] ), 
        .CO(\CARRYB[7][38] ), .S(\SUMB[7][38] ) );
  FA1A S2_7_37 ( .A(\ab[7][37] ), .B(\CARRYB[6][37] ), .CI(\SUMB[6][38] ), 
        .CO(\CARRYB[7][37] ), .S(\SUMB[7][37] ) );
  FA1A S2_7_36 ( .A(\ab[7][36] ), .B(\CARRYB[6][36] ), .CI(\SUMB[6][37] ), 
        .CO(\CARRYB[7][36] ), .S(\SUMB[7][36] ) );
  FA1A S2_6_38 ( .A(\ab[6][38] ), .B(\CARRYB[5][38] ), .CI(\SUMB[5][39] ), 
        .CO(\CARRYB[6][38] ), .S(\SUMB[6][38] ) );
  FA1A S2_6_37 ( .A(\ab[6][37] ), .B(\CARRYB[5][37] ), .CI(\SUMB[5][38] ), 
        .CO(\CARRYB[6][37] ), .S(\SUMB[6][37] ) );
  FA1A S2_6_36 ( .A(\ab[6][36] ), .B(\CARRYB[5][36] ), .CI(\SUMB[5][37] ), 
        .CO(\CARRYB[6][36] ), .S(\SUMB[6][36] ) );
  FA1A S2_5_38 ( .A(\ab[5][38] ), .B(\CARRYB[4][38] ), .CI(\SUMB[4][39] ), 
        .CO(\CARRYB[5][38] ), .S(\SUMB[5][38] ) );
  FA1A S2_5_37 ( .A(\ab[5][37] ), .B(\CARRYB[4][37] ), .CI(\SUMB[4][38] ), 
        .CO(\CARRYB[5][37] ), .S(\SUMB[5][37] ) );
  FA1A S2_5_36 ( .A(\ab[5][36] ), .B(\CARRYB[4][36] ), .CI(\SUMB[4][37] ), 
        .CO(\CARRYB[5][36] ), .S(\SUMB[5][36] ) );
  FA1A S2_4_38 ( .A(\ab[4][38] ), .B(\CARRYB[3][38] ), .CI(\SUMB[3][39] ), 
        .CO(\CARRYB[4][38] ), .S(\SUMB[4][38] ) );
  FA1A S2_4_37 ( .A(\ab[4][37] ), .B(\CARRYB[3][37] ), .CI(\SUMB[3][38] ), 
        .CO(\CARRYB[4][37] ), .S(\SUMB[4][37] ) );
  FA1A S2_4_36 ( .A(\ab[4][36] ), .B(\CARRYB[3][36] ), .CI(\SUMB[3][37] ), 
        .CO(\CARRYB[4][36] ), .S(\SUMB[4][36] ) );
  FA1A S2_3_38 ( .A(\ab[3][38] ), .B(\CARRYB[2][38] ), .CI(\SUMB[2][39] ), 
        .CO(\CARRYB[3][38] ), .S(\SUMB[3][38] ) );
  FA1A S2_3_37 ( .A(\ab[3][37] ), .B(\CARRYB[2][37] ), .CI(\SUMB[2][38] ), 
        .CO(\CARRYB[3][37] ), .S(\SUMB[3][37] ) );
  FA1A S2_3_36 ( .A(\ab[3][36] ), .B(\CARRYB[2][36] ), .CI(\SUMB[2][37] ), 
        .CO(\CARRYB[3][36] ), .S(\SUMB[3][36] ) );
  FA1A S2_2_38 ( .A(\ab[2][38] ), .B(\CARRYB[1][38] ), .CI(\SUMB[1][39] ), 
        .CO(\CARRYB[2][38] ), .S(\SUMB[2][38] ) );
  FA1A S2_2_37 ( .A(\ab[2][37] ), .B(\CARRYB[1][37] ), .CI(\SUMB[1][38] ), 
        .CO(\CARRYB[2][37] ), .S(\SUMB[2][37] ) );
  FA1A S2_2_36 ( .A(\ab[2][36] ), .B(\CARRYB[1][36] ), .CI(\SUMB[1][37] ), 
        .CO(\CARRYB[2][36] ), .S(\SUMB[2][36] ) );
  FA1A S4_38 ( .A(\ab[21][38] ), .B(\CARRYB[20][38] ), .CI(\SUMB[20][39] ), 
        .CO(\CARRYB[21][38] ), .S(\SUMB[21][38] ) );
  FA1A S4_33 ( .A(\ab[21][33] ), .B(\CARRYB[20][33] ), .CI(\SUMB[20][34] ), 
        .CO(\CARRYB[21][33] ), .S(\SUMB[21][33] ) );
  FA1A S4_32 ( .A(\ab[21][32] ), .B(\CARRYB[20][32] ), .CI(\SUMB[20][33] ), 
        .CO(\CARRYB[21][32] ), .S(\SUMB[21][32] ) );
  FA1A S2_20_34 ( .A(\ab[20][34] ), .B(\CARRYB[19][34] ), .CI(\SUMB[19][35] ), 
        .CO(\CARRYB[20][34] ), .S(\SUMB[20][34] ) );
  FA1A S2_20_33 ( .A(\ab[20][33] ), .B(\CARRYB[19][33] ), .CI(\SUMB[19][34] ), 
        .CO(\CARRYB[20][33] ), .S(\SUMB[20][33] ) );
  FA1A S2_19_34 ( .A(\ab[19][34] ), .B(\CARRYB[18][34] ), .CI(\SUMB[18][35] ), 
        .CO(\CARRYB[19][34] ), .S(\SUMB[19][34] ) );
  FA1A S2_20_35 ( .A(\ab[20][35] ), .B(\CARRYB[19][35] ), .CI(\SUMB[19][36] ), 
        .CO(\CARRYB[20][35] ), .S(\SUMB[20][35] ) );
  FA1A S2_19_35 ( .A(\ab[19][35] ), .B(\CARRYB[18][35] ), .CI(\SUMB[18][36] ), 
        .CO(\CARRYB[19][35] ), .S(\SUMB[19][35] ) );
  FA1A S2_18_35 ( .A(\ab[18][35] ), .B(\CARRYB[17][35] ), .CI(\SUMB[17][36] ), 
        .CO(\CARRYB[18][35] ), .S(\SUMB[18][35] ) );
  FA1A S2_20_32 ( .A(\ab[20][32] ), .B(\CARRYB[19][32] ), .CI(\SUMB[19][33] ), 
        .CO(\CARRYB[20][32] ), .S(\SUMB[20][32] ) );
  FA1A S2_19_33 ( .A(\ab[19][33] ), .B(\CARRYB[18][33] ), .CI(\SUMB[18][34] ), 
        .CO(\CARRYB[19][33] ), .S(\SUMB[19][33] ) );
  FA1A S2_19_32 ( .A(\ab[19][32] ), .B(\CARRYB[18][32] ), .CI(\SUMB[18][33] ), 
        .CO(\CARRYB[19][32] ), .S(\SUMB[19][32] ) );
  FA1A S2_18_34 ( .A(\ab[18][34] ), .B(\CARRYB[17][34] ), .CI(\SUMB[17][35] ), 
        .CO(\CARRYB[18][34] ), .S(\SUMB[18][34] ) );
  FA1A S2_18_33 ( .A(\ab[18][33] ), .B(\CARRYB[17][33] ), .CI(\SUMB[17][34] ), 
        .CO(\CARRYB[18][33] ), .S(\SUMB[18][33] ) );
  FA1A S2_18_32 ( .A(\ab[18][32] ), .B(\CARRYB[17][32] ), .CI(\SUMB[17][33] ), 
        .CO(\CARRYB[18][32] ), .S(\SUMB[18][32] ) );
  FA1A S2_17_35 ( .A(\ab[17][35] ), .B(\CARRYB[16][35] ), .CI(\SUMB[16][36] ), 
        .CO(\CARRYB[17][35] ), .S(\SUMB[17][35] ) );
  FA1A S2_17_34 ( .A(\ab[17][34] ), .B(\CARRYB[16][34] ), .CI(\SUMB[16][35] ), 
        .CO(\CARRYB[17][34] ), .S(\SUMB[17][34] ) );
  FA1A S2_17_33 ( .A(\ab[17][33] ), .B(\CARRYB[16][33] ), .CI(\SUMB[16][34] ), 
        .CO(\CARRYB[17][33] ), .S(\SUMB[17][33] ) );
  FA1A S2_16_35 ( .A(\ab[16][35] ), .B(\CARRYB[15][35] ), .CI(\SUMB[15][36] ), 
        .CO(\CARRYB[16][35] ), .S(\SUMB[16][35] ) );
  FA1A S2_16_34 ( .A(\ab[16][34] ), .B(\CARRYB[15][34] ), .CI(\SUMB[15][35] ), 
        .CO(\CARRYB[16][34] ), .S(\SUMB[16][34] ) );
  FA1A S2_17_32 ( .A(\ab[17][32] ), .B(\CARRYB[16][32] ), .CI(\SUMB[16][33] ), 
        .CO(\CARRYB[17][32] ), .S(\SUMB[17][32] ) );
  FA1A S2_15_35 ( .A(\ab[15][35] ), .B(\CARRYB[14][35] ), .CI(\SUMB[14][36] ), 
        .CO(\CARRYB[15][35] ), .S(\SUMB[15][35] ) );
  FA1A S2_16_33 ( .A(\ab[16][33] ), .B(\CARRYB[15][33] ), .CI(\SUMB[15][34] ), 
        .CO(\CARRYB[16][33] ), .S(\SUMB[16][33] ) );
  FA1A S2_16_32 ( .A(\ab[16][32] ), .B(\CARRYB[15][32] ), .CI(\SUMB[15][33] ), 
        .CO(\CARRYB[16][32] ), .S(\SUMB[16][32] ) );
  FA1A S2_15_34 ( .A(\ab[15][34] ), .B(\CARRYB[14][34] ), .CI(\SUMB[14][35] ), 
        .CO(\CARRYB[15][34] ), .S(\SUMB[15][34] ) );
  FA1A S2_15_33 ( .A(\ab[15][33] ), .B(\CARRYB[14][33] ), .CI(\SUMB[14][34] ), 
        .CO(\CARRYB[15][33] ), .S(\SUMB[15][33] ) );
  FA1A S2_15_32 ( .A(\ab[15][32] ), .B(\CARRYB[14][32] ), .CI(\SUMB[14][33] ), 
        .CO(\CARRYB[15][32] ), .S(\SUMB[15][32] ) );
  FA1A S2_14_35 ( .A(\ab[14][35] ), .B(\CARRYB[13][35] ), .CI(\SUMB[13][36] ), 
        .CO(\CARRYB[14][35] ), .S(\SUMB[14][35] ) );
  FA1A S2_14_34 ( .A(\ab[14][34] ), .B(\CARRYB[13][34] ), .CI(\SUMB[13][35] ), 
        .CO(\CARRYB[14][34] ), .S(\SUMB[14][34] ) );
  FA1A S2_14_33 ( .A(\ab[14][33] ), .B(\CARRYB[13][33] ), .CI(\SUMB[13][34] ), 
        .CO(\CARRYB[14][33] ), .S(\SUMB[14][33] ) );
  FA1A S2_14_32 ( .A(\ab[14][32] ), .B(\CARRYB[13][32] ), .CI(\SUMB[13][33] ), 
        .CO(\CARRYB[14][32] ), .S(\SUMB[14][32] ) );
  FA1A S2_13_35 ( .A(\ab[13][35] ), .B(\CARRYB[12][35] ), .CI(\SUMB[12][36] ), 
        .CO(\CARRYB[13][35] ), .S(\SUMB[13][35] ) );
  FA1A S2_13_34 ( .A(\ab[13][34] ), .B(\CARRYB[12][34] ), .CI(\SUMB[12][35] ), 
        .CO(\CARRYB[13][34] ), .S(\SUMB[13][34] ) );
  FA1A S2_13_33 ( .A(\ab[13][33] ), .B(\CARRYB[12][33] ), .CI(\SUMB[12][34] ), 
        .CO(\CARRYB[13][33] ), .S(\SUMB[13][33] ) );
  FA1A S2_13_32 ( .A(\ab[13][32] ), .B(\CARRYB[12][32] ), .CI(\SUMB[12][33] ), 
        .CO(\CARRYB[13][32] ), .S(\SUMB[13][32] ) );
  FA1A S2_12_35 ( .A(\ab[12][35] ), .B(\CARRYB[11][35] ), .CI(\SUMB[11][36] ), 
        .CO(\CARRYB[12][35] ), .S(\SUMB[12][35] ) );
  FA1A S2_12_34 ( .A(\ab[12][34] ), .B(\CARRYB[11][34] ), .CI(\SUMB[11][35] ), 
        .CO(\CARRYB[12][34] ), .S(\SUMB[12][34] ) );
  FA1A S2_12_33 ( .A(\ab[12][33] ), .B(\CARRYB[11][33] ), .CI(\SUMB[11][34] ), 
        .CO(\CARRYB[12][33] ), .S(\SUMB[12][33] ) );
  FA1A S2_12_32 ( .A(\ab[12][32] ), .B(\CARRYB[11][32] ), .CI(\SUMB[11][33] ), 
        .CO(\CARRYB[12][32] ), .S(\SUMB[12][32] ) );
  FA1A S2_11_35 ( .A(\ab[11][35] ), .B(\CARRYB[10][35] ), .CI(\SUMB[10][36] ), 
        .CO(\CARRYB[11][35] ), .S(\SUMB[11][35] ) );
  FA1A S2_11_34 ( .A(\ab[11][34] ), .B(\CARRYB[10][34] ), .CI(\SUMB[10][35] ), 
        .CO(\CARRYB[11][34] ), .S(\SUMB[11][34] ) );
  FA1A S2_11_33 ( .A(\ab[11][33] ), .B(\CARRYB[10][33] ), .CI(\SUMB[10][34] ), 
        .CO(\CARRYB[11][33] ), .S(\SUMB[11][33] ) );
  FA1A S2_11_32 ( .A(\ab[11][32] ), .B(\CARRYB[10][32] ), .CI(\SUMB[10][33] ), 
        .CO(\CARRYB[11][32] ), .S(\SUMB[11][32] ) );
  FA1A S2_10_35 ( .A(\ab[10][35] ), .B(\CARRYB[9][35] ), .CI(\SUMB[9][36] ), 
        .CO(\CARRYB[10][35] ), .S(\SUMB[10][35] ) );
  FA1A S2_10_34 ( .A(\ab[10][34] ), .B(\CARRYB[9][34] ), .CI(\SUMB[9][35] ), 
        .CO(\CARRYB[10][34] ), .S(\SUMB[10][34] ) );
  FA1A S2_10_33 ( .A(\ab[10][33] ), .B(\CARRYB[9][33] ), .CI(\SUMB[9][34] ), 
        .CO(\CARRYB[10][33] ), .S(\SUMB[10][33] ) );
  FA1A S2_10_32 ( .A(\ab[10][32] ), .B(\CARRYB[9][32] ), .CI(\SUMB[9][33] ), 
        .CO(\CARRYB[10][32] ), .S(\SUMB[10][32] ) );
  FA1A S2_9_35 ( .A(\ab[9][35] ), .B(\CARRYB[8][35] ), .CI(\SUMB[8][36] ), 
        .CO(\CARRYB[9][35] ), .S(\SUMB[9][35] ) );
  FA1A S2_9_34 ( .A(\ab[9][34] ), .B(\CARRYB[8][34] ), .CI(\SUMB[8][35] ), 
        .CO(\CARRYB[9][34] ), .S(\SUMB[9][34] ) );
  FA1A S2_9_33 ( .A(\ab[9][33] ), .B(\CARRYB[8][33] ), .CI(\SUMB[8][34] ), 
        .CO(\CARRYB[9][33] ), .S(\SUMB[9][33] ) );
  FA1A S2_9_32 ( .A(\ab[9][32] ), .B(\CARRYB[8][32] ), .CI(\SUMB[8][33] ), 
        .CO(\CARRYB[9][32] ), .S(\SUMB[9][32] ) );
  FA1A S2_8_35 ( .A(\ab[8][35] ), .B(\CARRYB[7][35] ), .CI(\SUMB[7][36] ), 
        .CO(\CARRYB[8][35] ), .S(\SUMB[8][35] ) );
  FA1A S2_8_34 ( .A(\ab[8][34] ), .B(\CARRYB[7][34] ), .CI(\SUMB[7][35] ), 
        .CO(\CARRYB[8][34] ), .S(\SUMB[8][34] ) );
  FA1A S2_8_33 ( .A(\ab[8][33] ), .B(\CARRYB[7][33] ), .CI(\SUMB[7][34] ), 
        .CO(\CARRYB[8][33] ), .S(\SUMB[8][33] ) );
  FA1A S2_8_32 ( .A(\ab[8][32] ), .B(\CARRYB[7][32] ), .CI(\SUMB[7][33] ), 
        .CO(\CARRYB[8][32] ), .S(\SUMB[8][32] ) );
  FA1A S2_7_35 ( .A(\ab[7][35] ), .B(\CARRYB[6][35] ), .CI(\SUMB[6][36] ), 
        .CO(\CARRYB[7][35] ), .S(\SUMB[7][35] ) );
  FA1A S2_7_34 ( .A(\ab[7][34] ), .B(\CARRYB[6][34] ), .CI(\SUMB[6][35] ), 
        .CO(\CARRYB[7][34] ), .S(\SUMB[7][34] ) );
  FA1A S2_7_33 ( .A(\ab[7][33] ), .B(\CARRYB[6][33] ), .CI(\SUMB[6][34] ), 
        .CO(\CARRYB[7][33] ), .S(\SUMB[7][33] ) );
  FA1A S2_7_32 ( .A(\ab[7][32] ), .B(\CARRYB[6][32] ), .CI(\SUMB[6][33] ), 
        .CO(\CARRYB[7][32] ), .S(\SUMB[7][32] ) );
  FA1A S2_6_35 ( .A(\ab[6][35] ), .B(\CARRYB[5][35] ), .CI(\SUMB[5][36] ), 
        .CO(\CARRYB[6][35] ), .S(\SUMB[6][35] ) );
  FA1A S2_6_34 ( .A(\ab[6][34] ), .B(\CARRYB[5][34] ), .CI(\SUMB[5][35] ), 
        .CO(\CARRYB[6][34] ), .S(\SUMB[6][34] ) );
  FA1A S2_6_33 ( .A(\ab[6][33] ), .B(\CARRYB[5][33] ), .CI(\SUMB[5][34] ), 
        .CO(\CARRYB[6][33] ), .S(\SUMB[6][33] ) );
  FA1A S2_6_32 ( .A(\ab[6][32] ), .B(\CARRYB[5][32] ), .CI(\SUMB[5][33] ), 
        .CO(\CARRYB[6][32] ), .S(\SUMB[6][32] ) );
  FA1A S2_5_35 ( .A(\ab[5][35] ), .B(\CARRYB[4][35] ), .CI(\SUMB[4][36] ), 
        .CO(\CARRYB[5][35] ), .S(\SUMB[5][35] ) );
  FA1A S2_5_34 ( .A(\ab[5][34] ), .B(\CARRYB[4][34] ), .CI(\SUMB[4][35] ), 
        .CO(\CARRYB[5][34] ), .S(\SUMB[5][34] ) );
  FA1A S2_5_33 ( .A(\ab[5][33] ), .B(\CARRYB[4][33] ), .CI(\SUMB[4][34] ), 
        .CO(\CARRYB[5][33] ), .S(\SUMB[5][33] ) );
  FA1A S2_5_32 ( .A(\ab[5][32] ), .B(\CARRYB[4][32] ), .CI(\SUMB[4][33] ), 
        .CO(\CARRYB[5][32] ), .S(\SUMB[5][32] ) );
  FA1A S2_4_35 ( .A(\ab[4][35] ), .B(\CARRYB[3][35] ), .CI(\SUMB[3][36] ), 
        .CO(\CARRYB[4][35] ), .S(\SUMB[4][35] ) );
  FA1A S2_4_34 ( .A(\ab[4][34] ), .B(\CARRYB[3][34] ), .CI(\SUMB[3][35] ), 
        .CO(\CARRYB[4][34] ), .S(\SUMB[4][34] ) );
  FA1A S2_4_33 ( .A(\ab[4][33] ), .B(\CARRYB[3][33] ), .CI(\SUMB[3][34] ), 
        .CO(\CARRYB[4][33] ), .S(\SUMB[4][33] ) );
  FA1A S2_4_32 ( .A(\ab[4][32] ), .B(\CARRYB[3][32] ), .CI(\SUMB[3][33] ), 
        .CO(\CARRYB[4][32] ), .S(\SUMB[4][32] ) );
  FA1A S2_3_35 ( .A(\ab[3][35] ), .B(\CARRYB[2][35] ), .CI(\SUMB[2][36] ), 
        .CO(\CARRYB[3][35] ), .S(\SUMB[3][35] ) );
  FA1A S2_3_34 ( .A(\ab[3][34] ), .B(\CARRYB[2][34] ), .CI(\SUMB[2][35] ), 
        .CO(\CARRYB[3][34] ), .S(\SUMB[3][34] ) );
  FA1A S2_3_33 ( .A(\ab[3][33] ), .B(\CARRYB[2][33] ), .CI(\SUMB[2][34] ), 
        .CO(\CARRYB[3][33] ), .S(\SUMB[3][33] ) );
  FA1A S2_3_32 ( .A(\ab[3][32] ), .B(\CARRYB[2][32] ), .CI(\SUMB[2][33] ), 
        .CO(\CARRYB[3][32] ), .S(\SUMB[3][32] ) );
  FA1A S2_2_35 ( .A(\ab[2][35] ), .B(\CARRYB[1][35] ), .CI(\SUMB[1][36] ), 
        .CO(\CARRYB[2][35] ), .S(\SUMB[2][35] ) );
  FA1A S2_2_34 ( .A(\ab[2][34] ), .B(\CARRYB[1][34] ), .CI(\SUMB[1][35] ), 
        .CO(\CARRYB[2][34] ), .S(\SUMB[2][34] ) );
  FA1A S2_2_33 ( .A(\ab[2][33] ), .B(\CARRYB[1][33] ), .CI(\SUMB[1][34] ), 
        .CO(\CARRYB[2][33] ), .S(\SUMB[2][33] ) );
  FA1A S2_2_32 ( .A(\ab[2][32] ), .B(\CARRYB[1][32] ), .CI(\SUMB[1][33] ), 
        .CO(\CARRYB[2][32] ), .S(\SUMB[2][32] ) );
  FA1A S4_34 ( .A(\ab[21][34] ), .B(\CARRYB[20][34] ), .CI(\SUMB[20][35] ), 
        .CO(\CARRYB[21][34] ), .S(\SUMB[21][34] ) );
  FA1A S4_35 ( .A(\ab[21][35] ), .B(\CARRYB[20][35] ), .CI(\SUMB[20][36] ), 
        .CO(\CARRYB[21][35] ), .S(\SUMB[21][35] ) );
  FA1A S4_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA1A S2_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\SUMB[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA1A S2_20_31 ( .A(\ab[20][31] ), .B(\CARRYB[19][31] ), .CI(\SUMB[19][32] ), 
        .CO(\CARRYB[20][31] ), .S(\SUMB[20][31] ) );
  FA1A S2_19_31 ( .A(\ab[19][31] ), .B(\CARRYB[18][31] ), .CI(\SUMB[18][32] ), 
        .CO(\CARRYB[19][31] ), .S(\SUMB[19][31] ) );
  FA1A S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA1A S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA1A S2_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\SUMB[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA1A S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA1A S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA1A S2_18_31 ( .A(\ab[18][31] ), .B(\CARRYB[17][31] ), .CI(\SUMB[17][32] ), 
        .CO(\CARRYB[18][31] ), .S(\SUMB[18][31] ) );
  FA1A S2_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\SUMB[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA1A S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA1A S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA1A S2_17_31 ( .A(\ab[17][31] ), .B(\CARRYB[16][31] ), .CI(\SUMB[16][32] ), 
        .CO(\CARRYB[17][31] ), .S(\SUMB[17][31] ) );
  FA1A S2_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\SUMB[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA1A S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA1A S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA1A S2_16_31 ( .A(\ab[16][31] ), .B(\CARRYB[15][31] ), .CI(\SUMB[15][32] ), 
        .CO(\CARRYB[16][31] ), .S(\SUMB[16][31] ) );
  FA1A S2_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\SUMB[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA1A S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA1A S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA1A S2_15_31 ( .A(\ab[15][31] ), .B(\CARRYB[14][31] ), .CI(\SUMB[14][32] ), 
        .CO(\CARRYB[15][31] ), .S(\SUMB[15][31] ) );
  FA1A S2_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\SUMB[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA1A S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA1A S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA1A S2_14_31 ( .A(\ab[14][31] ), .B(\CARRYB[13][31] ), .CI(\SUMB[13][32] ), 
        .CO(\CARRYB[14][31] ), .S(\SUMB[14][31] ) );
  FA1A S2_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\SUMB[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA1A S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA1A S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA1A S2_13_31 ( .A(\ab[13][31] ), .B(\CARRYB[12][31] ), .CI(\SUMB[12][32] ), 
        .CO(\CARRYB[13][31] ), .S(\SUMB[13][31] ) );
  FA1A S2_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\SUMB[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA1A S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA1A S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA1A S2_12_31 ( .A(\ab[12][31] ), .B(\CARRYB[11][31] ), .CI(\SUMB[11][32] ), 
        .CO(\CARRYB[12][31] ), .S(\SUMB[12][31] ) );
  FA1A S2_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\SUMB[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA1A S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA1A S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA1A S2_11_31 ( .A(\ab[11][31] ), .B(\CARRYB[10][31] ), .CI(\SUMB[10][32] ), 
        .CO(\CARRYB[11][31] ), .S(\SUMB[11][31] ) );
  FA1A S2_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\SUMB[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA1A S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1A S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1A S2_10_31 ( .A(\ab[10][31] ), .B(\CARRYB[9][31] ), .CI(\SUMB[9][32] ), 
        .CO(\CARRYB[10][31] ), .S(\SUMB[10][31] ) );
  FA1A S2_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\SUMB[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA1A S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1A S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1A S2_9_31 ( .A(\ab[9][31] ), .B(\CARRYB[8][31] ), .CI(\SUMB[8][32] ), 
        .CO(\CARRYB[9][31] ), .S(\SUMB[9][31] ) );
  FA1A S2_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\SUMB[8][31] ), 
        .CO(\CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA1A S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1A S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1A S2_8_31 ( .A(\ab[8][31] ), .B(\CARRYB[7][31] ), .CI(\SUMB[7][32] ), 
        .CO(\CARRYB[8][31] ), .S(\SUMB[8][31] ) );
  FA1A S2_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\SUMB[7][31] ), 
        .CO(\CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA1A S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1A S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA1A S2_7_31 ( .A(\ab[7][31] ), .B(\CARRYB[6][31] ), .CI(\SUMB[6][32] ), 
        .CO(\CARRYB[7][31] ), .S(\SUMB[7][31] ) );
  FA1A S2_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\SUMB[6][31] ), 
        .CO(\CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA1A S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1A S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA1A S2_6_31 ( .A(\ab[6][31] ), .B(\CARRYB[5][31] ), .CI(\SUMB[5][32] ), 
        .CO(\CARRYB[6][31] ), .S(\SUMB[6][31] ) );
  FA1A S2_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\SUMB[5][31] ), 
        .CO(\CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA1A S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA1A S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1A S2_5_31 ( .A(\ab[5][31] ), .B(\CARRYB[4][31] ), .CI(\SUMB[4][32] ), 
        .CO(\CARRYB[5][31] ), .S(\SUMB[5][31] ) );
  FA1A S2_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\SUMB[4][31] ), 
        .CO(\CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA1A S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA1A S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA1A S2_4_31 ( .A(\ab[4][31] ), .B(\CARRYB[3][31] ), .CI(\SUMB[3][32] ), 
        .CO(\CARRYB[4][31] ), .S(\SUMB[4][31] ) );
  FA1A S2_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\SUMB[3][31] ), 
        .CO(\CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA1A S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\SUMB[3][30] ), 
        .CO(\CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1A S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1A S2_3_31 ( .A(\ab[3][31] ), .B(\CARRYB[2][31] ), .CI(\SUMB[2][32] ), 
        .CO(\CARRYB[3][31] ), .S(\SUMB[3][31] ) );
  FA1A S2_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .CI(\SUMB[2][31] ), 
        .CO(\CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA1A S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1A S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA1A S2_2_31 ( .A(\ab[2][31] ), .B(\CARRYB[1][31] ), .CI(\SUMB[1][32] ), 
        .CO(\CARRYB[2][31] ), .S(\SUMB[2][31] ) );
  FA1A S2_2_30 ( .A(\ab[2][30] ), .B(\CARRYB[1][30] ), .CI(\SUMB[1][31] ), 
        .CO(\CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  FA1A S2_2_29 ( .A(\ab[2][29] ), .B(\CARRYB[1][29] ), .CI(\SUMB[1][30] ), 
        .CO(\CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1A S2_2_28 ( .A(\ab[2][28] ), .B(\CARRYB[1][28] ), .CI(\SUMB[1][29] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FA1A S4_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\SUMB[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA1A S4_31 ( .A(\ab[21][31] ), .B(\CARRYB[20][31] ), .CI(\SUMB[20][32] ), 
        .CO(\CARRYB[21][31] ), .S(\SUMB[21][31] ) );
  FA1A S4_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA1A S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA1A S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA1A S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA1A S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA1A S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA1A S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA1A S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA1A S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA1A S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA1A S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA1A S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA1A S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1A S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1A S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA1A S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA1A S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1A S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1A S2_2_27 ( .A(\ab[2][27] ), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1A S4_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA1A S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA1A S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA1A S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA1A S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA1A S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA1A S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA1A S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA1A S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA1A S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA1A S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1A S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA1A S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1A S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1A S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA1A S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA1A S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1A S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1A S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1A S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1A S4_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA1A S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA1A S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA1A S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA1A S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA1A S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA1A S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA1A S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA1A S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA1A S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA1A S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1A S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1A S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1A S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1A S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA1A S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA1A S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1A S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1A S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA1A S4_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA1A S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA1A S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA1A S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA1A S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA1A S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA1A S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA1A S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA1A S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA1A S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA1A S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1A S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1A S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1A S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1A S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA1A S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1A S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1A S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1A S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA1A S2_2_25 ( .A(\ab[2][25] ), .B(\CARRYB[1][25] ), .CI(\SUMB[1][26] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1A S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), 
        .CO(\CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA1A S4_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA1A S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA1A S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA1A S4_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA1A S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA1A S4_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA1A S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA1A S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA1A S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA1A S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA1A S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA1A S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA1A S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA1A S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA1A S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA1A S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA1A S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA1A S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA1A S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA1A S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA1A S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA1A S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA1A S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA1A S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA1A S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA1A S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA1A S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA1A S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA1A S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA1A S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA1A S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA1A S2_11_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1A S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1A S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1A S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA1A S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1A S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1A S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1A S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1A S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA1A S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1A S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1A S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA1A S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1A S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA1A S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA1A S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA1A S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1A S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1A S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA1A S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1A S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1A S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1A S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1A S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA1A S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1A S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1A S4_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA1A S4_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1A S4_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA1A S4_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA1A S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA1A S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA1A S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA1A S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA1A S4_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA1A S4_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA1A S4_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA1A S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA1A S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA1A S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA1A S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA1A S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA1A S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA1A S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA1A S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA1A S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA1A S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA1A S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA1A S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA1A S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA1A S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA1A S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA1A S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA1A S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA1A S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA1A S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA1A S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA1A S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA1A S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA1A S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA1A S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA1A S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA1A S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA1A S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA1A S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA1A S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA1A S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA1A S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA1A S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA1A S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA1A S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA1A S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA1A S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1A S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA1A S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA1A S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA1A S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA1A S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1A S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA1A S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA1A S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA1A S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1A S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1A S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA1A S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA1A S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA1A S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA1A S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA1A S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1A S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1A S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1A S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA1A S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA1A S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1A S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1A S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1A S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1A S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA1A S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA1A S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA1A S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1A S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1A S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA1A S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), 
        .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA1A S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA1A S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1A S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S4_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA1A S4_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA1A S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA1A S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA1A S4_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA1A S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA1A S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA1A S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA1A S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA1A S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA1A S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA1A S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA1A S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA1A S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA1A S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA1A S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA1A S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA1A S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA1A S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA1A S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA1A S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA1A S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA1A S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA1A S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA1A S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA1A S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA1A S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA1A S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA1A S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA1A S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA1A S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA1A S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA1A S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA1A S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA1A S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1A S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1A S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1A S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1A S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1A S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1A S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1A S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1A S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S4_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA1A S4_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA1A S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA1A S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA1A S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA1A S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S4_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), .CO(
        \CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1A S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1A S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA1A S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA1A S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA1A S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA1A S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1A S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S4_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), .CO(
        \CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1A S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1A S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1A S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S4_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), .CO(
        \CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA1A S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA1A S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1A S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1A S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1A S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA1A S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1A S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1A S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1A S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1A S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S4_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), .CO(
        \CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA1A S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1A S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1A S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1A S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S4_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), .CO(
        \CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1A S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1A S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA1A S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1A S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1A S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA1A S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA1A S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1A S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1A S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1A S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1A S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1A S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA1A S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1A S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA1A S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1A S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1A S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1A S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S4_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), .CO(
        \CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA1A S4_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), .CO(
        \CARRYB[21][0] ), .S(\SUMB[21][0] ) );
  FA1A S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA1A S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA1A S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA1A S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1A S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA1A S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1A S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1A S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1A S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1A S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1A S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1A S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1A S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1A S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1A S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S4_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), .CO(
        \CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1A S4_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), .CO(
        \CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1A S4_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), .CO(
        \CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1A S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1A S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA1A S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1A S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1A S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1A S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  IVP U2 ( .A(n40), .Z(n38) );
  IVP U3 ( .A(n40), .Z(n37) );
  IVP U4 ( .A(n40), .Z(n39) );
  IVP U5 ( .A(n40), .Z(n36) );
  IVP U6 ( .A(n112), .Z(n40) );
  IVP U7 ( .A(A[0]), .Z(n112) );
  IVP U8 ( .A(n45), .Z(n41) );
  IVP U9 ( .A(n45), .Z(n42) );
  IVP U10 ( .A(n45), .Z(n43) );
  IVP U11 ( .A(n50), .Z(n47) );
  IVP U12 ( .A(n50), .Z(n48) );
  IVP U13 ( .A(n50), .Z(n49) );
  IVP U14 ( .A(n50), .Z(n46) );
  IVP U15 ( .A(n45), .Z(n44) );
  IVP U16 ( .A(n55), .Z(n52) );
  IVP U17 ( .A(n55), .Z(n53) );
  IVP U18 ( .A(n55), .Z(n51) );
  IVP U19 ( .A(n55), .Z(n54) );
  IVP U20 ( .A(n60), .Z(n57) );
  IVP U21 ( .A(n60), .Z(n56) );
  IVP U22 ( .A(n60), .Z(n58) );
  IVP U23 ( .A(n60), .Z(n59) );
  IVP U24 ( .A(n65), .Z(n62) );
  IVP U25 ( .A(n65), .Z(n61) );
  IVP U26 ( .A(n65), .Z(n64) );
  IVP U27 ( .A(n65), .Z(n63) );
  IVP U28 ( .A(n70), .Z(n67) );
  IVP U29 ( .A(n70), .Z(n66) );
  IVP U30 ( .A(n70), .Z(n69) );
  IVP U31 ( .A(n70), .Z(n68) );
  IVP U32 ( .A(n75), .Z(n72) );
  IVP U33 ( .A(n75), .Z(n71) );
  IVP U34 ( .A(n75), .Z(n73) );
  IVP U35 ( .A(n75), .Z(n74) );
  IVP U36 ( .A(n80), .Z(n76) );
  IVP U37 ( .A(n80), .Z(n77) );
  IVP U38 ( .A(n80), .Z(n78) );
  IVP U39 ( .A(n80), .Z(n79) );
  IVP U40 ( .A(n85), .Z(n82) );
  IVP U41 ( .A(n85), .Z(n83) );
  IVP U42 ( .A(n85), .Z(n81) );
  IVP U43 ( .A(n85), .Z(n84) );
  IVP U44 ( .A(n90), .Z(n87) );
  IVP U45 ( .A(n90), .Z(n88) );
  IVP U46 ( .A(n90), .Z(n86) );
  IVP U47 ( .A(n90), .Z(n89) );
  IVP U48 ( .A(n95), .Z(n92) );
  IVP U49 ( .A(n95), .Z(n93) );
  IVP U50 ( .A(n95), .Z(n91) );
  IVP U51 ( .A(n95), .Z(n94) );
  IVP U52 ( .A(n100), .Z(n97) );
  IVP U53 ( .A(n100), .Z(n98) );
  IVP U54 ( .A(n100), .Z(n96) );
  IVP U55 ( .A(n100), .Z(n99) );
  IVP U56 ( .A(n113), .Z(n45) );
  IVP U57 ( .A(A[1]), .Z(n113) );
  IVP U58 ( .A(n114), .Z(n50) );
  IVP U59 ( .A(A[2]), .Z(n114) );
  IVP U60 ( .A(n115), .Z(n55) );
  IVP U61 ( .A(A[3]), .Z(n115) );
  IVP U62 ( .A(n116), .Z(n60) );
  IVP U63 ( .A(A[4]), .Z(n116) );
  IVP U64 ( .A(n117), .Z(n65) );
  IVP U65 ( .A(A[5]), .Z(n117) );
  IVP U66 ( .A(n118), .Z(n70) );
  IVP U67 ( .A(A[6]), .Z(n118) );
  IVP U68 ( .A(n119), .Z(n75) );
  IVP U69 ( .A(A[7]), .Z(n119) );
  IVP U70 ( .A(n120), .Z(n80) );
  IVP U71 ( .A(A[8]), .Z(n120) );
  IVP U72 ( .A(n121), .Z(n85) );
  IVP U73 ( .A(A[9]), .Z(n121) );
  IVP U74 ( .A(n122), .Z(n90) );
  IVP U75 ( .A(A[10]), .Z(n122) );
  IVP U76 ( .A(n123), .Z(n95) );
  IVP U77 ( .A(A[11]), .Z(n123) );
  IVP U78 ( .A(n124), .Z(n100) );
  IVP U79 ( .A(A[12]), .Z(n124) );
  IVP U80 ( .A(n35), .Z(n32) );
  IVP U81 ( .A(n35), .Z(n33) );
  IVP U82 ( .A(n35), .Z(n31) );
  IVP U83 ( .A(n35), .Z(n34) );
  IVP U84 ( .A(n7), .Z(n4) );
  IVP U85 ( .A(n7), .Z(n3) );
  IVP U86 ( .A(n30), .Z(n27) );
  IVP U87 ( .A(n7), .Z(n5) );
  IVP U88 ( .A(n30), .Z(n26) );
  IVP U89 ( .A(n7), .Z(n6) );
  IVP U90 ( .A(n30), .Z(n28) );
  IVP U91 ( .A(n30), .Z(n29) );
  IVP U92 ( .A(A[16]), .Z(n23) );
  IVP U93 ( .A(A[16]), .Z(n24) );
  IVP U94 ( .A(A[16]), .Z(n25) );
  IVP U95 ( .A(A[17]), .Z(n22) );
  IVP U96 ( .A(A[18]), .Z(n20) );
  IVP U97 ( .A(A[18]), .Z(n21) );
  IVP U98 ( .A(A[19]), .Z(n17) );
  IVP U99 ( .A(A[19]), .Z(n16) );
  IVP U100 ( .A(A[19]), .Z(n18) );
  IVP U101 ( .A(A[19]), .Z(n19) );
  IVP U102 ( .A(A[20]), .Z(n13) );
  IVP U103 ( .A(A[20]), .Z(n12) );
  IVP U104 ( .A(A[20]), .Z(n14) );
  IVP U105 ( .A(A[20]), .Z(n15) );
  IVP U106 ( .A(A[21]), .Z(n9) );
  IVP U107 ( .A(A[21]), .Z(n10) );
  IVP U108 ( .A(A[21]), .Z(n8) );
  IVP U109 ( .A(A[21]), .Z(n11) );
  IVP U110 ( .A(n111), .Z(n35) );
  IVP U111 ( .A(A[13]), .Z(n111) );
  IVP U112 ( .A(n109), .Z(n7) );
  IVP U113 ( .A(A[14]), .Z(n109) );
  IVP U114 ( .A(n110), .Z(n30) );
  IVP U115 ( .A(A[15]), .Z(n110) );
  EO U116 ( .A(\CARRYB[21][4] ), .B(\SUMB[21][5] ), .Z(\A1[24] ) );
  EO U117 ( .A(\CARRYB[21][9] ), .B(\SUMB[21][10] ), .Z(\A1[29] ) );
  EO U118 ( .A(\CARRYB[21][1] ), .B(\SUMB[21][2] ), .Z(\A1[21] ) );
  EO U119 ( .A(\CARRYB[21][2] ), .B(\SUMB[21][3] ), .Z(\A1[22] ) );
  EO U120 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  EO U121 ( .A(\CARRYB[21][3] ), .B(\SUMB[21][4] ), .Z(\A1[23] ) );
  EO U122 ( .A(\CARRYB[21][5] ), .B(\SUMB[21][6] ), .Z(\A1[25] ) );
  EO U123 ( .A(\CARRYB[21][6] ), .B(\SUMB[21][7] ), .Z(\A1[26] ) );
  EO U124 ( .A(\CARRYB[21][7] ), .B(\SUMB[21][8] ), .Z(\A1[27] ) );
  EO U125 ( .A(\CARRYB[21][8] ), .B(\SUMB[21][9] ), .Z(\A1[28] ) );
  EO U126 ( .A(\CARRYB[21][17] ), .B(\SUMB[21][18] ), .Z(\A1[37] ) );
  EO U127 ( .A(\CARRYB[21][13] ), .B(\SUMB[21][14] ), .Z(\A1[33] ) );
  EO U128 ( .A(\CARRYB[21][12] ), .B(\SUMB[21][13] ), .Z(\A1[32] ) );
  EO U129 ( .A(\CARRYB[21][16] ), .B(\SUMB[21][17] ), .Z(\A1[36] ) );
  EO U130 ( .A(\CARRYB[21][18] ), .B(\SUMB[21][19] ), .Z(\A1[38] ) );
  EO U131 ( .A(\CARRYB[21][21] ), .B(\SUMB[21][22] ), .Z(\A1[41] ) );
  EO U132 ( .A(\CARRYB[21][19] ), .B(\SUMB[21][20] ), .Z(\A1[39] ) );
  EO U133 ( .A(\CARRYB[21][20] ), .B(\SUMB[21][21] ), .Z(\A1[40] ) );
  EO U134 ( .A(\CARRYB[21][15] ), .B(\SUMB[21][16] ), .Z(\A1[35] ) );
  EO U135 ( .A(\CARRYB[21][14] ), .B(\SUMB[21][15] ), .Z(\A1[34] ) );
  EO U136 ( .A(\CARRYB[21][22] ), .B(\SUMB[21][23] ), .Z(\A1[42] ) );
  EO U137 ( .A(\CARRYB[21][10] ), .B(\SUMB[21][11] ), .Z(\A1[30] ) );
  EO U138 ( .A(\CARRYB[21][23] ), .B(\SUMB[21][24] ), .Z(\A1[43] ) );
  EO U139 ( .A(\CARRYB[21][11] ), .B(\SUMB[21][12] ), .Z(\A1[31] ) );
  EO U140 ( .A(\CARRYB[21][24] ), .B(\SUMB[21][25] ), .Z(\A1[44] ) );
  EO U141 ( .A(\CARRYB[21][25] ), .B(\SUMB[21][26] ), .Z(\A1[45] ) );
  EO U142 ( .A(\CARRYB[21][26] ), .B(\SUMB[21][27] ), .Z(\A1[46] ) );
  EO U143 ( .A(\CARRYB[21][29] ), .B(\SUMB[21][30] ), .Z(\A1[49] ) );
  EO U144 ( .A(\CARRYB[21][27] ), .B(\SUMB[21][28] ), .Z(\A1[47] ) );
  EO U145 ( .A(\CARRYB[21][30] ), .B(\SUMB[21][31] ), .Z(\A1[50] ) );
  EO U146 ( .A(\CARRYB[21][28] ), .B(\SUMB[21][29] ), .Z(\A1[48] ) );
  EO U147 ( .A(\CARRYB[21][33] ), .B(\SUMB[21][34] ), .Z(\A1[53] ) );
  EO U148 ( .A(\CARRYB[21][34] ), .B(\SUMB[21][35] ), .Z(\A1[54] ) );
  EO U149 ( .A(\CARRYB[21][32] ), .B(\SUMB[21][33] ), .Z(\A1[52] ) );
  EO U150 ( .A(\CARRYB[21][37] ), .B(\SUMB[21][38] ), .Z(\A1[57] ) );
  EO U151 ( .A(\CARRYB[21][31] ), .B(\SUMB[21][32] ), .Z(\A1[51] ) );
  EO U152 ( .A(\CARRYB[21][35] ), .B(\SUMB[21][36] ), .Z(\A1[55] ) );
  EO U153 ( .A(\CARRYB[21][38] ), .B(\SUMB[21][39] ), .Z(\A1[58] ) );
  EO U154 ( .A(\CARRYB[21][36] ), .B(\SUMB[21][37] ), .Z(\A1[56] ) );
  EO U155 ( .A(\CARRYB[21][39] ), .B(\SUMB[21][40] ), .Z(\A1[59] ) );
  EO U156 ( .A(\CARRYB[21][40] ), .B(\SUMB[21][41] ), .Z(\A1[60] ) );
  EO U157 ( .A(\CARRYB[21][41] ), .B(\SUMB[21][42] ), .Z(\A1[61] ) );
  EO U158 ( .A(\CARRYB[21][42] ), .B(\SUMB[21][43] ), .Z(\A1[62] ) );
  EO U159 ( .A(\CARRYB[21][43] ), .B(\SUMB[21][44] ), .Z(\A1[63] ) );
  EO U160 ( .A(\CARRYB[21][44] ), .B(\SUMB[21][45] ), .Z(\A1[64] ) );
  EO U161 ( .A(\CARRYB[21][45] ), .B(\SUMB[21][46] ), .Z(\A1[65] ) );
  EO U162 ( .A(\CARRYB[21][0] ), .B(\SUMB[21][1] ), .Z(\A1[20] ) );
  EO U163 ( .A(\CARRYB[21][46] ), .B(\ab[21][47] ), .Z(\A1[66] ) );
  EO U164 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U165 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U166 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U167 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U168 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U169 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U170 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U171 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U172 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U173 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U174 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U175 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U176 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U177 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U178 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Z(\SUMB[1][18] ) );
  EO U179 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Z(\SUMB[1][19] ) );
  EO U180 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Z(\SUMB[1][16] ) );
  EO U181 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Z(\SUMB[1][17] ) );
  EO U182 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Z(\SUMB[1][20] ) );
  EO U183 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Z(\SUMB[1][22] ) );
  EO U184 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Z(\SUMB[1][23] ) );
  EO U185 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Z(\SUMB[1][21] ) );
  EO U186 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Z(\SUMB[1][24] ) );
  EO U187 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Z(\SUMB[1][25] ) );
  EO U188 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Z(\SUMB[1][26] ) );
  EO U189 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Z(\SUMB[1][27] ) );
  EO U190 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Z(\SUMB[1][28] ) );
  EO U191 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Z(\SUMB[1][29] ) );
  EO U192 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Z(\SUMB[1][30] ) );
  EO U193 ( .A(\ab[0][32] ), .B(\ab[1][31] ), .Z(\SUMB[1][31] ) );
  EO U194 ( .A(\ab[0][33] ), .B(\ab[1][32] ), .Z(\SUMB[1][32] ) );
  EO U195 ( .A(\ab[0][34] ), .B(\ab[1][33] ), .Z(\SUMB[1][33] ) );
  EO U196 ( .A(\ab[0][35] ), .B(\ab[1][34] ), .Z(\SUMB[1][34] ) );
  EO U197 ( .A(\ab[0][36] ), .B(\ab[1][35] ), .Z(\SUMB[1][35] ) );
  EO U198 ( .A(\ab[0][37] ), .B(\ab[1][36] ), .Z(\SUMB[1][36] ) );
  EO U199 ( .A(\ab[0][38] ), .B(\ab[1][37] ), .Z(\SUMB[1][37] ) );
  EO U200 ( .A(\ab[0][39] ), .B(\ab[1][38] ), .Z(\SUMB[1][38] ) );
  EO U201 ( .A(\ab[0][40] ), .B(\ab[1][39] ), .Z(\SUMB[1][39] ) );
  EO U202 ( .A(\ab[0][41] ), .B(\ab[1][40] ), .Z(\SUMB[1][40] ) );
  EO U203 ( .A(\ab[0][42] ), .B(\ab[1][41] ), .Z(\SUMB[1][41] ) );
  EO U204 ( .A(\ab[0][43] ), .B(\ab[1][42] ), .Z(\SUMB[1][42] ) );
  EO U205 ( .A(\ab[0][44] ), .B(\ab[1][43] ), .Z(\SUMB[1][43] ) );
  EO U206 ( .A(\ab[0][45] ), .B(\ab[1][44] ), .Z(\SUMB[1][44] ) );
  EO U207 ( .A(\ab[0][46] ), .B(\ab[1][45] ), .Z(\SUMB[1][45] ) );
  EO U208 ( .A(\ab[0][47] ), .B(\ab[1][46] ), .Z(\SUMB[1][46] ) );
  IVP U209 ( .A(B[2]), .Z(n162) );
  IVP U210 ( .A(B[3]), .Z(n161) );
  IVP U211 ( .A(B[4]), .Z(n160) );
  IVP U212 ( .A(B[1]), .Z(n163) );
  IVP U213 ( .A(B[5]), .Z(n159) );
  IVP U214 ( .A(B[0]), .Z(n164) );
  IVP U215 ( .A(B[6]), .Z(n158) );
  IVP U216 ( .A(B[7]), .Z(n157) );
  IVP U217 ( .A(B[8]), .Z(n156) );
  IVP U218 ( .A(B[9]), .Z(n155) );
  IVP U219 ( .A(B[10]), .Z(n154) );
  IVP U220 ( .A(B[11]), .Z(n153) );
  IVP U221 ( .A(B[12]), .Z(n152) );
  IVP U222 ( .A(B[13]), .Z(n151) );
  IVP U223 ( .A(B[14]), .Z(n150) );
  IVP U224 ( .A(B[15]), .Z(n149) );
  IVP U225 ( .A(B[16]), .Z(n148) );
  IVP U226 ( .A(B[17]), .Z(n147) );
  IVP U227 ( .A(B[18]), .Z(n146) );
  IVP U228 ( .A(B[19]), .Z(n145) );
  IVP U229 ( .A(B[20]), .Z(n144) );
  IVP U230 ( .A(B[21]), .Z(n143) );
  IVP U231 ( .A(B[22]), .Z(n142) );
  IVP U232 ( .A(B[23]), .Z(n141) );
  IVP U233 ( .A(B[24]), .Z(n140) );
  IVP U234 ( .A(B[25]), .Z(n139) );
  IVP U235 ( .A(B[26]), .Z(n138) );
  IVP U236 ( .A(B[27]), .Z(n137) );
  IVP U237 ( .A(B[28]), .Z(n136) );
  IVP U238 ( .A(B[29]), .Z(n135) );
  IVP U239 ( .A(B[30]), .Z(n134) );
  IVP U240 ( .A(B[31]), .Z(n133) );
  IVP U241 ( .A(B[32]), .Z(n132) );
  IVP U242 ( .A(B[33]), .Z(n131) );
  IVP U243 ( .A(B[34]), .Z(n130) );
  IVP U244 ( .A(B[35]), .Z(n129) );
  IVP U245 ( .A(B[36]), .Z(n128) );
  IVP U246 ( .A(B[37]), .Z(n127) );
  IVP U247 ( .A(B[38]), .Z(n126) );
  IVP U248 ( .A(B[39]), .Z(n125) );
  IVP U249 ( .A(B[40]), .Z(n101) );
  IVP U250 ( .A(B[41]), .Z(n102) );
  IVP U251 ( .A(B[42]), .Z(n103) );
  IVP U252 ( .A(B[43]), .Z(n104) );
  IVP U253 ( .A(B[44]), .Z(n105) );
  IVP U254 ( .A(B[45]), .Z(n106) );
  IVP U255 ( .A(B[47]), .Z(n108) );
  IVP U256 ( .A(B[46]), .Z(n107) );
  AN2P U257 ( .A(\CARRYB[21][0] ), .B(\SUMB[21][1] ), .Z(\A2[21] ) );
  AN2P U258 ( .A(\CARRYB[21][1] ), .B(\SUMB[21][2] ), .Z(\A2[22] ) );
  AN2P U259 ( .A(\CARRYB[21][2] ), .B(\SUMB[21][3] ), .Z(\A2[23] ) );
  AN2P U260 ( .A(\CARRYB[21][3] ), .B(\SUMB[21][4] ), .Z(\A2[24] ) );
  AN2P U261 ( .A(\CARRYB[21][4] ), .B(\SUMB[21][5] ), .Z(\A2[25] ) );
  AN2P U262 ( .A(\CARRYB[21][5] ), .B(\SUMB[21][6] ), .Z(\A2[26] ) );
  AN2P U263 ( .A(\CARRYB[21][6] ), .B(\SUMB[21][7] ), .Z(\A2[27] ) );
  AN2P U264 ( .A(\CARRYB[21][7] ), .B(\SUMB[21][8] ), .Z(\A2[28] ) );
  AN2P U265 ( .A(\CARRYB[21][8] ), .B(\SUMB[21][9] ), .Z(\A2[29] ) );
  AN2P U266 ( .A(\CARRYB[21][9] ), .B(\SUMB[21][10] ), .Z(\A2[30] ) );
  AN2P U267 ( .A(\CARRYB[21][10] ), .B(\SUMB[21][11] ), .Z(\A2[31] ) );
  AN2P U268 ( .A(\CARRYB[21][11] ), .B(\SUMB[21][12] ), .Z(\A2[32] ) );
  AN2P U269 ( .A(\CARRYB[21][12] ), .B(\SUMB[21][13] ), .Z(\A2[33] ) );
  AN2P U270 ( .A(\CARRYB[21][13] ), .B(\SUMB[21][14] ), .Z(\A2[34] ) );
  AN2P U271 ( .A(\CARRYB[21][14] ), .B(\SUMB[21][15] ), .Z(\A2[35] ) );
  AN2P U272 ( .A(\CARRYB[21][15] ), .B(\SUMB[21][16] ), .Z(\A2[36] ) );
  AN2P U273 ( .A(\CARRYB[21][16] ), .B(\SUMB[21][17] ), .Z(\A2[37] ) );
  AN2P U274 ( .A(\CARRYB[21][17] ), .B(\SUMB[21][18] ), .Z(\A2[38] ) );
  AN2P U275 ( .A(\CARRYB[21][18] ), .B(\SUMB[21][19] ), .Z(\A2[39] ) );
  AN2P U276 ( .A(\CARRYB[21][19] ), .B(\SUMB[21][20] ), .Z(\A2[40] ) );
  AN2P U277 ( .A(\CARRYB[21][20] ), .B(\SUMB[21][21] ), .Z(\A2[41] ) );
  AN2P U278 ( .A(\CARRYB[21][21] ), .B(\SUMB[21][22] ), .Z(\A2[42] ) );
  AN2P U279 ( .A(\CARRYB[21][22] ), .B(\SUMB[21][23] ), .Z(\A2[43] ) );
  AN2P U280 ( .A(\CARRYB[21][23] ), .B(\SUMB[21][24] ), .Z(\A2[44] ) );
  AN2P U281 ( .A(\CARRYB[21][24] ), .B(\SUMB[21][25] ), .Z(\A2[45] ) );
  AN2P U282 ( .A(\CARRYB[21][26] ), .B(\SUMB[21][27] ), .Z(\A2[47] ) );
  AN2P U283 ( .A(\CARRYB[21][27] ), .B(\SUMB[21][28] ), .Z(\A2[48] ) );
  AN2P U284 ( .A(\CARRYB[21][28] ), .B(\SUMB[21][29] ), .Z(\A2[49] ) );
  AN2P U285 ( .A(\CARRYB[21][29] ), .B(\SUMB[21][30] ), .Z(\A2[50] ) );
  AN2P U286 ( .A(\CARRYB[21][30] ), .B(\SUMB[21][31] ), .Z(\A2[51] ) );
  AN2P U287 ( .A(\CARRYB[21][31] ), .B(\SUMB[21][32] ), .Z(\A2[52] ) );
  AN2P U288 ( .A(\CARRYB[21][32] ), .B(\SUMB[21][33] ), .Z(\A2[53] ) );
  AN2P U289 ( .A(\CARRYB[21][33] ), .B(\SUMB[21][34] ), .Z(\A2[54] ) );
  AN2P U290 ( .A(\CARRYB[21][34] ), .B(\SUMB[21][35] ), .Z(\A2[55] ) );
  AN2P U291 ( .A(\CARRYB[21][35] ), .B(\SUMB[21][36] ), .Z(\A2[56] ) );
  AN2P U292 ( .A(\CARRYB[21][36] ), .B(\SUMB[21][37] ), .Z(\A2[57] ) );
  AN2P U293 ( .A(\CARRYB[21][37] ), .B(\SUMB[21][38] ), .Z(\A2[58] ) );
  AN2P U294 ( .A(\CARRYB[21][38] ), .B(\SUMB[21][39] ), .Z(\A2[59] ) );
  AN2P U295 ( .A(\CARRYB[21][39] ), .B(\SUMB[21][40] ), .Z(\A2[60] ) );
  AN2P U296 ( .A(\CARRYB[21][40] ), .B(\SUMB[21][41] ), .Z(\A2[61] ) );
  AN2P U297 ( .A(\CARRYB[21][41] ), .B(\SUMB[21][42] ), .Z(\A2[62] ) );
  AN2P U298 ( .A(\CARRYB[21][42] ), .B(\SUMB[21][43] ), .Z(\A2[63] ) );
  AN2P U299 ( .A(\CARRYB[21][43] ), .B(\SUMB[21][44] ), .Z(\A2[64] ) );
  AN2P U300 ( .A(\CARRYB[21][44] ), .B(\SUMB[21][45] ), .Z(\A2[65] ) );
  AN2P U301 ( .A(\CARRYB[21][45] ), .B(\SUMB[21][46] ), .Z(\A2[66] ) );
  AN2P U302 ( .A(\CARRYB[21][46] ), .B(\ab[21][47] ), .Z(\A2[67] ) );
  AN2P U303 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U304 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U305 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U306 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U307 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U308 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U309 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U310 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U311 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U312 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U313 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U314 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U315 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U316 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U317 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U318 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\CARRYB[1][16] ) );
  AN2P U319 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\CARRYB[1][17] ) );
  AN2P U320 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\CARRYB[1][18] ) );
  AN2P U321 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\CARRYB[1][19] ) );
  AN2P U322 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\CARRYB[1][20] ) );
  AN2P U323 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\CARRYB[1][21] ) );
  AN2P U324 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(\CARRYB[1][22] ) );
  AN2P U325 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(\CARRYB[1][23] ) );
  AN2P U326 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(\CARRYB[1][24] ) );
  AN2P U327 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(\CARRYB[1][25] ) );
  AN2P U328 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\CARRYB[1][26] ) );
  AN2P U329 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(\CARRYB[1][27] ) );
  AN2P U330 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(\CARRYB[1][28] ) );
  AN2P U331 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(\CARRYB[1][29] ) );
  AN2P U332 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(\CARRYB[1][30] ) );
  AN2P U333 ( .A(\ab[1][31] ), .B(\ab[0][32] ), .Z(\CARRYB[1][31] ) );
  AN2P U334 ( .A(\ab[1][32] ), .B(\ab[0][33] ), .Z(\CARRYB[1][32] ) );
  AN2P U335 ( .A(\ab[1][33] ), .B(\ab[0][34] ), .Z(\CARRYB[1][33] ) );
  AN2P U336 ( .A(\ab[1][34] ), .B(\ab[0][35] ), .Z(\CARRYB[1][34] ) );
  AN2P U337 ( .A(\ab[1][35] ), .B(\ab[0][36] ), .Z(\CARRYB[1][35] ) );
  AN2P U338 ( .A(\ab[1][36] ), .B(\ab[0][37] ), .Z(\CARRYB[1][36] ) );
  AN2P U339 ( .A(\ab[1][37] ), .B(\ab[0][38] ), .Z(\CARRYB[1][37] ) );
  AN2P U340 ( .A(\ab[1][38] ), .B(\ab[0][39] ), .Z(\CARRYB[1][38] ) );
  AN2P U341 ( .A(\ab[1][39] ), .B(\ab[0][40] ), .Z(\CARRYB[1][39] ) );
  AN2P U342 ( .A(\ab[1][40] ), .B(\ab[0][41] ), .Z(\CARRYB[1][40] ) );
  AN2P U343 ( .A(\ab[1][41] ), .B(\ab[0][42] ), .Z(\CARRYB[1][41] ) );
  AN2P U344 ( .A(\ab[1][42] ), .B(\ab[0][43] ), .Z(\CARRYB[1][42] ) );
  AN2P U345 ( .A(\ab[1][43] ), .B(\ab[0][44] ), .Z(\CARRYB[1][43] ) );
  AN2P U346 ( .A(\ab[1][44] ), .B(\ab[0][45] ), .Z(\CARRYB[1][44] ) );
  AN2P U347 ( .A(\ab[1][45] ), .B(\ab[0][46] ), .Z(\CARRYB[1][45] ) );
  AN2P U348 ( .A(\ab[1][46] ), .B(\ab[0][47] ), .Z(\CARRYB[1][46] ) );
  AN2P U349 ( .A(\CARRYB[21][25] ), .B(\SUMB[21][26] ), .Z(\A2[46] ) );
  NR2 U351 ( .A(n84), .B(n155), .Z(\ab[9][9] ) );
  NR2 U352 ( .A(n84), .B(n156), .Z(\ab[9][8] ) );
  NR2 U353 ( .A(n84), .B(n157), .Z(\ab[9][7] ) );
  NR2 U354 ( .A(n84), .B(n158), .Z(\ab[9][6] ) );
  NR2 U355 ( .A(n84), .B(n159), .Z(\ab[9][5] ) );
  NR2 U356 ( .A(n84), .B(n160), .Z(\ab[9][4] ) );
  NR2 U357 ( .A(n84), .B(n108), .Z(\ab[9][47] ) );
  NR2 U358 ( .A(n84), .B(n107), .Z(\ab[9][46] ) );
  NR2 U359 ( .A(n84), .B(n106), .Z(\ab[9][45] ) );
  NR2 U360 ( .A(n84), .B(n105), .Z(\ab[9][44] ) );
  NR2 U361 ( .A(n84), .B(n104), .Z(\ab[9][43] ) );
  NR2 U362 ( .A(n84), .B(n103), .Z(\ab[9][42] ) );
  NR2 U363 ( .A(n83), .B(n102), .Z(\ab[9][41] ) );
  NR2 U364 ( .A(n83), .B(n101), .Z(\ab[9][40] ) );
  NR2 U365 ( .A(n83), .B(n161), .Z(\ab[9][3] ) );
  NR2 U366 ( .A(n83), .B(n125), .Z(\ab[9][39] ) );
  NR2 U367 ( .A(n83), .B(n126), .Z(\ab[9][38] ) );
  NR2 U368 ( .A(n83), .B(n127), .Z(\ab[9][37] ) );
  NR2 U369 ( .A(n83), .B(n128), .Z(\ab[9][36] ) );
  NR2 U370 ( .A(n83), .B(n129), .Z(\ab[9][35] ) );
  NR2 U371 ( .A(n83), .B(n130), .Z(\ab[9][34] ) );
  NR2 U372 ( .A(n83), .B(n131), .Z(\ab[9][33] ) );
  NR2 U373 ( .A(n83), .B(n132), .Z(\ab[9][32] ) );
  NR2 U374 ( .A(n83), .B(n133), .Z(\ab[9][31] ) );
  NR2 U375 ( .A(n82), .B(n134), .Z(\ab[9][30] ) );
  NR2 U376 ( .A(n82), .B(n162), .Z(\ab[9][2] ) );
  NR2 U377 ( .A(n82), .B(n135), .Z(\ab[9][29] ) );
  NR2 U378 ( .A(n82), .B(n136), .Z(\ab[9][28] ) );
  NR2 U379 ( .A(n82), .B(n137), .Z(\ab[9][27] ) );
  NR2 U380 ( .A(n82), .B(n138), .Z(\ab[9][26] ) );
  NR2 U381 ( .A(n82), .B(n139), .Z(\ab[9][25] ) );
  NR2 U382 ( .A(n82), .B(n140), .Z(\ab[9][24] ) );
  NR2 U383 ( .A(n82), .B(n141), .Z(\ab[9][23] ) );
  NR2 U384 ( .A(n82), .B(n142), .Z(\ab[9][22] ) );
  NR2 U385 ( .A(n82), .B(n143), .Z(\ab[9][21] ) );
  NR2 U386 ( .A(n82), .B(n144), .Z(\ab[9][20] ) );
  NR2 U387 ( .A(n81), .B(n163), .Z(\ab[9][1] ) );
  NR2 U388 ( .A(n81), .B(n145), .Z(\ab[9][19] ) );
  NR2 U389 ( .A(n81), .B(n146), .Z(\ab[9][18] ) );
  NR2 U390 ( .A(n81), .B(n147), .Z(\ab[9][17] ) );
  NR2 U391 ( .A(n81), .B(n148), .Z(\ab[9][16] ) );
  NR2 U392 ( .A(n81), .B(n149), .Z(\ab[9][15] ) );
  NR2 U393 ( .A(n81), .B(n150), .Z(\ab[9][14] ) );
  NR2 U394 ( .A(n81), .B(n151), .Z(\ab[9][13] ) );
  NR2 U395 ( .A(n81), .B(n152), .Z(\ab[9][12] ) );
  NR2 U396 ( .A(n81), .B(n153), .Z(\ab[9][11] ) );
  NR2 U397 ( .A(n81), .B(n154), .Z(\ab[9][10] ) );
  NR2 U398 ( .A(n81), .B(n164), .Z(\ab[9][0] ) );
  NR2 U399 ( .A(n155), .B(n79), .Z(\ab[8][9] ) );
  NR2 U400 ( .A(n156), .B(n79), .Z(\ab[8][8] ) );
  NR2 U401 ( .A(n157), .B(n79), .Z(\ab[8][7] ) );
  NR2 U402 ( .A(n158), .B(n79), .Z(\ab[8][6] ) );
  NR2 U403 ( .A(n159), .B(n79), .Z(\ab[8][5] ) );
  NR2 U404 ( .A(n160), .B(n79), .Z(\ab[8][4] ) );
  NR2 U405 ( .A(n108), .B(n79), .Z(\ab[8][47] ) );
  NR2 U406 ( .A(n107), .B(n79), .Z(\ab[8][46] ) );
  NR2 U407 ( .A(n106), .B(n79), .Z(\ab[8][45] ) );
  NR2 U408 ( .A(n105), .B(n79), .Z(\ab[8][44] ) );
  NR2 U409 ( .A(n104), .B(n79), .Z(\ab[8][43] ) );
  NR2 U410 ( .A(n103), .B(n79), .Z(\ab[8][42] ) );
  NR2 U411 ( .A(n102), .B(n78), .Z(\ab[8][41] ) );
  NR2 U412 ( .A(n101), .B(n78), .Z(\ab[8][40] ) );
  NR2 U413 ( .A(n161), .B(n78), .Z(\ab[8][3] ) );
  NR2 U414 ( .A(n125), .B(n78), .Z(\ab[8][39] ) );
  NR2 U415 ( .A(n126), .B(n78), .Z(\ab[8][38] ) );
  NR2 U416 ( .A(n127), .B(n78), .Z(\ab[8][37] ) );
  NR2 U417 ( .A(n128), .B(n78), .Z(\ab[8][36] ) );
  NR2 U418 ( .A(n129), .B(n78), .Z(\ab[8][35] ) );
  NR2 U419 ( .A(n130), .B(n78), .Z(\ab[8][34] ) );
  NR2 U420 ( .A(n131), .B(n78), .Z(\ab[8][33] ) );
  NR2 U421 ( .A(n132), .B(n78), .Z(\ab[8][32] ) );
  NR2 U422 ( .A(n133), .B(n78), .Z(\ab[8][31] ) );
  NR2 U423 ( .A(n134), .B(n77), .Z(\ab[8][30] ) );
  NR2 U424 ( .A(n162), .B(n77), .Z(\ab[8][2] ) );
  NR2 U425 ( .A(n135), .B(n77), .Z(\ab[8][29] ) );
  NR2 U426 ( .A(n136), .B(n77), .Z(\ab[8][28] ) );
  NR2 U427 ( .A(n137), .B(n77), .Z(\ab[8][27] ) );
  NR2 U428 ( .A(n138), .B(n77), .Z(\ab[8][26] ) );
  NR2 U429 ( .A(n139), .B(n77), .Z(\ab[8][25] ) );
  NR2 U430 ( .A(n140), .B(n77), .Z(\ab[8][24] ) );
  NR2 U431 ( .A(n141), .B(n77), .Z(\ab[8][23] ) );
  NR2 U432 ( .A(n142), .B(n77), .Z(\ab[8][22] ) );
  NR2 U433 ( .A(n143), .B(n77), .Z(\ab[8][21] ) );
  NR2 U434 ( .A(n144), .B(n77), .Z(\ab[8][20] ) );
  NR2 U435 ( .A(n163), .B(n76), .Z(\ab[8][1] ) );
  NR2 U436 ( .A(n145), .B(n76), .Z(\ab[8][19] ) );
  NR2 U437 ( .A(n146), .B(n76), .Z(\ab[8][18] ) );
  NR2 U438 ( .A(n147), .B(n76), .Z(\ab[8][17] ) );
  NR2 U439 ( .A(n148), .B(n76), .Z(\ab[8][16] ) );
  NR2 U440 ( .A(n149), .B(n76), .Z(\ab[8][15] ) );
  NR2 U441 ( .A(n150), .B(n76), .Z(\ab[8][14] ) );
  NR2 U442 ( .A(n151), .B(n76), .Z(\ab[8][13] ) );
  NR2 U443 ( .A(n152), .B(n76), .Z(\ab[8][12] ) );
  NR2 U444 ( .A(n153), .B(n76), .Z(\ab[8][11] ) );
  NR2 U445 ( .A(n154), .B(n76), .Z(\ab[8][10] ) );
  NR2 U446 ( .A(n164), .B(n76), .Z(\ab[8][0] ) );
  NR2 U447 ( .A(n155), .B(n74), .Z(\ab[7][9] ) );
  NR2 U448 ( .A(n156), .B(n74), .Z(\ab[7][8] ) );
  NR2 U449 ( .A(n157), .B(n74), .Z(\ab[7][7] ) );
  NR2 U450 ( .A(n158), .B(n74), .Z(\ab[7][6] ) );
  NR2 U451 ( .A(n159), .B(n74), .Z(\ab[7][5] ) );
  NR2 U452 ( .A(n160), .B(n74), .Z(\ab[7][4] ) );
  NR2 U453 ( .A(n108), .B(n74), .Z(\ab[7][47] ) );
  NR2 U454 ( .A(n107), .B(n74), .Z(\ab[7][46] ) );
  NR2 U455 ( .A(n106), .B(n74), .Z(\ab[7][45] ) );
  NR2 U456 ( .A(n105), .B(n74), .Z(\ab[7][44] ) );
  NR2 U457 ( .A(n104), .B(n74), .Z(\ab[7][43] ) );
  NR2 U458 ( .A(n103), .B(n74), .Z(\ab[7][42] ) );
  NR2 U459 ( .A(n102), .B(n73), .Z(\ab[7][41] ) );
  NR2 U460 ( .A(n101), .B(n73), .Z(\ab[7][40] ) );
  NR2 U461 ( .A(n161), .B(n73), .Z(\ab[7][3] ) );
  NR2 U462 ( .A(n125), .B(n73), .Z(\ab[7][39] ) );
  NR2 U463 ( .A(n126), .B(n73), .Z(\ab[7][38] ) );
  NR2 U464 ( .A(n127), .B(n73), .Z(\ab[7][37] ) );
  NR2 U465 ( .A(n128), .B(n73), .Z(\ab[7][36] ) );
  NR2 U466 ( .A(n129), .B(n73), .Z(\ab[7][35] ) );
  NR2 U467 ( .A(n130), .B(n73), .Z(\ab[7][34] ) );
  NR2 U468 ( .A(n131), .B(n73), .Z(\ab[7][33] ) );
  NR2 U469 ( .A(n132), .B(n73), .Z(\ab[7][32] ) );
  NR2 U470 ( .A(n133), .B(n73), .Z(\ab[7][31] ) );
  NR2 U471 ( .A(n134), .B(n72), .Z(\ab[7][30] ) );
  NR2 U472 ( .A(n162), .B(n72), .Z(\ab[7][2] ) );
  NR2 U473 ( .A(n135), .B(n72), .Z(\ab[7][29] ) );
  NR2 U474 ( .A(n136), .B(n72), .Z(\ab[7][28] ) );
  NR2 U475 ( .A(n137), .B(n72), .Z(\ab[7][27] ) );
  NR2 U476 ( .A(n138), .B(n72), .Z(\ab[7][26] ) );
  NR2 U477 ( .A(n139), .B(n72), .Z(\ab[7][25] ) );
  NR2 U478 ( .A(n140), .B(n72), .Z(\ab[7][24] ) );
  NR2 U479 ( .A(n141), .B(n72), .Z(\ab[7][23] ) );
  NR2 U480 ( .A(n142), .B(n72), .Z(\ab[7][22] ) );
  NR2 U481 ( .A(n143), .B(n72), .Z(\ab[7][21] ) );
  NR2 U482 ( .A(n144), .B(n72), .Z(\ab[7][20] ) );
  NR2 U483 ( .A(n163), .B(n71), .Z(\ab[7][1] ) );
  NR2 U484 ( .A(n145), .B(n71), .Z(\ab[7][19] ) );
  NR2 U485 ( .A(n146), .B(n71), .Z(\ab[7][18] ) );
  NR2 U486 ( .A(n147), .B(n71), .Z(\ab[7][17] ) );
  NR2 U487 ( .A(n148), .B(n71), .Z(\ab[7][16] ) );
  NR2 U488 ( .A(n149), .B(n71), .Z(\ab[7][15] ) );
  NR2 U489 ( .A(n150), .B(n71), .Z(\ab[7][14] ) );
  NR2 U490 ( .A(n151), .B(n71), .Z(\ab[7][13] ) );
  NR2 U491 ( .A(n152), .B(n71), .Z(\ab[7][12] ) );
  NR2 U492 ( .A(n153), .B(n71), .Z(\ab[7][11] ) );
  NR2 U493 ( .A(n154), .B(n71), .Z(\ab[7][10] ) );
  NR2 U494 ( .A(n164), .B(n71), .Z(\ab[7][0] ) );
  NR2 U495 ( .A(n155), .B(n69), .Z(\ab[6][9] ) );
  NR2 U496 ( .A(n156), .B(n69), .Z(\ab[6][8] ) );
  NR2 U497 ( .A(n157), .B(n69), .Z(\ab[6][7] ) );
  NR2 U498 ( .A(n158), .B(n69), .Z(\ab[6][6] ) );
  NR2 U499 ( .A(n159), .B(n69), .Z(\ab[6][5] ) );
  NR2 U500 ( .A(n160), .B(n69), .Z(\ab[6][4] ) );
  NR2 U501 ( .A(n108), .B(n69), .Z(\ab[6][47] ) );
  NR2 U502 ( .A(n107), .B(n69), .Z(\ab[6][46] ) );
  NR2 U503 ( .A(n106), .B(n69), .Z(\ab[6][45] ) );
  NR2 U504 ( .A(n105), .B(n69), .Z(\ab[6][44] ) );
  NR2 U505 ( .A(n104), .B(n69), .Z(\ab[6][43] ) );
  NR2 U506 ( .A(n103), .B(n69), .Z(\ab[6][42] ) );
  NR2 U507 ( .A(n102), .B(n68), .Z(\ab[6][41] ) );
  NR2 U508 ( .A(n101), .B(n68), .Z(\ab[6][40] ) );
  NR2 U509 ( .A(n161), .B(n68), .Z(\ab[6][3] ) );
  NR2 U510 ( .A(n125), .B(n68), .Z(\ab[6][39] ) );
  NR2 U511 ( .A(n126), .B(n68), .Z(\ab[6][38] ) );
  NR2 U512 ( .A(n127), .B(n68), .Z(\ab[6][37] ) );
  NR2 U513 ( .A(n128), .B(n68), .Z(\ab[6][36] ) );
  NR2 U514 ( .A(n129), .B(n68), .Z(\ab[6][35] ) );
  NR2 U515 ( .A(n130), .B(n68), .Z(\ab[6][34] ) );
  NR2 U516 ( .A(n131), .B(n68), .Z(\ab[6][33] ) );
  NR2 U517 ( .A(n132), .B(n68), .Z(\ab[6][32] ) );
  NR2 U518 ( .A(n133), .B(n68), .Z(\ab[6][31] ) );
  NR2 U519 ( .A(n134), .B(n67), .Z(\ab[6][30] ) );
  NR2 U520 ( .A(n162), .B(n67), .Z(\ab[6][2] ) );
  NR2 U521 ( .A(n135), .B(n67), .Z(\ab[6][29] ) );
  NR2 U522 ( .A(n136), .B(n67), .Z(\ab[6][28] ) );
  NR2 U523 ( .A(n137), .B(n67), .Z(\ab[6][27] ) );
  NR2 U524 ( .A(n138), .B(n67), .Z(\ab[6][26] ) );
  NR2 U525 ( .A(n139), .B(n67), .Z(\ab[6][25] ) );
  NR2 U526 ( .A(n140), .B(n67), .Z(\ab[6][24] ) );
  NR2 U527 ( .A(n141), .B(n67), .Z(\ab[6][23] ) );
  NR2 U528 ( .A(n142), .B(n67), .Z(\ab[6][22] ) );
  NR2 U529 ( .A(n143), .B(n67), .Z(\ab[6][21] ) );
  NR2 U530 ( .A(n144), .B(n67), .Z(\ab[6][20] ) );
  NR2 U531 ( .A(n163), .B(n66), .Z(\ab[6][1] ) );
  NR2 U532 ( .A(n145), .B(n66), .Z(\ab[6][19] ) );
  NR2 U533 ( .A(n146), .B(n66), .Z(\ab[6][18] ) );
  NR2 U534 ( .A(n147), .B(n66), .Z(\ab[6][17] ) );
  NR2 U535 ( .A(n148), .B(n66), .Z(\ab[6][16] ) );
  NR2 U536 ( .A(n149), .B(n66), .Z(\ab[6][15] ) );
  NR2 U537 ( .A(n150), .B(n66), .Z(\ab[6][14] ) );
  NR2 U538 ( .A(n151), .B(n66), .Z(\ab[6][13] ) );
  NR2 U539 ( .A(n152), .B(n66), .Z(\ab[6][12] ) );
  NR2 U540 ( .A(n153), .B(n66), .Z(\ab[6][11] ) );
  NR2 U541 ( .A(n154), .B(n66), .Z(\ab[6][10] ) );
  NR2 U542 ( .A(n164), .B(n66), .Z(\ab[6][0] ) );
  NR2 U543 ( .A(n155), .B(n64), .Z(\ab[5][9] ) );
  NR2 U544 ( .A(n156), .B(n64), .Z(\ab[5][8] ) );
  NR2 U545 ( .A(n157), .B(n64), .Z(\ab[5][7] ) );
  NR2 U546 ( .A(n158), .B(n64), .Z(\ab[5][6] ) );
  NR2 U547 ( .A(n159), .B(n64), .Z(\ab[5][5] ) );
  NR2 U548 ( .A(n160), .B(n64), .Z(\ab[5][4] ) );
  NR2 U549 ( .A(n108), .B(n64), .Z(\ab[5][47] ) );
  NR2 U550 ( .A(n107), .B(n64), .Z(\ab[5][46] ) );
  NR2 U551 ( .A(n106), .B(n64), .Z(\ab[5][45] ) );
  NR2 U552 ( .A(n105), .B(n64), .Z(\ab[5][44] ) );
  NR2 U553 ( .A(n104), .B(n64), .Z(\ab[5][43] ) );
  NR2 U554 ( .A(n103), .B(n64), .Z(\ab[5][42] ) );
  NR2 U555 ( .A(n102), .B(n63), .Z(\ab[5][41] ) );
  NR2 U556 ( .A(n101), .B(n63), .Z(\ab[5][40] ) );
  NR2 U557 ( .A(n161), .B(n63), .Z(\ab[5][3] ) );
  NR2 U558 ( .A(n125), .B(n63), .Z(\ab[5][39] ) );
  NR2 U559 ( .A(n126), .B(n63), .Z(\ab[5][38] ) );
  NR2 U560 ( .A(n127), .B(n63), .Z(\ab[5][37] ) );
  NR2 U561 ( .A(n128), .B(n63), .Z(\ab[5][36] ) );
  NR2 U562 ( .A(n129), .B(n63), .Z(\ab[5][35] ) );
  NR2 U563 ( .A(n130), .B(n63), .Z(\ab[5][34] ) );
  NR2 U564 ( .A(n131), .B(n63), .Z(\ab[5][33] ) );
  NR2 U565 ( .A(n132), .B(n63), .Z(\ab[5][32] ) );
  NR2 U566 ( .A(n133), .B(n63), .Z(\ab[5][31] ) );
  NR2 U567 ( .A(n134), .B(n62), .Z(\ab[5][30] ) );
  NR2 U568 ( .A(n162), .B(n62), .Z(\ab[5][2] ) );
  NR2 U569 ( .A(n135), .B(n62), .Z(\ab[5][29] ) );
  NR2 U570 ( .A(n136), .B(n62), .Z(\ab[5][28] ) );
  NR2 U571 ( .A(n137), .B(n62), .Z(\ab[5][27] ) );
  NR2 U572 ( .A(n138), .B(n62), .Z(\ab[5][26] ) );
  NR2 U573 ( .A(n139), .B(n62), .Z(\ab[5][25] ) );
  NR2 U574 ( .A(n140), .B(n62), .Z(\ab[5][24] ) );
  NR2 U575 ( .A(n141), .B(n62), .Z(\ab[5][23] ) );
  NR2 U576 ( .A(n142), .B(n62), .Z(\ab[5][22] ) );
  NR2 U577 ( .A(n143), .B(n62), .Z(\ab[5][21] ) );
  NR2 U578 ( .A(n144), .B(n62), .Z(\ab[5][20] ) );
  NR2 U579 ( .A(n163), .B(n61), .Z(\ab[5][1] ) );
  NR2 U580 ( .A(n145), .B(n61), .Z(\ab[5][19] ) );
  NR2 U581 ( .A(n146), .B(n61), .Z(\ab[5][18] ) );
  NR2 U582 ( .A(n147), .B(n61), .Z(\ab[5][17] ) );
  NR2 U583 ( .A(n148), .B(n61), .Z(\ab[5][16] ) );
  NR2 U584 ( .A(n149), .B(n61), .Z(\ab[5][15] ) );
  NR2 U585 ( .A(n150), .B(n61), .Z(\ab[5][14] ) );
  NR2 U586 ( .A(n151), .B(n61), .Z(\ab[5][13] ) );
  NR2 U587 ( .A(n152), .B(n61), .Z(\ab[5][12] ) );
  NR2 U588 ( .A(n153), .B(n61), .Z(\ab[5][11] ) );
  NR2 U589 ( .A(n154), .B(n61), .Z(\ab[5][10] ) );
  NR2 U590 ( .A(n164), .B(n61), .Z(\ab[5][0] ) );
  NR2 U591 ( .A(n155), .B(n59), .Z(\ab[4][9] ) );
  NR2 U592 ( .A(n156), .B(n59), .Z(\ab[4][8] ) );
  NR2 U593 ( .A(n157), .B(n59), .Z(\ab[4][7] ) );
  NR2 U594 ( .A(n158), .B(n59), .Z(\ab[4][6] ) );
  NR2 U595 ( .A(n159), .B(n59), .Z(\ab[4][5] ) );
  NR2 U596 ( .A(n160), .B(n59), .Z(\ab[4][4] ) );
  NR2 U597 ( .A(n108), .B(n59), .Z(\ab[4][47] ) );
  NR2 U598 ( .A(n107), .B(n59), .Z(\ab[4][46] ) );
  NR2 U599 ( .A(n106), .B(n59), .Z(\ab[4][45] ) );
  NR2 U600 ( .A(n105), .B(n59), .Z(\ab[4][44] ) );
  NR2 U601 ( .A(n104), .B(n59), .Z(\ab[4][43] ) );
  NR2 U602 ( .A(n103), .B(n59), .Z(\ab[4][42] ) );
  NR2 U603 ( .A(n102), .B(n58), .Z(\ab[4][41] ) );
  NR2 U604 ( .A(n101), .B(n58), .Z(\ab[4][40] ) );
  NR2 U605 ( .A(n161), .B(n58), .Z(\ab[4][3] ) );
  NR2 U606 ( .A(n125), .B(n58), .Z(\ab[4][39] ) );
  NR2 U607 ( .A(n126), .B(n58), .Z(\ab[4][38] ) );
  NR2 U608 ( .A(n127), .B(n58), .Z(\ab[4][37] ) );
  NR2 U609 ( .A(n128), .B(n58), .Z(\ab[4][36] ) );
  NR2 U610 ( .A(n129), .B(n58), .Z(\ab[4][35] ) );
  NR2 U611 ( .A(n130), .B(n58), .Z(\ab[4][34] ) );
  NR2 U612 ( .A(n131), .B(n58), .Z(\ab[4][33] ) );
  NR2 U613 ( .A(n132), .B(n58), .Z(\ab[4][32] ) );
  NR2 U614 ( .A(n133), .B(n58), .Z(\ab[4][31] ) );
  NR2 U615 ( .A(n134), .B(n57), .Z(\ab[4][30] ) );
  NR2 U616 ( .A(n162), .B(n57), .Z(\ab[4][2] ) );
  NR2 U617 ( .A(n135), .B(n57), .Z(\ab[4][29] ) );
  NR2 U618 ( .A(n136), .B(n57), .Z(\ab[4][28] ) );
  NR2 U619 ( .A(n137), .B(n57), .Z(\ab[4][27] ) );
  NR2 U620 ( .A(n138), .B(n57), .Z(\ab[4][26] ) );
  NR2 U621 ( .A(n139), .B(n57), .Z(\ab[4][25] ) );
  NR2 U622 ( .A(n140), .B(n57), .Z(\ab[4][24] ) );
  NR2 U623 ( .A(n141), .B(n57), .Z(\ab[4][23] ) );
  NR2 U624 ( .A(n142), .B(n57), .Z(\ab[4][22] ) );
  NR2 U625 ( .A(n143), .B(n57), .Z(\ab[4][21] ) );
  NR2 U626 ( .A(n144), .B(n57), .Z(\ab[4][20] ) );
  NR2 U627 ( .A(n163), .B(n56), .Z(\ab[4][1] ) );
  NR2 U628 ( .A(n145), .B(n56), .Z(\ab[4][19] ) );
  NR2 U629 ( .A(n146), .B(n56), .Z(\ab[4][18] ) );
  NR2 U630 ( .A(n147), .B(n56), .Z(\ab[4][17] ) );
  NR2 U631 ( .A(n148), .B(n56), .Z(\ab[4][16] ) );
  NR2 U632 ( .A(n149), .B(n56), .Z(\ab[4][15] ) );
  NR2 U633 ( .A(n150), .B(n56), .Z(\ab[4][14] ) );
  NR2 U634 ( .A(n151), .B(n56), .Z(\ab[4][13] ) );
  NR2 U635 ( .A(n152), .B(n56), .Z(\ab[4][12] ) );
  NR2 U636 ( .A(n153), .B(n56), .Z(\ab[4][11] ) );
  NR2 U637 ( .A(n154), .B(n56), .Z(\ab[4][10] ) );
  NR2 U638 ( .A(n164), .B(n56), .Z(\ab[4][0] ) );
  NR2 U639 ( .A(n155), .B(n54), .Z(\ab[3][9] ) );
  NR2 U640 ( .A(n156), .B(n54), .Z(\ab[3][8] ) );
  NR2 U641 ( .A(n157), .B(n54), .Z(\ab[3][7] ) );
  NR2 U642 ( .A(n158), .B(n54), .Z(\ab[3][6] ) );
  NR2 U643 ( .A(n159), .B(n54), .Z(\ab[3][5] ) );
  NR2 U644 ( .A(n160), .B(n54), .Z(\ab[3][4] ) );
  NR2 U645 ( .A(n108), .B(n54), .Z(\ab[3][47] ) );
  NR2 U646 ( .A(n107), .B(n54), .Z(\ab[3][46] ) );
  NR2 U647 ( .A(n106), .B(n54), .Z(\ab[3][45] ) );
  NR2 U648 ( .A(n105), .B(n54), .Z(\ab[3][44] ) );
  NR2 U649 ( .A(n104), .B(n54), .Z(\ab[3][43] ) );
  NR2 U650 ( .A(n103), .B(n54), .Z(\ab[3][42] ) );
  NR2 U651 ( .A(n102), .B(n53), .Z(\ab[3][41] ) );
  NR2 U652 ( .A(n101), .B(n53), .Z(\ab[3][40] ) );
  NR2 U653 ( .A(n161), .B(n53), .Z(\ab[3][3] ) );
  NR2 U654 ( .A(n125), .B(n53), .Z(\ab[3][39] ) );
  NR2 U655 ( .A(n126), .B(n53), .Z(\ab[3][38] ) );
  NR2 U656 ( .A(n127), .B(n53), .Z(\ab[3][37] ) );
  NR2 U657 ( .A(n128), .B(n53), .Z(\ab[3][36] ) );
  NR2 U658 ( .A(n129), .B(n53), .Z(\ab[3][35] ) );
  NR2 U659 ( .A(n130), .B(n53), .Z(\ab[3][34] ) );
  NR2 U660 ( .A(n131), .B(n53), .Z(\ab[3][33] ) );
  NR2 U661 ( .A(n132), .B(n53), .Z(\ab[3][32] ) );
  NR2 U662 ( .A(n133), .B(n53), .Z(\ab[3][31] ) );
  NR2 U663 ( .A(n134), .B(n52), .Z(\ab[3][30] ) );
  NR2 U664 ( .A(n162), .B(n52), .Z(\ab[3][2] ) );
  NR2 U665 ( .A(n135), .B(n52), .Z(\ab[3][29] ) );
  NR2 U666 ( .A(n136), .B(n52), .Z(\ab[3][28] ) );
  NR2 U667 ( .A(n137), .B(n52), .Z(\ab[3][27] ) );
  NR2 U668 ( .A(n138), .B(n52), .Z(\ab[3][26] ) );
  NR2 U669 ( .A(n139), .B(n52), .Z(\ab[3][25] ) );
  NR2 U670 ( .A(n140), .B(n52), .Z(\ab[3][24] ) );
  NR2 U671 ( .A(n141), .B(n52), .Z(\ab[3][23] ) );
  NR2 U672 ( .A(n142), .B(n52), .Z(\ab[3][22] ) );
  NR2 U673 ( .A(n143), .B(n52), .Z(\ab[3][21] ) );
  NR2 U674 ( .A(n144), .B(n52), .Z(\ab[3][20] ) );
  NR2 U675 ( .A(n163), .B(n51), .Z(\ab[3][1] ) );
  NR2 U676 ( .A(n145), .B(n51), .Z(\ab[3][19] ) );
  NR2 U677 ( .A(n146), .B(n51), .Z(\ab[3][18] ) );
  NR2 U678 ( .A(n147), .B(n51), .Z(\ab[3][17] ) );
  NR2 U679 ( .A(n148), .B(n51), .Z(\ab[3][16] ) );
  NR2 U680 ( .A(n149), .B(n51), .Z(\ab[3][15] ) );
  NR2 U681 ( .A(n150), .B(n51), .Z(\ab[3][14] ) );
  NR2 U682 ( .A(n151), .B(n51), .Z(\ab[3][13] ) );
  NR2 U683 ( .A(n152), .B(n51), .Z(\ab[3][12] ) );
  NR2 U684 ( .A(n153), .B(n51), .Z(\ab[3][11] ) );
  NR2 U685 ( .A(n154), .B(n51), .Z(\ab[3][10] ) );
  NR2 U686 ( .A(n164), .B(n51), .Z(\ab[3][0] ) );
  NR2 U687 ( .A(n155), .B(n49), .Z(\ab[2][9] ) );
  NR2 U688 ( .A(n156), .B(n49), .Z(\ab[2][8] ) );
  NR2 U689 ( .A(n157), .B(n49), .Z(\ab[2][7] ) );
  NR2 U690 ( .A(n158), .B(n49), .Z(\ab[2][6] ) );
  NR2 U691 ( .A(n159), .B(n49), .Z(\ab[2][5] ) );
  NR2 U692 ( .A(n160), .B(n49), .Z(\ab[2][4] ) );
  NR2 U693 ( .A(n108), .B(n49), .Z(\ab[2][47] ) );
  NR2 U694 ( .A(n107), .B(n49), .Z(\ab[2][46] ) );
  NR2 U695 ( .A(n106), .B(n49), .Z(\ab[2][45] ) );
  NR2 U696 ( .A(n105), .B(n49), .Z(\ab[2][44] ) );
  NR2 U697 ( .A(n104), .B(n49), .Z(\ab[2][43] ) );
  NR2 U698 ( .A(n103), .B(n49), .Z(\ab[2][42] ) );
  NR2 U699 ( .A(n102), .B(n48), .Z(\ab[2][41] ) );
  NR2 U700 ( .A(n101), .B(n48), .Z(\ab[2][40] ) );
  NR2 U701 ( .A(n161), .B(n48), .Z(\ab[2][3] ) );
  NR2 U702 ( .A(n125), .B(n48), .Z(\ab[2][39] ) );
  NR2 U703 ( .A(n126), .B(n48), .Z(\ab[2][38] ) );
  NR2 U704 ( .A(n127), .B(n48), .Z(\ab[2][37] ) );
  NR2 U705 ( .A(n128), .B(n48), .Z(\ab[2][36] ) );
  NR2 U706 ( .A(n129), .B(n48), .Z(\ab[2][35] ) );
  NR2 U707 ( .A(n130), .B(n48), .Z(\ab[2][34] ) );
  NR2 U708 ( .A(n131), .B(n48), .Z(\ab[2][33] ) );
  NR2 U709 ( .A(n132), .B(n48), .Z(\ab[2][32] ) );
  NR2 U710 ( .A(n133), .B(n48), .Z(\ab[2][31] ) );
  NR2 U711 ( .A(n134), .B(n47), .Z(\ab[2][30] ) );
  NR2 U712 ( .A(n162), .B(n47), .Z(\ab[2][2] ) );
  NR2 U713 ( .A(n135), .B(n47), .Z(\ab[2][29] ) );
  NR2 U714 ( .A(n136), .B(n47), .Z(\ab[2][28] ) );
  NR2 U715 ( .A(n137), .B(n47), .Z(\ab[2][27] ) );
  NR2 U716 ( .A(n138), .B(n47), .Z(\ab[2][26] ) );
  NR2 U717 ( .A(n139), .B(n47), .Z(\ab[2][25] ) );
  NR2 U718 ( .A(n140), .B(n47), .Z(\ab[2][24] ) );
  NR2 U719 ( .A(n141), .B(n47), .Z(\ab[2][23] ) );
  NR2 U720 ( .A(n142), .B(n47), .Z(\ab[2][22] ) );
  NR2 U721 ( .A(n143), .B(n47), .Z(\ab[2][21] ) );
  NR2 U722 ( .A(n144), .B(n47), .Z(\ab[2][20] ) );
  NR2 U723 ( .A(n163), .B(n46), .Z(\ab[2][1] ) );
  NR2 U724 ( .A(n145), .B(n46), .Z(\ab[2][19] ) );
  NR2 U725 ( .A(n146), .B(n46), .Z(\ab[2][18] ) );
  NR2 U726 ( .A(n147), .B(n46), .Z(\ab[2][17] ) );
  NR2 U727 ( .A(n148), .B(n46), .Z(\ab[2][16] ) );
  NR2 U728 ( .A(n149), .B(n46), .Z(\ab[2][15] ) );
  NR2 U729 ( .A(n150), .B(n46), .Z(\ab[2][14] ) );
  NR2 U730 ( .A(n151), .B(n46), .Z(\ab[2][13] ) );
  NR2 U731 ( .A(n152), .B(n46), .Z(\ab[2][12] ) );
  NR2 U732 ( .A(n153), .B(n46), .Z(\ab[2][11] ) );
  NR2 U733 ( .A(n154), .B(n46), .Z(\ab[2][10] ) );
  NR2 U734 ( .A(n164), .B(n46), .Z(\ab[2][0] ) );
  NR2 U735 ( .A(n155), .B(n11), .Z(\ab[21][9] ) );
  NR2 U736 ( .A(n156), .B(n11), .Z(\ab[21][8] ) );
  NR2 U737 ( .A(n157), .B(n11), .Z(\ab[21][7] ) );
  NR2 U738 ( .A(n158), .B(n11), .Z(\ab[21][6] ) );
  NR2 U739 ( .A(n159), .B(n11), .Z(\ab[21][5] ) );
  NR2 U740 ( .A(n160), .B(n11), .Z(\ab[21][4] ) );
  NR2 U741 ( .A(n108), .B(n11), .Z(\ab[21][47] ) );
  NR2 U742 ( .A(n107), .B(n11), .Z(\ab[21][46] ) );
  NR2 U743 ( .A(n106), .B(n11), .Z(\ab[21][45] ) );
  NR2 U744 ( .A(n105), .B(n11), .Z(\ab[21][44] ) );
  NR2 U745 ( .A(n104), .B(n11), .Z(\ab[21][43] ) );
  NR2 U746 ( .A(n103), .B(n11), .Z(\ab[21][42] ) );
  NR2 U747 ( .A(n102), .B(n10), .Z(\ab[21][41] ) );
  NR2 U748 ( .A(n101), .B(n10), .Z(\ab[21][40] ) );
  NR2 U749 ( .A(n161), .B(n10), .Z(\ab[21][3] ) );
  NR2 U750 ( .A(n125), .B(n10), .Z(\ab[21][39] ) );
  NR2 U751 ( .A(n126), .B(n10), .Z(\ab[21][38] ) );
  NR2 U752 ( .A(n127), .B(n10), .Z(\ab[21][37] ) );
  NR2 U753 ( .A(n128), .B(n10), .Z(\ab[21][36] ) );
  NR2 U754 ( .A(n129), .B(n10), .Z(\ab[21][35] ) );
  NR2 U755 ( .A(n130), .B(n10), .Z(\ab[21][34] ) );
  NR2 U756 ( .A(n131), .B(n10), .Z(\ab[21][33] ) );
  NR2 U757 ( .A(n132), .B(n10), .Z(\ab[21][32] ) );
  NR2 U758 ( .A(n133), .B(n10), .Z(\ab[21][31] ) );
  NR2 U759 ( .A(n134), .B(n9), .Z(\ab[21][30] ) );
  NR2 U760 ( .A(n162), .B(n9), .Z(\ab[21][2] ) );
  NR2 U761 ( .A(n135), .B(n9), .Z(\ab[21][29] ) );
  NR2 U762 ( .A(n136), .B(n9), .Z(\ab[21][28] ) );
  NR2 U763 ( .A(n137), .B(n9), .Z(\ab[21][27] ) );
  NR2 U764 ( .A(n138), .B(n9), .Z(\ab[21][26] ) );
  NR2 U765 ( .A(n139), .B(n9), .Z(\ab[21][25] ) );
  NR2 U766 ( .A(n140), .B(n9), .Z(\ab[21][24] ) );
  NR2 U767 ( .A(n141), .B(n9), .Z(\ab[21][23] ) );
  NR2 U768 ( .A(n142), .B(n9), .Z(\ab[21][22] ) );
  NR2 U769 ( .A(n143), .B(n9), .Z(\ab[21][21] ) );
  NR2 U770 ( .A(n144), .B(n9), .Z(\ab[21][20] ) );
  NR2 U771 ( .A(n163), .B(n8), .Z(\ab[21][1] ) );
  NR2 U772 ( .A(n145), .B(n8), .Z(\ab[21][19] ) );
  NR2 U773 ( .A(n146), .B(n8), .Z(\ab[21][18] ) );
  NR2 U774 ( .A(n147), .B(n8), .Z(\ab[21][17] ) );
  NR2 U775 ( .A(n148), .B(n8), .Z(\ab[21][16] ) );
  NR2 U776 ( .A(n149), .B(n8), .Z(\ab[21][15] ) );
  NR2 U777 ( .A(n150), .B(n8), .Z(\ab[21][14] ) );
  NR2 U778 ( .A(n151), .B(n8), .Z(\ab[21][13] ) );
  NR2 U779 ( .A(n152), .B(n8), .Z(\ab[21][12] ) );
  NR2 U780 ( .A(n153), .B(n8), .Z(\ab[21][11] ) );
  NR2 U781 ( .A(n154), .B(n8), .Z(\ab[21][10] ) );
  NR2 U782 ( .A(n164), .B(n8), .Z(\ab[21][0] ) );
  NR2 U783 ( .A(n155), .B(n15), .Z(\ab[20][9] ) );
  NR2 U784 ( .A(n156), .B(n15), .Z(\ab[20][8] ) );
  NR2 U785 ( .A(n157), .B(n15), .Z(\ab[20][7] ) );
  NR2 U786 ( .A(n158), .B(n15), .Z(\ab[20][6] ) );
  NR2 U787 ( .A(n159), .B(n15), .Z(\ab[20][5] ) );
  NR2 U788 ( .A(n160), .B(n15), .Z(\ab[20][4] ) );
  NR2 U789 ( .A(n108), .B(n15), .Z(\ab[20][47] ) );
  NR2 U790 ( .A(n107), .B(n15), .Z(\ab[20][46] ) );
  NR2 U791 ( .A(n106), .B(n15), .Z(\ab[20][45] ) );
  NR2 U792 ( .A(n105), .B(n15), .Z(\ab[20][44] ) );
  NR2 U793 ( .A(n104), .B(n15), .Z(\ab[20][43] ) );
  NR2 U794 ( .A(n103), .B(n15), .Z(\ab[20][42] ) );
  NR2 U795 ( .A(n102), .B(n14), .Z(\ab[20][41] ) );
  NR2 U796 ( .A(n101), .B(n14), .Z(\ab[20][40] ) );
  NR2 U797 ( .A(n161), .B(n14), .Z(\ab[20][3] ) );
  NR2 U798 ( .A(n125), .B(n14), .Z(\ab[20][39] ) );
  NR2 U799 ( .A(n126), .B(n14), .Z(\ab[20][38] ) );
  NR2 U800 ( .A(n127), .B(n14), .Z(\ab[20][37] ) );
  NR2 U801 ( .A(n128), .B(n14), .Z(\ab[20][36] ) );
  NR2 U802 ( .A(n129), .B(n14), .Z(\ab[20][35] ) );
  NR2 U803 ( .A(n130), .B(n14), .Z(\ab[20][34] ) );
  NR2 U804 ( .A(n131), .B(n14), .Z(\ab[20][33] ) );
  NR2 U805 ( .A(n132), .B(n14), .Z(\ab[20][32] ) );
  NR2 U806 ( .A(n133), .B(n14), .Z(\ab[20][31] ) );
  NR2 U807 ( .A(n134), .B(n13), .Z(\ab[20][30] ) );
  NR2 U808 ( .A(n162), .B(n13), .Z(\ab[20][2] ) );
  NR2 U809 ( .A(n135), .B(n13), .Z(\ab[20][29] ) );
  NR2 U810 ( .A(n136), .B(n13), .Z(\ab[20][28] ) );
  NR2 U811 ( .A(n137), .B(n13), .Z(\ab[20][27] ) );
  NR2 U812 ( .A(n138), .B(n13), .Z(\ab[20][26] ) );
  NR2 U813 ( .A(n139), .B(n13), .Z(\ab[20][25] ) );
  NR2 U814 ( .A(n140), .B(n13), .Z(\ab[20][24] ) );
  NR2 U815 ( .A(n141), .B(n13), .Z(\ab[20][23] ) );
  NR2 U816 ( .A(n142), .B(n13), .Z(\ab[20][22] ) );
  NR2 U817 ( .A(n143), .B(n13), .Z(\ab[20][21] ) );
  NR2 U818 ( .A(n144), .B(n13), .Z(\ab[20][20] ) );
  NR2 U819 ( .A(n163), .B(n12), .Z(\ab[20][1] ) );
  NR2 U820 ( .A(n145), .B(n12), .Z(\ab[20][19] ) );
  NR2 U821 ( .A(n146), .B(n12), .Z(\ab[20][18] ) );
  NR2 U822 ( .A(n147), .B(n12), .Z(\ab[20][17] ) );
  NR2 U823 ( .A(n148), .B(n12), .Z(\ab[20][16] ) );
  NR2 U824 ( .A(n149), .B(n12), .Z(\ab[20][15] ) );
  NR2 U825 ( .A(n150), .B(n12), .Z(\ab[20][14] ) );
  NR2 U826 ( .A(n151), .B(n12), .Z(\ab[20][13] ) );
  NR2 U827 ( .A(n152), .B(n12), .Z(\ab[20][12] ) );
  NR2 U828 ( .A(n153), .B(n12), .Z(\ab[20][11] ) );
  NR2 U829 ( .A(n154), .B(n12), .Z(\ab[20][10] ) );
  NR2 U830 ( .A(n164), .B(n12), .Z(\ab[20][0] ) );
  NR2 U831 ( .A(n155), .B(n44), .Z(\ab[1][9] ) );
  NR2 U832 ( .A(n156), .B(n44), .Z(\ab[1][8] ) );
  NR2 U833 ( .A(n157), .B(n44), .Z(\ab[1][7] ) );
  NR2 U834 ( .A(n158), .B(n44), .Z(\ab[1][6] ) );
  NR2 U835 ( .A(n159), .B(n44), .Z(\ab[1][5] ) );
  NR2 U836 ( .A(n160), .B(n44), .Z(\ab[1][4] ) );
  NR2 U837 ( .A(n108), .B(n44), .Z(\ab[1][47] ) );
  NR2 U838 ( .A(n107), .B(n44), .Z(\ab[1][46] ) );
  NR2 U839 ( .A(n106), .B(n44), .Z(\ab[1][45] ) );
  NR2 U840 ( .A(n105), .B(n44), .Z(\ab[1][44] ) );
  NR2 U841 ( .A(n104), .B(n44), .Z(\ab[1][43] ) );
  NR2 U842 ( .A(n103), .B(n43), .Z(\ab[1][42] ) );
  NR2 U843 ( .A(n102), .B(n43), .Z(\ab[1][41] ) );
  NR2 U844 ( .A(n101), .B(n43), .Z(\ab[1][40] ) );
  NR2 U845 ( .A(n161), .B(n43), .Z(\ab[1][3] ) );
  NR2 U846 ( .A(n125), .B(n43), .Z(\ab[1][39] ) );
  NR2 U847 ( .A(n126), .B(n43), .Z(\ab[1][38] ) );
  NR2 U848 ( .A(n127), .B(n43), .Z(\ab[1][37] ) );
  NR2 U849 ( .A(n128), .B(n43), .Z(\ab[1][36] ) );
  NR2 U850 ( .A(n129), .B(n43), .Z(\ab[1][35] ) );
  NR2 U851 ( .A(n130), .B(n43), .Z(\ab[1][34] ) );
  NR2 U852 ( .A(n131), .B(n43), .Z(\ab[1][33] ) );
  NR2 U853 ( .A(n132), .B(n43), .Z(\ab[1][32] ) );
  NR2 U854 ( .A(n133), .B(n42), .Z(\ab[1][31] ) );
  NR2 U855 ( .A(n134), .B(n42), .Z(\ab[1][30] ) );
  NR2 U856 ( .A(n162), .B(n42), .Z(\ab[1][2] ) );
  NR2 U857 ( .A(n135), .B(n42), .Z(\ab[1][29] ) );
  NR2 U858 ( .A(n136), .B(n42), .Z(\ab[1][28] ) );
  NR2 U859 ( .A(n137), .B(n42), .Z(\ab[1][27] ) );
  NR2 U860 ( .A(n138), .B(n42), .Z(\ab[1][26] ) );
  NR2 U861 ( .A(n139), .B(n42), .Z(\ab[1][25] ) );
  NR2 U862 ( .A(n140), .B(n42), .Z(\ab[1][24] ) );
  NR2 U863 ( .A(n141), .B(n42), .Z(\ab[1][23] ) );
  NR2 U864 ( .A(n142), .B(n42), .Z(\ab[1][22] ) );
  NR2 U865 ( .A(n143), .B(n42), .Z(\ab[1][21] ) );
  NR2 U866 ( .A(n144), .B(n41), .Z(\ab[1][20] ) );
  NR2 U867 ( .A(n145), .B(n41), .Z(\ab[1][19] ) );
  NR2 U868 ( .A(n146), .B(n41), .Z(\ab[1][18] ) );
  NR2 U869 ( .A(n147), .B(n41), .Z(\ab[1][17] ) );
  NR2 U870 ( .A(n148), .B(n41), .Z(\ab[1][16] ) );
  NR2 U871 ( .A(n149), .B(n41), .Z(\ab[1][15] ) );
  NR2 U872 ( .A(n150), .B(n41), .Z(\ab[1][14] ) );
  NR2 U873 ( .A(n151), .B(n41), .Z(\ab[1][13] ) );
  NR2 U874 ( .A(n152), .B(n41), .Z(\ab[1][12] ) );
  NR2 U875 ( .A(n153), .B(n41), .Z(\ab[1][11] ) );
  NR2 U876 ( .A(n154), .B(n41), .Z(\ab[1][10] ) );
  NR2 U877 ( .A(n155), .B(n19), .Z(\ab[19][9] ) );
  NR2 U878 ( .A(n156), .B(n19), .Z(\ab[19][8] ) );
  NR2 U879 ( .A(n157), .B(n19), .Z(\ab[19][7] ) );
  NR2 U880 ( .A(n158), .B(n19), .Z(\ab[19][6] ) );
  NR2 U881 ( .A(n159), .B(n19), .Z(\ab[19][5] ) );
  NR2 U882 ( .A(n160), .B(n19), .Z(\ab[19][4] ) );
  NR2 U883 ( .A(n108), .B(n19), .Z(\ab[19][47] ) );
  NR2 U884 ( .A(n107), .B(n19), .Z(\ab[19][46] ) );
  NR2 U885 ( .A(n106), .B(n19), .Z(\ab[19][45] ) );
  NR2 U886 ( .A(n105), .B(n19), .Z(\ab[19][44] ) );
  NR2 U887 ( .A(n104), .B(n19), .Z(\ab[19][43] ) );
  NR2 U888 ( .A(n103), .B(n19), .Z(\ab[19][42] ) );
  NR2 U889 ( .A(n102), .B(n18), .Z(\ab[19][41] ) );
  NR2 U890 ( .A(n101), .B(n18), .Z(\ab[19][40] ) );
  NR2 U891 ( .A(n161), .B(n18), .Z(\ab[19][3] ) );
  NR2 U892 ( .A(n125), .B(n18), .Z(\ab[19][39] ) );
  NR2 U893 ( .A(n126), .B(n18), .Z(\ab[19][38] ) );
  NR2 U894 ( .A(n127), .B(n18), .Z(\ab[19][37] ) );
  NR2 U895 ( .A(n128), .B(n18), .Z(\ab[19][36] ) );
  NR2 U896 ( .A(n129), .B(n18), .Z(\ab[19][35] ) );
  NR2 U897 ( .A(n130), .B(n18), .Z(\ab[19][34] ) );
  NR2 U898 ( .A(n131), .B(n18), .Z(\ab[19][33] ) );
  NR2 U899 ( .A(n132), .B(n18), .Z(\ab[19][32] ) );
  NR2 U900 ( .A(n133), .B(n18), .Z(\ab[19][31] ) );
  NR2 U901 ( .A(n134), .B(n17), .Z(\ab[19][30] ) );
  NR2 U902 ( .A(n162), .B(n17), .Z(\ab[19][2] ) );
  NR2 U903 ( .A(n135), .B(n17), .Z(\ab[19][29] ) );
  NR2 U904 ( .A(n136), .B(n17), .Z(\ab[19][28] ) );
  NR2 U905 ( .A(n137), .B(n17), .Z(\ab[19][27] ) );
  NR2 U906 ( .A(n138), .B(n17), .Z(\ab[19][26] ) );
  NR2 U907 ( .A(n139), .B(n17), .Z(\ab[19][25] ) );
  NR2 U908 ( .A(n140), .B(n17), .Z(\ab[19][24] ) );
  NR2 U909 ( .A(n141), .B(n17), .Z(\ab[19][23] ) );
  NR2 U910 ( .A(n142), .B(n17), .Z(\ab[19][22] ) );
  NR2 U911 ( .A(n143), .B(n17), .Z(\ab[19][21] ) );
  NR2 U912 ( .A(n144), .B(n17), .Z(\ab[19][20] ) );
  NR2 U913 ( .A(n163), .B(n16), .Z(\ab[19][1] ) );
  NR2 U914 ( .A(n145), .B(n16), .Z(\ab[19][19] ) );
  NR2 U915 ( .A(n146), .B(n16), .Z(\ab[19][18] ) );
  NR2 U916 ( .A(n147), .B(n16), .Z(\ab[19][17] ) );
  NR2 U917 ( .A(n148), .B(n16), .Z(\ab[19][16] ) );
  NR2 U918 ( .A(n149), .B(n16), .Z(\ab[19][15] ) );
  NR2 U919 ( .A(n150), .B(n16), .Z(\ab[19][14] ) );
  NR2 U920 ( .A(n151), .B(n16), .Z(\ab[19][13] ) );
  NR2 U921 ( .A(n152), .B(n16), .Z(\ab[19][12] ) );
  NR2 U922 ( .A(n153), .B(n16), .Z(\ab[19][11] ) );
  NR2 U923 ( .A(n154), .B(n16), .Z(\ab[19][10] ) );
  NR2 U924 ( .A(n164), .B(n16), .Z(\ab[19][0] ) );
  NR2 U925 ( .A(n155), .B(n21), .Z(\ab[18][9] ) );
  NR2 U926 ( .A(n156), .B(n21), .Z(\ab[18][8] ) );
  NR2 U927 ( .A(n157), .B(n21), .Z(\ab[18][7] ) );
  NR2 U928 ( .A(n158), .B(n21), .Z(\ab[18][6] ) );
  NR2 U929 ( .A(n159), .B(n21), .Z(\ab[18][5] ) );
  NR2 U930 ( .A(n160), .B(n21), .Z(\ab[18][4] ) );
  NR2 U931 ( .A(n108), .B(n21), .Z(\ab[18][47] ) );
  NR2 U932 ( .A(n107), .B(n21), .Z(\ab[18][46] ) );
  NR2 U933 ( .A(n106), .B(n21), .Z(\ab[18][45] ) );
  NR2 U934 ( .A(n105), .B(n21), .Z(\ab[18][44] ) );
  NR2 U935 ( .A(n104), .B(n21), .Z(\ab[18][43] ) );
  NR2 U936 ( .A(n103), .B(n21), .Z(\ab[18][42] ) );
  NR2 U937 ( .A(n102), .B(n20), .Z(\ab[18][41] ) );
  NR2 U938 ( .A(n101), .B(n20), .Z(\ab[18][40] ) );
  NR2 U939 ( .A(n161), .B(n20), .Z(\ab[18][3] ) );
  NR2 U940 ( .A(n125), .B(n20), .Z(\ab[18][39] ) );
  NR2 U941 ( .A(n126), .B(n20), .Z(\ab[18][38] ) );
  NR2 U942 ( .A(n127), .B(n20), .Z(\ab[18][37] ) );
  NR2 U943 ( .A(n128), .B(n20), .Z(\ab[18][36] ) );
  NR2 U944 ( .A(n129), .B(n20), .Z(\ab[18][35] ) );
  NR2 U945 ( .A(n130), .B(n20), .Z(\ab[18][34] ) );
  NR2 U946 ( .A(n131), .B(n20), .Z(\ab[18][33] ) );
  NR2 U947 ( .A(n132), .B(n20), .Z(\ab[18][32] ) );
  NR2 U948 ( .A(n133), .B(n20), .Z(\ab[18][31] ) );
  NR2 U949 ( .A(n134), .B(n21), .Z(\ab[18][30] ) );
  NR2 U950 ( .A(n162), .B(n20), .Z(\ab[18][2] ) );
  NR2 U951 ( .A(n135), .B(n20), .Z(\ab[18][29] ) );
  NR2 U952 ( .A(n136), .B(n21), .Z(\ab[18][28] ) );
  NR2 U953 ( .A(n137), .B(n21), .Z(\ab[18][27] ) );
  NR2 U954 ( .A(n138), .B(n21), .Z(\ab[18][26] ) );
  NR2 U955 ( .A(n139), .B(n21), .Z(\ab[18][25] ) );
  NR2 U956 ( .A(n140), .B(n21), .Z(\ab[18][24] ) );
  NR2 U957 ( .A(n141), .B(n21), .Z(\ab[18][23] ) );
  NR2 U958 ( .A(n142), .B(n21), .Z(\ab[18][22] ) );
  NR2 U959 ( .A(n143), .B(n21), .Z(\ab[18][21] ) );
  NR2 U960 ( .A(n144), .B(n21), .Z(\ab[18][20] ) );
  NR2 U961 ( .A(n163), .B(n20), .Z(\ab[18][1] ) );
  NR2 U962 ( .A(n145), .B(n21), .Z(\ab[18][19] ) );
  NR2 U963 ( .A(n146), .B(n21), .Z(\ab[18][18] ) );
  NR2 U964 ( .A(n147), .B(n21), .Z(\ab[18][17] ) );
  NR2 U965 ( .A(n148), .B(n21), .Z(\ab[18][16] ) );
  NR2 U966 ( .A(n149), .B(n21), .Z(\ab[18][15] ) );
  NR2 U967 ( .A(n150), .B(n21), .Z(\ab[18][14] ) );
  NR2 U968 ( .A(n151), .B(n21), .Z(\ab[18][13] ) );
  NR2 U969 ( .A(n152), .B(n21), .Z(\ab[18][12] ) );
  NR2 U970 ( .A(n153), .B(n21), .Z(\ab[18][11] ) );
  NR2 U971 ( .A(n154), .B(n21), .Z(\ab[18][10] ) );
  NR2 U972 ( .A(n164), .B(n21), .Z(\ab[18][0] ) );
  NR2 U973 ( .A(n155), .B(n22), .Z(\ab[17][9] ) );
  NR2 U974 ( .A(n156), .B(n22), .Z(\ab[17][8] ) );
  NR2 U975 ( .A(n157), .B(n22), .Z(\ab[17][7] ) );
  NR2 U976 ( .A(n158), .B(n22), .Z(\ab[17][6] ) );
  NR2 U977 ( .A(n159), .B(n22), .Z(\ab[17][5] ) );
  NR2 U978 ( .A(n160), .B(n22), .Z(\ab[17][4] ) );
  NR2 U979 ( .A(n108), .B(n22), .Z(\ab[17][47] ) );
  NR2 U980 ( .A(n107), .B(n22), .Z(\ab[17][46] ) );
  NR2 U981 ( .A(n106), .B(n22), .Z(\ab[17][45] ) );
  NR2 U982 ( .A(n105), .B(n22), .Z(\ab[17][44] ) );
  NR2 U983 ( .A(n104), .B(n22), .Z(\ab[17][43] ) );
  NR2 U984 ( .A(n103), .B(n22), .Z(\ab[17][42] ) );
  NR2 U985 ( .A(n102), .B(n22), .Z(\ab[17][41] ) );
  NR2 U986 ( .A(n101), .B(n22), .Z(\ab[17][40] ) );
  NR2 U987 ( .A(n161), .B(n22), .Z(\ab[17][3] ) );
  NR2 U988 ( .A(n125), .B(n22), .Z(\ab[17][39] ) );
  NR2 U989 ( .A(n126), .B(n22), .Z(\ab[17][38] ) );
  NR2 U990 ( .A(n127), .B(n22), .Z(\ab[17][37] ) );
  NR2 U991 ( .A(n128), .B(n22), .Z(\ab[17][36] ) );
  NR2 U992 ( .A(n129), .B(n22), .Z(\ab[17][35] ) );
  NR2 U993 ( .A(n130), .B(n22), .Z(\ab[17][34] ) );
  NR2 U994 ( .A(n131), .B(n22), .Z(\ab[17][33] ) );
  NR2 U995 ( .A(n132), .B(n22), .Z(\ab[17][32] ) );
  NR2 U996 ( .A(n133), .B(n22), .Z(\ab[17][31] ) );
  NR2 U997 ( .A(n134), .B(n22), .Z(\ab[17][30] ) );
  NR2 U998 ( .A(n162), .B(n22), .Z(\ab[17][2] ) );
  NR2 U999 ( .A(n135), .B(n22), .Z(\ab[17][29] ) );
  NR2 U1000 ( .A(n136), .B(n22), .Z(\ab[17][28] ) );
  NR2 U1001 ( .A(n137), .B(n22), .Z(\ab[17][27] ) );
  NR2 U1002 ( .A(n138), .B(n22), .Z(\ab[17][26] ) );
  NR2 U1003 ( .A(n139), .B(n22), .Z(\ab[17][25] ) );
  NR2 U1004 ( .A(n140), .B(n22), .Z(\ab[17][24] ) );
  NR2 U1005 ( .A(n141), .B(n22), .Z(\ab[17][23] ) );
  NR2 U1006 ( .A(n142), .B(n22), .Z(\ab[17][22] ) );
  NR2 U1007 ( .A(n143), .B(n22), .Z(\ab[17][21] ) );
  NR2 U1008 ( .A(n144), .B(n22), .Z(\ab[17][20] ) );
  NR2 U1009 ( .A(n163), .B(n22), .Z(\ab[17][1] ) );
  NR2 U1010 ( .A(n145), .B(n22), .Z(\ab[17][19] ) );
  NR2 U1011 ( .A(n146), .B(n22), .Z(\ab[17][18] ) );
  NR2 U1012 ( .A(n147), .B(n22), .Z(\ab[17][17] ) );
  NR2 U1013 ( .A(n148), .B(n22), .Z(\ab[17][16] ) );
  NR2 U1014 ( .A(n149), .B(n22), .Z(\ab[17][15] ) );
  NR2 U1015 ( .A(n150), .B(n22), .Z(\ab[17][14] ) );
  NR2 U1016 ( .A(n151), .B(n22), .Z(\ab[17][13] ) );
  NR2 U1017 ( .A(n152), .B(n22), .Z(\ab[17][12] ) );
  NR2 U1018 ( .A(n153), .B(n22), .Z(\ab[17][11] ) );
  NR2 U1019 ( .A(n154), .B(n22), .Z(\ab[17][10] ) );
  NR2 U1020 ( .A(n164), .B(n22), .Z(\ab[17][0] ) );
  NR2 U1021 ( .A(n155), .B(n25), .Z(\ab[16][9] ) );
  NR2 U1022 ( .A(n156), .B(n25), .Z(\ab[16][8] ) );
  NR2 U1023 ( .A(n157), .B(n25), .Z(\ab[16][7] ) );
  NR2 U1024 ( .A(n158), .B(n25), .Z(\ab[16][6] ) );
  NR2 U1025 ( .A(n159), .B(n25), .Z(\ab[16][5] ) );
  NR2 U1026 ( .A(n160), .B(n25), .Z(\ab[16][4] ) );
  NR2 U1027 ( .A(n108), .B(n25), .Z(\ab[16][47] ) );
  NR2 U1028 ( .A(n107), .B(n25), .Z(\ab[16][46] ) );
  NR2 U1029 ( .A(n106), .B(n25), .Z(\ab[16][45] ) );
  NR2 U1030 ( .A(n105), .B(n25), .Z(\ab[16][44] ) );
  NR2 U1031 ( .A(n104), .B(n25), .Z(\ab[16][43] ) );
  NR2 U1032 ( .A(n103), .B(n25), .Z(\ab[16][42] ) );
  NR2 U1033 ( .A(n102), .B(n24), .Z(\ab[16][41] ) );
  NR2 U1034 ( .A(n101), .B(n24), .Z(\ab[16][40] ) );
  NR2 U1035 ( .A(n161), .B(n24), .Z(\ab[16][3] ) );
  NR2 U1036 ( .A(n125), .B(n24), .Z(\ab[16][39] ) );
  NR2 U1037 ( .A(n126), .B(n24), .Z(\ab[16][38] ) );
  NR2 U1038 ( .A(n127), .B(n24), .Z(\ab[16][37] ) );
  NR2 U1039 ( .A(n128), .B(n24), .Z(\ab[16][36] ) );
  NR2 U1040 ( .A(n129), .B(n24), .Z(\ab[16][35] ) );
  NR2 U1041 ( .A(n130), .B(n24), .Z(\ab[16][34] ) );
  NR2 U1042 ( .A(n131), .B(n24), .Z(\ab[16][33] ) );
  NR2 U1043 ( .A(n132), .B(n24), .Z(\ab[16][32] ) );
  NR2 U1044 ( .A(n133), .B(n24), .Z(\ab[16][31] ) );
  NR2 U1045 ( .A(n134), .B(n25), .Z(\ab[16][30] ) );
  NR2 U1046 ( .A(n162), .B(n23), .Z(\ab[16][2] ) );
  NR2 U1047 ( .A(n135), .B(n25), .Z(\ab[16][29] ) );
  NR2 U1048 ( .A(n136), .B(n25), .Z(\ab[16][28] ) );
  NR2 U1049 ( .A(n137), .B(n25), .Z(\ab[16][27] ) );
  NR2 U1050 ( .A(n138), .B(n25), .Z(\ab[16][26] ) );
  NR2 U1051 ( .A(n139), .B(n25), .Z(\ab[16][25] ) );
  NR2 U1052 ( .A(n140), .B(n25), .Z(\ab[16][24] ) );
  NR2 U1053 ( .A(n141), .B(n25), .Z(\ab[16][23] ) );
  NR2 U1054 ( .A(n142), .B(n25), .Z(\ab[16][22] ) );
  NR2 U1055 ( .A(n143), .B(n25), .Z(\ab[16][21] ) );
  NR2 U1056 ( .A(n144), .B(n25), .Z(\ab[16][20] ) );
  NR2 U1057 ( .A(n163), .B(n23), .Z(\ab[16][1] ) );
  NR2 U1058 ( .A(n145), .B(n23), .Z(\ab[16][19] ) );
  NR2 U1059 ( .A(n146), .B(n23), .Z(\ab[16][18] ) );
  NR2 U1060 ( .A(n147), .B(n23), .Z(\ab[16][17] ) );
  NR2 U1061 ( .A(n148), .B(n23), .Z(\ab[16][16] ) );
  NR2 U1062 ( .A(n149), .B(n23), .Z(\ab[16][15] ) );
  NR2 U1063 ( .A(n150), .B(n23), .Z(\ab[16][14] ) );
  NR2 U1064 ( .A(n151), .B(n23), .Z(\ab[16][13] ) );
  NR2 U1065 ( .A(n152), .B(n23), .Z(\ab[16][12] ) );
  NR2 U1066 ( .A(n153), .B(n23), .Z(\ab[16][11] ) );
  NR2 U1067 ( .A(n154), .B(n23), .Z(\ab[16][10] ) );
  NR2 U1068 ( .A(n164), .B(n23), .Z(\ab[16][0] ) );
  NR2 U1069 ( .A(n155), .B(n29), .Z(\ab[15][9] ) );
  NR2 U1070 ( .A(n156), .B(n29), .Z(\ab[15][8] ) );
  NR2 U1071 ( .A(n157), .B(n29), .Z(\ab[15][7] ) );
  NR2 U1072 ( .A(n158), .B(n29), .Z(\ab[15][6] ) );
  NR2 U1073 ( .A(n159), .B(n29), .Z(\ab[15][5] ) );
  NR2 U1074 ( .A(n160), .B(n29), .Z(\ab[15][4] ) );
  NR2 U1075 ( .A(n108), .B(n29), .Z(\ab[15][47] ) );
  NR2 U1076 ( .A(n107), .B(n29), .Z(\ab[15][46] ) );
  NR2 U1077 ( .A(n106), .B(n29), .Z(\ab[15][45] ) );
  NR2 U1078 ( .A(n105), .B(n29), .Z(\ab[15][44] ) );
  NR2 U1079 ( .A(n104), .B(n29), .Z(\ab[15][43] ) );
  NR2 U1080 ( .A(n103), .B(n29), .Z(\ab[15][42] ) );
  NR2 U1081 ( .A(n102), .B(n28), .Z(\ab[15][41] ) );
  NR2 U1082 ( .A(n101), .B(n28), .Z(\ab[15][40] ) );
  NR2 U1083 ( .A(n161), .B(n28), .Z(\ab[15][3] ) );
  NR2 U1084 ( .A(n125), .B(n28), .Z(\ab[15][39] ) );
  NR2 U1085 ( .A(n126), .B(n28), .Z(\ab[15][38] ) );
  NR2 U1086 ( .A(n127), .B(n28), .Z(\ab[15][37] ) );
  NR2 U1087 ( .A(n128), .B(n28), .Z(\ab[15][36] ) );
  NR2 U1088 ( .A(n129), .B(n28), .Z(\ab[15][35] ) );
  NR2 U1089 ( .A(n130), .B(n28), .Z(\ab[15][34] ) );
  NR2 U1090 ( .A(n131), .B(n28), .Z(\ab[15][33] ) );
  NR2 U1091 ( .A(n132), .B(n28), .Z(\ab[15][32] ) );
  NR2 U1092 ( .A(n133), .B(n28), .Z(\ab[15][31] ) );
  NR2 U1093 ( .A(n134), .B(n27), .Z(\ab[15][30] ) );
  NR2 U1094 ( .A(n162), .B(n27), .Z(\ab[15][2] ) );
  NR2 U1095 ( .A(n135), .B(n27), .Z(\ab[15][29] ) );
  NR2 U1096 ( .A(n136), .B(n27), .Z(\ab[15][28] ) );
  NR2 U1097 ( .A(n137), .B(n27), .Z(\ab[15][27] ) );
  NR2 U1098 ( .A(n138), .B(n27), .Z(\ab[15][26] ) );
  NR2 U1099 ( .A(n139), .B(n27), .Z(\ab[15][25] ) );
  NR2 U1100 ( .A(n140), .B(n27), .Z(\ab[15][24] ) );
  NR2 U1101 ( .A(n141), .B(n27), .Z(\ab[15][23] ) );
  NR2 U1102 ( .A(n142), .B(n27), .Z(\ab[15][22] ) );
  NR2 U1103 ( .A(n143), .B(n27), .Z(\ab[15][21] ) );
  NR2 U1104 ( .A(n144), .B(n27), .Z(\ab[15][20] ) );
  NR2 U1105 ( .A(n163), .B(n26), .Z(\ab[15][1] ) );
  NR2 U1106 ( .A(n145), .B(n26), .Z(\ab[15][19] ) );
  NR2 U1107 ( .A(n146), .B(n26), .Z(\ab[15][18] ) );
  NR2 U1108 ( .A(n147), .B(n26), .Z(\ab[15][17] ) );
  NR2 U1109 ( .A(n148), .B(n26), .Z(\ab[15][16] ) );
  NR2 U1110 ( .A(n149), .B(n26), .Z(\ab[15][15] ) );
  NR2 U1111 ( .A(n150), .B(n26), .Z(\ab[15][14] ) );
  NR2 U1112 ( .A(n151), .B(n26), .Z(\ab[15][13] ) );
  NR2 U1113 ( .A(n152), .B(n26), .Z(\ab[15][12] ) );
  NR2 U1114 ( .A(n153), .B(n26), .Z(\ab[15][11] ) );
  NR2 U1115 ( .A(n154), .B(n26), .Z(\ab[15][10] ) );
  NR2 U1116 ( .A(n164), .B(n26), .Z(\ab[15][0] ) );
  NR2 U1117 ( .A(n155), .B(n6), .Z(\ab[14][9] ) );
  NR2 U1118 ( .A(n156), .B(n6), .Z(\ab[14][8] ) );
  NR2 U1119 ( .A(n157), .B(n6), .Z(\ab[14][7] ) );
  NR2 U1120 ( .A(n158), .B(n6), .Z(\ab[14][6] ) );
  NR2 U1121 ( .A(n159), .B(n6), .Z(\ab[14][5] ) );
  NR2 U1122 ( .A(n160), .B(n6), .Z(\ab[14][4] ) );
  NR2 U1123 ( .A(n108), .B(n6), .Z(\ab[14][47] ) );
  NR2 U1124 ( .A(n107), .B(n6), .Z(\ab[14][46] ) );
  NR2 U1125 ( .A(n106), .B(n6), .Z(\ab[14][45] ) );
  NR2 U1126 ( .A(n105), .B(n6), .Z(\ab[14][44] ) );
  NR2 U1127 ( .A(n104), .B(n6), .Z(\ab[14][43] ) );
  NR2 U1128 ( .A(n103), .B(n6), .Z(\ab[14][42] ) );
  NR2 U1129 ( .A(n102), .B(n5), .Z(\ab[14][41] ) );
  NR2 U1130 ( .A(n101), .B(n5), .Z(\ab[14][40] ) );
  NR2 U1131 ( .A(n161), .B(n5), .Z(\ab[14][3] ) );
  NR2 U1132 ( .A(n125), .B(n5), .Z(\ab[14][39] ) );
  NR2 U1133 ( .A(n126), .B(n5), .Z(\ab[14][38] ) );
  NR2 U1134 ( .A(n127), .B(n5), .Z(\ab[14][37] ) );
  NR2 U1135 ( .A(n128), .B(n5), .Z(\ab[14][36] ) );
  NR2 U1136 ( .A(n129), .B(n5), .Z(\ab[14][35] ) );
  NR2 U1137 ( .A(n130), .B(n5), .Z(\ab[14][34] ) );
  NR2 U1138 ( .A(n131), .B(n5), .Z(\ab[14][33] ) );
  NR2 U1139 ( .A(n132), .B(n5), .Z(\ab[14][32] ) );
  NR2 U1140 ( .A(n133), .B(n5), .Z(\ab[14][31] ) );
  NR2 U1141 ( .A(n134), .B(n4), .Z(\ab[14][30] ) );
  NR2 U1142 ( .A(n162), .B(n4), .Z(\ab[14][2] ) );
  NR2 U1143 ( .A(n135), .B(n4), .Z(\ab[14][29] ) );
  NR2 U1144 ( .A(n136), .B(n4), .Z(\ab[14][28] ) );
  NR2 U1145 ( .A(n137), .B(n4), .Z(\ab[14][27] ) );
  NR2 U1146 ( .A(n138), .B(n4), .Z(\ab[14][26] ) );
  NR2 U1147 ( .A(n139), .B(n4), .Z(\ab[14][25] ) );
  NR2 U1148 ( .A(n140), .B(n4), .Z(\ab[14][24] ) );
  NR2 U1149 ( .A(n141), .B(n4), .Z(\ab[14][23] ) );
  NR2 U1150 ( .A(n142), .B(n4), .Z(\ab[14][22] ) );
  NR2 U1151 ( .A(n143), .B(n4), .Z(\ab[14][21] ) );
  NR2 U1152 ( .A(n144), .B(n4), .Z(\ab[14][20] ) );
  NR2 U1153 ( .A(n163), .B(n3), .Z(\ab[14][1] ) );
  NR2 U1154 ( .A(n145), .B(n3), .Z(\ab[14][19] ) );
  NR2 U1155 ( .A(n146), .B(n3), .Z(\ab[14][18] ) );
  NR2 U1156 ( .A(n147), .B(n3), .Z(\ab[14][17] ) );
  NR2 U1157 ( .A(n148), .B(n3), .Z(\ab[14][16] ) );
  NR2 U1158 ( .A(n149), .B(n3), .Z(\ab[14][15] ) );
  NR2 U1159 ( .A(n150), .B(n3), .Z(\ab[14][14] ) );
  NR2 U1160 ( .A(n151), .B(n3), .Z(\ab[14][13] ) );
  NR2 U1161 ( .A(n152), .B(n3), .Z(\ab[14][12] ) );
  NR2 U1162 ( .A(n153), .B(n3), .Z(\ab[14][11] ) );
  NR2 U1163 ( .A(n154), .B(n3), .Z(\ab[14][10] ) );
  NR2 U1164 ( .A(n164), .B(n3), .Z(\ab[14][0] ) );
  NR2 U1165 ( .A(n155), .B(n34), .Z(\ab[13][9] ) );
  NR2 U1166 ( .A(n156), .B(n34), .Z(\ab[13][8] ) );
  NR2 U1167 ( .A(n157), .B(n34), .Z(\ab[13][7] ) );
  NR2 U1168 ( .A(n158), .B(n34), .Z(\ab[13][6] ) );
  NR2 U1169 ( .A(n159), .B(n34), .Z(\ab[13][5] ) );
  NR2 U1170 ( .A(n160), .B(n34), .Z(\ab[13][4] ) );
  NR2 U1171 ( .A(n108), .B(n34), .Z(\ab[13][47] ) );
  NR2 U1172 ( .A(n107), .B(n34), .Z(\ab[13][46] ) );
  NR2 U1173 ( .A(n106), .B(n34), .Z(\ab[13][45] ) );
  NR2 U1174 ( .A(n105), .B(n34), .Z(\ab[13][44] ) );
  NR2 U1175 ( .A(n104), .B(n34), .Z(\ab[13][43] ) );
  NR2 U1176 ( .A(n103), .B(n34), .Z(\ab[13][42] ) );
  NR2 U1177 ( .A(n102), .B(n33), .Z(\ab[13][41] ) );
  NR2 U1178 ( .A(n101), .B(n33), .Z(\ab[13][40] ) );
  NR2 U1179 ( .A(n161), .B(n33), .Z(\ab[13][3] ) );
  NR2 U1180 ( .A(n125), .B(n33), .Z(\ab[13][39] ) );
  NR2 U1181 ( .A(n126), .B(n33), .Z(\ab[13][38] ) );
  NR2 U1182 ( .A(n127), .B(n33), .Z(\ab[13][37] ) );
  NR2 U1183 ( .A(n128), .B(n33), .Z(\ab[13][36] ) );
  NR2 U1184 ( .A(n129), .B(n33), .Z(\ab[13][35] ) );
  NR2 U1185 ( .A(n130), .B(n33), .Z(\ab[13][34] ) );
  NR2 U1186 ( .A(n131), .B(n33), .Z(\ab[13][33] ) );
  NR2 U1187 ( .A(n132), .B(n33), .Z(\ab[13][32] ) );
  NR2 U1188 ( .A(n133), .B(n33), .Z(\ab[13][31] ) );
  NR2 U1189 ( .A(n134), .B(n32), .Z(\ab[13][30] ) );
  NR2 U1190 ( .A(n162), .B(n32), .Z(\ab[13][2] ) );
  NR2 U1191 ( .A(n135), .B(n32), .Z(\ab[13][29] ) );
  NR2 U1192 ( .A(n136), .B(n32), .Z(\ab[13][28] ) );
  NR2 U1193 ( .A(n137), .B(n32), .Z(\ab[13][27] ) );
  NR2 U1194 ( .A(n138), .B(n32), .Z(\ab[13][26] ) );
  NR2 U1195 ( .A(n139), .B(n32), .Z(\ab[13][25] ) );
  NR2 U1196 ( .A(n140), .B(n32), .Z(\ab[13][24] ) );
  NR2 U1197 ( .A(n141), .B(n32), .Z(\ab[13][23] ) );
  NR2 U1198 ( .A(n142), .B(n32), .Z(\ab[13][22] ) );
  NR2 U1199 ( .A(n143), .B(n32), .Z(\ab[13][21] ) );
  NR2 U1200 ( .A(n144), .B(n32), .Z(\ab[13][20] ) );
  NR2 U1201 ( .A(n163), .B(n31), .Z(\ab[13][1] ) );
  NR2 U1202 ( .A(n145), .B(n31), .Z(\ab[13][19] ) );
  NR2 U1203 ( .A(n146), .B(n31), .Z(\ab[13][18] ) );
  NR2 U1204 ( .A(n147), .B(n31), .Z(\ab[13][17] ) );
  NR2 U1205 ( .A(n148), .B(n31), .Z(\ab[13][16] ) );
  NR2 U1206 ( .A(n149), .B(n31), .Z(\ab[13][15] ) );
  NR2 U1207 ( .A(n150), .B(n31), .Z(\ab[13][14] ) );
  NR2 U1208 ( .A(n151), .B(n31), .Z(\ab[13][13] ) );
  NR2 U1209 ( .A(n152), .B(n31), .Z(\ab[13][12] ) );
  NR2 U1210 ( .A(n153), .B(n31), .Z(\ab[13][11] ) );
  NR2 U1211 ( .A(n154), .B(n31), .Z(\ab[13][10] ) );
  NR2 U1212 ( .A(n164), .B(n31), .Z(\ab[13][0] ) );
  NR2 U1213 ( .A(n155), .B(n99), .Z(\ab[12][9] ) );
  NR2 U1214 ( .A(n156), .B(n99), .Z(\ab[12][8] ) );
  NR2 U1215 ( .A(n157), .B(n99), .Z(\ab[12][7] ) );
  NR2 U1216 ( .A(n158), .B(n99), .Z(\ab[12][6] ) );
  NR2 U1217 ( .A(n159), .B(n99), .Z(\ab[12][5] ) );
  NR2 U1218 ( .A(n160), .B(n99), .Z(\ab[12][4] ) );
  NR2 U1219 ( .A(n108), .B(n99), .Z(\ab[12][47] ) );
  NR2 U1220 ( .A(n107), .B(n99), .Z(\ab[12][46] ) );
  NR2 U1221 ( .A(n106), .B(n99), .Z(\ab[12][45] ) );
  NR2 U1222 ( .A(n105), .B(n99), .Z(\ab[12][44] ) );
  NR2 U1223 ( .A(n104), .B(n99), .Z(\ab[12][43] ) );
  NR2 U1224 ( .A(n103), .B(n99), .Z(\ab[12][42] ) );
  NR2 U1225 ( .A(n102), .B(n98), .Z(\ab[12][41] ) );
  NR2 U1226 ( .A(n101), .B(n98), .Z(\ab[12][40] ) );
  NR2 U1227 ( .A(n161), .B(n98), .Z(\ab[12][3] ) );
  NR2 U1228 ( .A(n125), .B(n98), .Z(\ab[12][39] ) );
  NR2 U1229 ( .A(n126), .B(n98), .Z(\ab[12][38] ) );
  NR2 U1230 ( .A(n127), .B(n98), .Z(\ab[12][37] ) );
  NR2 U1231 ( .A(n128), .B(n98), .Z(\ab[12][36] ) );
  NR2 U1232 ( .A(n129), .B(n98), .Z(\ab[12][35] ) );
  NR2 U1233 ( .A(n130), .B(n98), .Z(\ab[12][34] ) );
  NR2 U1234 ( .A(n131), .B(n98), .Z(\ab[12][33] ) );
  NR2 U1235 ( .A(n132), .B(n98), .Z(\ab[12][32] ) );
  NR2 U1236 ( .A(n133), .B(n98), .Z(\ab[12][31] ) );
  NR2 U1237 ( .A(n134), .B(n97), .Z(\ab[12][30] ) );
  NR2 U1238 ( .A(n162), .B(n97), .Z(\ab[12][2] ) );
  NR2 U1239 ( .A(n135), .B(n97), .Z(\ab[12][29] ) );
  NR2 U1240 ( .A(n136), .B(n97), .Z(\ab[12][28] ) );
  NR2 U1241 ( .A(n137), .B(n97), .Z(\ab[12][27] ) );
  NR2 U1242 ( .A(n138), .B(n97), .Z(\ab[12][26] ) );
  NR2 U1243 ( .A(n139), .B(n97), .Z(\ab[12][25] ) );
  NR2 U1244 ( .A(n140), .B(n97), .Z(\ab[12][24] ) );
  NR2 U1245 ( .A(n141), .B(n97), .Z(\ab[12][23] ) );
  NR2 U1246 ( .A(n142), .B(n97), .Z(\ab[12][22] ) );
  NR2 U1247 ( .A(n143), .B(n97), .Z(\ab[12][21] ) );
  NR2 U1248 ( .A(n144), .B(n97), .Z(\ab[12][20] ) );
  NR2 U1249 ( .A(n163), .B(n96), .Z(\ab[12][1] ) );
  NR2 U1250 ( .A(n145), .B(n96), .Z(\ab[12][19] ) );
  NR2 U1251 ( .A(n146), .B(n96), .Z(\ab[12][18] ) );
  NR2 U1252 ( .A(n147), .B(n96), .Z(\ab[12][17] ) );
  NR2 U1253 ( .A(n148), .B(n96), .Z(\ab[12][16] ) );
  NR2 U1254 ( .A(n149), .B(n96), .Z(\ab[12][15] ) );
  NR2 U1255 ( .A(n150), .B(n96), .Z(\ab[12][14] ) );
  NR2 U1256 ( .A(n151), .B(n96), .Z(\ab[12][13] ) );
  NR2 U1257 ( .A(n152), .B(n96), .Z(\ab[12][12] ) );
  NR2 U1258 ( .A(n153), .B(n96), .Z(\ab[12][11] ) );
  NR2 U1259 ( .A(n154), .B(n96), .Z(\ab[12][10] ) );
  NR2 U1260 ( .A(n164), .B(n96), .Z(\ab[12][0] ) );
  NR2 U1261 ( .A(n155), .B(n94), .Z(\ab[11][9] ) );
  NR2 U1262 ( .A(n156), .B(n94), .Z(\ab[11][8] ) );
  NR2 U1263 ( .A(n157), .B(n94), .Z(\ab[11][7] ) );
  NR2 U1264 ( .A(n158), .B(n94), .Z(\ab[11][6] ) );
  NR2 U1265 ( .A(n159), .B(n94), .Z(\ab[11][5] ) );
  NR2 U1266 ( .A(n160), .B(n94), .Z(\ab[11][4] ) );
  NR2 U1267 ( .A(n108), .B(n94), .Z(\ab[11][47] ) );
  NR2 U1268 ( .A(n107), .B(n94), .Z(\ab[11][46] ) );
  NR2 U1269 ( .A(n106), .B(n94), .Z(\ab[11][45] ) );
  NR2 U1270 ( .A(n105), .B(n94), .Z(\ab[11][44] ) );
  NR2 U1271 ( .A(n104), .B(n94), .Z(\ab[11][43] ) );
  NR2 U1272 ( .A(n103), .B(n94), .Z(\ab[11][42] ) );
  NR2 U1273 ( .A(n102), .B(n93), .Z(\ab[11][41] ) );
  NR2 U1274 ( .A(n101), .B(n93), .Z(\ab[11][40] ) );
  NR2 U1275 ( .A(n161), .B(n93), .Z(\ab[11][3] ) );
  NR2 U1276 ( .A(n125), .B(n93), .Z(\ab[11][39] ) );
  NR2 U1277 ( .A(n126), .B(n93), .Z(\ab[11][38] ) );
  NR2 U1278 ( .A(n127), .B(n93), .Z(\ab[11][37] ) );
  NR2 U1279 ( .A(n128), .B(n93), .Z(\ab[11][36] ) );
  NR2 U1280 ( .A(n129), .B(n93), .Z(\ab[11][35] ) );
  NR2 U1281 ( .A(n130), .B(n93), .Z(\ab[11][34] ) );
  NR2 U1282 ( .A(n131), .B(n93), .Z(\ab[11][33] ) );
  NR2 U1283 ( .A(n132), .B(n93), .Z(\ab[11][32] ) );
  NR2 U1284 ( .A(n133), .B(n93), .Z(\ab[11][31] ) );
  NR2 U1285 ( .A(n134), .B(n92), .Z(\ab[11][30] ) );
  NR2 U1286 ( .A(n162), .B(n92), .Z(\ab[11][2] ) );
  NR2 U1287 ( .A(n135), .B(n92), .Z(\ab[11][29] ) );
  NR2 U1288 ( .A(n136), .B(n92), .Z(\ab[11][28] ) );
  NR2 U1289 ( .A(n137), .B(n92), .Z(\ab[11][27] ) );
  NR2 U1290 ( .A(n138), .B(n92), .Z(\ab[11][26] ) );
  NR2 U1291 ( .A(n139), .B(n92), .Z(\ab[11][25] ) );
  NR2 U1292 ( .A(n140), .B(n92), .Z(\ab[11][24] ) );
  NR2 U1293 ( .A(n141), .B(n92), .Z(\ab[11][23] ) );
  NR2 U1294 ( .A(n142), .B(n92), .Z(\ab[11][22] ) );
  NR2 U1295 ( .A(n143), .B(n92), .Z(\ab[11][21] ) );
  NR2 U1296 ( .A(n144), .B(n92), .Z(\ab[11][20] ) );
  NR2 U1297 ( .A(n163), .B(n91), .Z(\ab[11][1] ) );
  NR2 U1298 ( .A(n145), .B(n91), .Z(\ab[11][19] ) );
  NR2 U1299 ( .A(n146), .B(n91), .Z(\ab[11][18] ) );
  NR2 U1300 ( .A(n147), .B(n91), .Z(\ab[11][17] ) );
  NR2 U1301 ( .A(n148), .B(n91), .Z(\ab[11][16] ) );
  NR2 U1302 ( .A(n149), .B(n91), .Z(\ab[11][15] ) );
  NR2 U1303 ( .A(n150), .B(n91), .Z(\ab[11][14] ) );
  NR2 U1304 ( .A(n151), .B(n91), .Z(\ab[11][13] ) );
  NR2 U1305 ( .A(n152), .B(n91), .Z(\ab[11][12] ) );
  NR2 U1306 ( .A(n153), .B(n91), .Z(\ab[11][11] ) );
  NR2 U1307 ( .A(n154), .B(n91), .Z(\ab[11][10] ) );
  NR2 U1308 ( .A(n164), .B(n91), .Z(\ab[11][0] ) );
  NR2 U1309 ( .A(n155), .B(n89), .Z(\ab[10][9] ) );
  NR2 U1310 ( .A(n156), .B(n89), .Z(\ab[10][8] ) );
  NR2 U1311 ( .A(n157), .B(n89), .Z(\ab[10][7] ) );
  NR2 U1312 ( .A(n158), .B(n89), .Z(\ab[10][6] ) );
  NR2 U1313 ( .A(n159), .B(n89), .Z(\ab[10][5] ) );
  NR2 U1314 ( .A(n160), .B(n89), .Z(\ab[10][4] ) );
  NR2 U1315 ( .A(n108), .B(n89), .Z(\ab[10][47] ) );
  NR2 U1316 ( .A(n107), .B(n89), .Z(\ab[10][46] ) );
  NR2 U1317 ( .A(n106), .B(n89), .Z(\ab[10][45] ) );
  NR2 U1318 ( .A(n105), .B(n89), .Z(\ab[10][44] ) );
  NR2 U1319 ( .A(n104), .B(n89), .Z(\ab[10][43] ) );
  NR2 U1320 ( .A(n103), .B(n89), .Z(\ab[10][42] ) );
  NR2 U1321 ( .A(n102), .B(n88), .Z(\ab[10][41] ) );
  NR2 U1322 ( .A(n101), .B(n88), .Z(\ab[10][40] ) );
  NR2 U1323 ( .A(n161), .B(n88), .Z(\ab[10][3] ) );
  NR2 U1324 ( .A(n125), .B(n88), .Z(\ab[10][39] ) );
  NR2 U1325 ( .A(n126), .B(n88), .Z(\ab[10][38] ) );
  NR2 U1326 ( .A(n127), .B(n88), .Z(\ab[10][37] ) );
  NR2 U1327 ( .A(n128), .B(n88), .Z(\ab[10][36] ) );
  NR2 U1328 ( .A(n129), .B(n88), .Z(\ab[10][35] ) );
  NR2 U1329 ( .A(n130), .B(n88), .Z(\ab[10][34] ) );
  NR2 U1330 ( .A(n131), .B(n88), .Z(\ab[10][33] ) );
  NR2 U1331 ( .A(n132), .B(n88), .Z(\ab[10][32] ) );
  NR2 U1332 ( .A(n133), .B(n88), .Z(\ab[10][31] ) );
  NR2 U1333 ( .A(n134), .B(n87), .Z(\ab[10][30] ) );
  NR2 U1334 ( .A(n162), .B(n87), .Z(\ab[10][2] ) );
  NR2 U1335 ( .A(n135), .B(n87), .Z(\ab[10][29] ) );
  NR2 U1336 ( .A(n136), .B(n87), .Z(\ab[10][28] ) );
  NR2 U1337 ( .A(n137), .B(n87), .Z(\ab[10][27] ) );
  NR2 U1338 ( .A(n138), .B(n87), .Z(\ab[10][26] ) );
  NR2 U1339 ( .A(n139), .B(n87), .Z(\ab[10][25] ) );
  NR2 U1340 ( .A(n140), .B(n87), .Z(\ab[10][24] ) );
  NR2 U1341 ( .A(n141), .B(n87), .Z(\ab[10][23] ) );
  NR2 U1342 ( .A(n142), .B(n87), .Z(\ab[10][22] ) );
  NR2 U1343 ( .A(n143), .B(n87), .Z(\ab[10][21] ) );
  NR2 U1344 ( .A(n144), .B(n87), .Z(\ab[10][20] ) );
  NR2 U1345 ( .A(n163), .B(n86), .Z(\ab[10][1] ) );
  NR2 U1346 ( .A(n145), .B(n86), .Z(\ab[10][19] ) );
  NR2 U1347 ( .A(n146), .B(n86), .Z(\ab[10][18] ) );
  NR2 U1348 ( .A(n147), .B(n86), .Z(\ab[10][17] ) );
  NR2 U1349 ( .A(n148), .B(n86), .Z(\ab[10][16] ) );
  NR2 U1350 ( .A(n149), .B(n86), .Z(\ab[10][15] ) );
  NR2 U1351 ( .A(n150), .B(n86), .Z(\ab[10][14] ) );
  NR2 U1352 ( .A(n151), .B(n86), .Z(\ab[10][13] ) );
  NR2 U1353 ( .A(n152), .B(n86), .Z(\ab[10][12] ) );
  NR2 U1354 ( .A(n153), .B(n86), .Z(\ab[10][11] ) );
  NR2 U1355 ( .A(n154), .B(n86), .Z(\ab[10][10] ) );
  NR2 U1356 ( .A(n164), .B(n86), .Z(\ab[10][0] ) );
  NR2 U1357 ( .A(n155), .B(n39), .Z(\ab[0][9] ) );
  NR2 U1358 ( .A(n156), .B(n39), .Z(\ab[0][8] ) );
  NR2 U1359 ( .A(n157), .B(n39), .Z(\ab[0][7] ) );
  NR2 U1360 ( .A(n158), .B(n39), .Z(\ab[0][6] ) );
  NR2 U1361 ( .A(n159), .B(n39), .Z(\ab[0][5] ) );
  NR2 U1362 ( .A(n160), .B(n39), .Z(\ab[0][4] ) );
  NR2 U1363 ( .A(n108), .B(n39), .Z(\ab[0][47] ) );
  NR2 U1364 ( .A(n107), .B(n39), .Z(\ab[0][46] ) );
  NR2 U1365 ( .A(n106), .B(n39), .Z(\ab[0][45] ) );
  NR2 U1366 ( .A(n105), .B(n39), .Z(\ab[0][44] ) );
  NR2 U1367 ( .A(n104), .B(n38), .Z(\ab[0][43] ) );
  NR2 U1368 ( .A(n103), .B(n38), .Z(\ab[0][42] ) );
  NR2 U1369 ( .A(n102), .B(n38), .Z(\ab[0][41] ) );
  NR2 U1370 ( .A(n101), .B(n38), .Z(\ab[0][40] ) );
  NR2 U1371 ( .A(n161), .B(n38), .Z(\ab[0][3] ) );
  NR2 U1372 ( .A(n125), .B(n38), .Z(\ab[0][39] ) );
  NR2 U1373 ( .A(n126), .B(n38), .Z(\ab[0][38] ) );
  NR2 U1374 ( .A(n127), .B(n38), .Z(\ab[0][37] ) );
  NR2 U1375 ( .A(n128), .B(n38), .Z(\ab[0][36] ) );
  NR2 U1376 ( .A(n129), .B(n38), .Z(\ab[0][35] ) );
  NR2 U1377 ( .A(n130), .B(n38), .Z(\ab[0][34] ) );
  NR2 U1378 ( .A(n131), .B(n38), .Z(\ab[0][33] ) );
  NR2 U1379 ( .A(n132), .B(n37), .Z(\ab[0][32] ) );
  NR2 U1380 ( .A(n133), .B(n37), .Z(\ab[0][31] ) );
  NR2 U1381 ( .A(n134), .B(n37), .Z(\ab[0][30] ) );
  NR2 U1382 ( .A(n162), .B(n37), .Z(\ab[0][2] ) );
  NR2 U1383 ( .A(n135), .B(n37), .Z(\ab[0][29] ) );
  NR2 U1384 ( .A(n136), .B(n37), .Z(\ab[0][28] ) );
  NR2 U1385 ( .A(n137), .B(n37), .Z(\ab[0][27] ) );
  NR2 U1386 ( .A(n138), .B(n37), .Z(\ab[0][26] ) );
  NR2 U1387 ( .A(n139), .B(n37), .Z(\ab[0][25] ) );
  NR2 U1388 ( .A(n140), .B(n37), .Z(\ab[0][24] ) );
  NR2 U1389 ( .A(n141), .B(n37), .Z(\ab[0][23] ) );
  NR2 U1390 ( .A(n142), .B(n37), .Z(\ab[0][22] ) );
  NR2 U1391 ( .A(n143), .B(n36), .Z(\ab[0][21] ) );
  NR2 U1392 ( .A(n144), .B(n36), .Z(\ab[0][20] ) );
  NR2 U1393 ( .A(n145), .B(n36), .Z(\ab[0][19] ) );
  NR2 U1394 ( .A(n146), .B(n36), .Z(\ab[0][18] ) );
  NR2 U1395 ( .A(n147), .B(n36), .Z(\ab[0][17] ) );
  NR2 U1396 ( .A(n148), .B(n36), .Z(\ab[0][16] ) );
  NR2 U1397 ( .A(n149), .B(n36), .Z(\ab[0][15] ) );
  NR2 U1398 ( .A(n150), .B(n36), .Z(\ab[0][14] ) );
  NR2 U1399 ( .A(n151), .B(n36), .Z(\ab[0][13] ) );
  NR2 U1400 ( .A(n152), .B(n36), .Z(\ab[0][12] ) );
  NR2 U1401 ( .A(n153), .B(n36), .Z(\ab[0][11] ) );
  NR2 U1402 ( .A(n154), .B(n36), .Z(\ab[0][10] ) );
  AN3 U1403 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U1404 ( .A(n41), .B(n163), .Z(\ab[1][1] ) );
endmodule


module LOG_POLY_DW01_add_6 ( A, B, CI, SUM, CO );
  input [123:0] A;
  input [123:0] B;
  output [123:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  AN4P U2 ( .A(n502), .B(n467), .C(n465), .D(n472), .Z(n1) );
  OR2P U3 ( .A(n335), .B(n336), .Z(n2) );
  AN2P U4 ( .A(B[47]), .B(A[47]), .Z(n3) );
  AN2P U5 ( .A(B[67]), .B(A[67]), .Z(n4) );
  AO7 U6 ( .A(n38), .B(n169), .C(n226), .Z(n254) );
  NR2 U7 ( .A(n2), .B(n295), .Z(n279) );
  IVP U8 ( .A(n296), .Z(n295) );
  ND2 U9 ( .A(n265), .B(n266), .Z(n43) );
  ND2 U10 ( .A(n267), .B(n87), .Z(n266) );
  ND4 U11 ( .A(n272), .B(n273), .C(n274), .D(n383), .Z(n271) );
  NR2 U12 ( .A(n368), .B(n369), .Z(n272) );
  NR3 U13 ( .A(n361), .B(n362), .C(n363), .Z(n273) );
  ND2 U14 ( .A(n275), .B(n276), .Z(n274) );
  NR2 U15 ( .A(n297), .B(n3), .Z(n277) );
  ND4 U16 ( .A(n279), .B(n280), .C(n281), .D(n282), .Z(n278) );
  AO7 U17 ( .A(n62), .B(n63), .C(n64), .Z(n60) );
  AO7 U18 ( .A(n189), .B(n158), .C(n190), .Z(n186) );
  ND2 U19 ( .A(n220), .B(n221), .Z(n217) );
  AO6 U20 ( .A(n224), .B(n167), .C(n225), .Z(n220) );
  ND2 U21 ( .A(n87), .B(n222), .Z(n221) );
  NR2 U22 ( .A(n163), .B(n169), .Z(n224) );
  IVP U23 ( .A(n375), .Z(n383) );
  AO2 U24 ( .A(n166), .B(n167), .C(n168), .D(n87), .Z(n126) );
  IVP U25 ( .A(n169), .Z(n166) );
  NR2 U26 ( .A(n169), .B(n170), .Z(n168) );
  IVP U27 ( .A(n339), .Z(n346) );
  IVP U28 ( .A(n364), .Z(n409) );
  IVP U29 ( .A(n399), .Z(n393) );
  AO7 U30 ( .A(n400), .B(n401), .C(n402), .Z(n399) );
  IVP U31 ( .A(n369), .Z(n402) );
  AO7 U32 ( .A(n409), .B(n410), .C(n411), .Z(n401) );
  IVP U33 ( .A(n367), .Z(n361) );
  IVP U34 ( .A(n370), .Z(n368) );
  NR3 U35 ( .A(n89), .B(n63), .C(n523), .Z(n532) );
  ND2 U36 ( .A(n521), .B(n522), .Z(n170) );
  NR2 U37 ( .A(n523), .B(n63), .Z(n522) );
  NR2 U38 ( .A(n89), .B(n88), .Z(n521) );
  NR2 U39 ( .A(n223), .B(n170), .Z(n222) );
  ND2 U40 ( .A(n365), .B(n366), .Z(n362) );
  NR2 U41 ( .A(n523), .B(n63), .Z(n553) );
  NR2 U42 ( .A(n88), .B(n89), .Z(n86) );
  ND2 U43 ( .A(n162), .B(n159), .Z(n134) );
  NR2 U44 ( .A(n146), .B(n158), .Z(n162) );
  ND4 U45 ( .A(n268), .B(n269), .C(n270), .D(n271), .Z(n87) );
  AO7 U46 ( .A(n443), .B(n444), .C(n445), .Z(n269) );
  ND3 U47 ( .A(A[63]), .B(B[63]), .C(n383), .Z(n268) );
  NR2 U48 ( .A(n371), .B(n372), .Z(n270) );
  NR2 U49 ( .A(n306), .B(n307), .Z(n296) );
  ND2 U50 ( .A(n301), .B(n303), .Z(n306) );
  AO7 U51 ( .A(A[44]), .B(B[44]), .C(n302), .Z(n307) );
  AO7 U52 ( .A(n246), .B(n247), .C(n234), .Z(n243) );
  AO7 U53 ( .A(n251), .B(n252), .C(n253), .Z(n248) );
  ND2 U54 ( .A(n308), .B(n309), .Z(n302) );
  IVP U55 ( .A(B[47]), .Z(n308) );
  IVP U56 ( .A(A[47]), .Z(n309) );
  EN U57 ( .A(n238), .B(n239), .Z(SUM[103]) );
  ND2 U58 ( .A(n233), .B(n228), .Z(n239) );
  ND2 U59 ( .A(n235), .B(n242), .Z(n238) );
  ND2 U60 ( .A(n232), .B(n243), .Z(n242) );
  NR2 U61 ( .A(n353), .B(n354), .Z(n282) );
  ND2 U62 ( .A(n319), .B(n323), .Z(n353) );
  AO7 U63 ( .A(A[40]), .B(B[40]), .C(n320), .Z(n354) );
  ND3 U64 ( .A(n487), .B(n1), .C(n488), .Z(n375) );
  NR2 U65 ( .A(n511), .B(n512), .Z(n487) );
  IVP U66 ( .A(n446), .Z(n488) );
  AO7 U67 ( .A(n52), .B(n53), .C(n54), .Z(n51) );
  AO7 U68 ( .A(n179), .B(n180), .C(n153), .Z(n176) );
  AO2 U69 ( .A(B[62]), .B(A[62]), .C(B[61]), .D(A[61]), .Z(n373) );
  ND2 U70 ( .A(n377), .B(n378), .Z(n376) );
  ND3 U71 ( .A(A[60]), .B(B[60]), .C(n379), .Z(n374) );
  AO7 U72 ( .A(n57), .B(n58), .C(n59), .Z(n55) );
  AO7 U73 ( .A(n184), .B(n185), .C(n147), .Z(n181) );
  ND2 U74 ( .A(n349), .B(n350), .Z(n339) );
  IVP U75 ( .A(B[37]), .Z(n349) );
  IVP U76 ( .A(A[37]), .Z(n350) );
  AO3 U77 ( .A(n324), .B(n325), .C(n293), .D(n282), .Z(n314) );
  AO3 U78 ( .A(n328), .B(n332), .C(n333), .D(n334), .Z(n324) );
  NR2 U79 ( .A(n328), .B(n329), .Z(n325) );
  ND2 U80 ( .A(A[33]), .B(B[33]), .Z(n332) );
  AO7 U81 ( .A(n304), .B(n305), .C(n296), .Z(n275) );
  ND2 U82 ( .A(n340), .B(n341), .Z(n304) );
  AO3 U83 ( .A(n2), .B(n314), .C(n315), .D(n316), .Z(n305) );
  ND3 U84 ( .A(A[39]), .B(B[39]), .C(n282), .Z(n340) );
  AO6 U85 ( .A(n380), .B(n381), .C(n382), .Z(n371) );
  AO2 U86 ( .A(B[59]), .B(A[59]), .C(n433), .D(n396), .Z(n380) );
  AO7 U87 ( .A(n392), .B(n393), .C(n370), .Z(n381) );
  ND2 U88 ( .A(n383), .B(n367), .Z(n382) );
  ND2 U89 ( .A(n343), .B(n344), .Z(n337) );
  IVP U90 ( .A(B[39]), .Z(n343) );
  IVP U91 ( .A(A[39]), .Z(n344) );
  ND2 U92 ( .A(n351), .B(n352), .Z(n338) );
  IVP U93 ( .A(B[38]), .Z(n351) );
  IVP U94 ( .A(A[38]), .Z(n352) );
  ND2 U95 ( .A(n355), .B(n356), .Z(n320) );
  IVP U96 ( .A(B[43]), .Z(n355) );
  IVP U97 ( .A(A[43]), .Z(n356) );
  ND2 U98 ( .A(n359), .B(n360), .Z(n319) );
  IVP U99 ( .A(B[42]), .Z(n359) );
  IVP U100 ( .A(A[42]), .Z(n360) );
  ND2 U101 ( .A(n330), .B(n331), .Z(n294) );
  IVP U102 ( .A(B[33]), .Z(n330) );
  IVP U103 ( .A(A[33]), .Z(n331) );
  ND2 U104 ( .A(n310), .B(n311), .Z(n303) );
  IVP U105 ( .A(B[45]), .Z(n310) );
  IVP U106 ( .A(A[45]), .Z(n311) );
  ND2 U107 ( .A(n312), .B(n313), .Z(n301) );
  IVP U108 ( .A(B[46]), .Z(n312) );
  IVP U109 ( .A(A[46]), .Z(n313) );
  ND2 U110 ( .A(n357), .B(n358), .Z(n323) );
  IVP U111 ( .A(B[41]), .Z(n357) );
  IVP U112 ( .A(A[41]), .Z(n358) );
  ND2 U113 ( .A(n84), .B(n85), .Z(n82) );
  ND2 U114 ( .A(n86), .B(n87), .Z(n85) );
  ND2 U115 ( .A(n92), .B(n93), .Z(n90) );
  ND4 U116 ( .A(n338), .B(n342), .C(n337), .D(n282), .Z(n341) );
  AO3 U117 ( .A(n345), .B(n346), .C(n347), .D(n348), .Z(n342) );
  ND2 U118 ( .A(A[36]), .B(B[36]), .Z(n345) );
  ND2 U119 ( .A(B[37]), .B(A[37]), .Z(n347) );
  ND2 U120 ( .A(n338), .B(n339), .Z(n335) );
  AO7 U121 ( .A(A[36]), .B(B[36]), .C(n337), .Z(n336) );
  ND3 U122 ( .A(B[32]), .B(A[32]), .C(n294), .Z(n329) );
  EN U123 ( .A(n51), .B(n5), .Z(SUM[94]) );
  ND2 U124 ( .A(n50), .B(n48), .Z(n5) );
  EN U125 ( .A(n44), .B(n45), .Z(SUM[95]) );
  ND2 U126 ( .A(n46), .B(n47), .Z(n45) );
  ND2 U127 ( .A(n48), .B(n49), .Z(n44) );
  ND2 U128 ( .A(n50), .B(n51), .Z(n49) );
  EN U129 ( .A(n243), .B(n6), .Z(SUM[102]) );
  ND2 U130 ( .A(n232), .B(n235), .Z(n6) );
  EN U131 ( .A(n176), .B(n7), .Z(SUM[110]) );
  ND2 U132 ( .A(n150), .B(n157), .Z(n7) );
  EN U133 ( .A(n171), .B(n172), .Z(SUM[111]) );
  ND2 U134 ( .A(n151), .B(n156), .Z(n172) );
  ND2 U135 ( .A(n157), .B(n175), .Z(n171) );
  ND2 U136 ( .A(n150), .B(n176), .Z(n175) );
  NR2 U137 ( .A(n384), .B(n385), .Z(n367) );
  ND2 U138 ( .A(n379), .B(n377), .Z(n384) );
  AO7 U139 ( .A(A[60]), .B(B[60]), .C(n378), .Z(n385) );
  NR2 U140 ( .A(n394), .B(n395), .Z(n370) );
  ND2 U141 ( .A(n397), .B(n398), .Z(n394) );
  AO7 U142 ( .A(A[56]), .B(B[56]), .C(n396), .Z(n395) );
  ND2 U143 ( .A(n419), .B(n420), .Z(n364) );
  IVP U144 ( .A(B[51]), .Z(n419) );
  IVP U145 ( .A(A[51]), .Z(n420) );
  AO7 U146 ( .A(n126), .B(n127), .C(n128), .Z(n122) );
  AO6 U147 ( .A(n129), .B(n130), .C(n131), .Z(n128) );
  AO7 U148 ( .A(n33), .B(n34), .C(n35), .Z(n32) );
  AO7 U149 ( .A(n113), .B(n114), .C(n115), .Z(n109) );
  NR3 U150 ( .A(n289), .B(n290), .C(n291), .Z(n280) );
  NR2 U151 ( .A(A[31]), .B(B[31]), .Z(n290) );
  ND2 U152 ( .A(n293), .B(n294), .Z(n289) );
  AO7 U153 ( .A(A[32]), .B(B[32]), .C(n292), .Z(n291) );
  ND2 U154 ( .A(n417), .B(n418), .Z(n365) );
  IVP U155 ( .A(B[50]), .Z(n417) );
  IVP U156 ( .A(A[50]), .Z(n418) );
  ND3 U157 ( .A(n529), .B(n530), .C(n531), .Z(n167) );
  ND2 U158 ( .A(n553), .B(n554), .Z(n530) );
  AO6 U159 ( .A(n93), .B(n532), .C(n533), .Z(n531) );
  AO2 U160 ( .A(n566), .B(n65), .C(n567), .D(n566), .Z(n529) );
  ND4 U161 ( .A(n403), .B(n404), .C(n405), .D(n406), .Z(n369) );
  ND2 U162 ( .A(n407), .B(n408), .Z(n403) );
  IVP U163 ( .A(B[52]), .Z(n407) );
  IVP U164 ( .A(A[52]), .Z(n408) );
  AO7 U165 ( .A(n80), .B(n62), .C(n81), .Z(n78) );
  AO7 U166 ( .A(n38), .B(n39), .C(n40), .Z(n36) );
  AO7 U167 ( .A(n216), .B(n189), .C(n197), .Z(n213) );
  AO7 U168 ( .A(n75), .B(n76), .C(n77), .Z(n73) );
  AO7 U169 ( .A(n199), .B(n212), .C(n198), .Z(n209) );
  AO7 U170 ( .A(n412), .B(n413), .C(n414), .Z(n400) );
  ND2 U171 ( .A(n365), .B(n366), .Z(n413) );
  ND3 U172 ( .A(B[48]), .B(A[48]), .C(n364), .Z(n412) );
  ND4 U173 ( .A(B[49]), .B(A[49]), .C(n364), .D(n365), .Z(n414) );
  AO6 U174 ( .A(n298), .B(n299), .C(n300), .Z(n297) );
  AO2 U175 ( .A(B[46]), .B(A[46]), .C(B[45]), .D(A[45]), .Z(n298) );
  ND2 U176 ( .A(n301), .B(n302), .Z(n300) );
  ND3 U177 ( .A(A[44]), .B(B[44]), .C(n303), .Z(n299) );
  AO3 U178 ( .A(n317), .B(n318), .C(n319), .D(n320), .Z(n316) );
  ND2 U179 ( .A(n321), .B(n322), .Z(n318) );
  AN3 U180 ( .A(A[40]), .B(B[40]), .C(n323), .Z(n317) );
  ND2 U181 ( .A(B[41]), .B(A[41]), .Z(n321) );
  AO3 U182 ( .A(A[64]), .B(B[64]), .C(n445), .D(n456), .Z(n512) );
  ND2 U183 ( .A(n415), .B(n416), .Z(n366) );
  IVP U184 ( .A(B[49]), .Z(n415) );
  IVP U185 ( .A(A[49]), .Z(n416) );
  ND2 U186 ( .A(n326), .B(n327), .Z(n293) );
  IVP U187 ( .A(B[35]), .Z(n326) );
  IVP U188 ( .A(A[35]), .Z(n327) );
  ND2 U189 ( .A(n425), .B(n426), .Z(n404) );
  IVP U190 ( .A(B[55]), .Z(n425) );
  IVP U191 ( .A(A[55]), .Z(n426) );
  ND2 U192 ( .A(n427), .B(n428), .Z(n405) );
  IVP U193 ( .A(B[54]), .Z(n427) );
  IVP U194 ( .A(A[54]), .Z(n428) );
  ND2 U195 ( .A(n513), .B(n514), .Z(n456) );
  IVP U196 ( .A(B[65]), .Z(n513) );
  IVP U197 ( .A(A[65]), .Z(n514) );
  ND2 U198 ( .A(n434), .B(n435), .Z(n396) );
  IVP U199 ( .A(B[59]), .Z(n434) );
  IVP U200 ( .A(A[59]), .Z(n435) );
  ND2 U201 ( .A(n390), .B(n391), .Z(n379) );
  IVP U202 ( .A(B[61]), .Z(n390) );
  IVP U203 ( .A(A[61]), .Z(n391) );
  ND2 U204 ( .A(n386), .B(n387), .Z(n378) );
  IVP U205 ( .A(B[62]), .Z(n386) );
  IVP U206 ( .A(A[62]), .Z(n387) );
  ND2 U207 ( .A(n388), .B(n389), .Z(n377) );
  IVP U208 ( .A(B[63]), .Z(n388) );
  IVP U209 ( .A(A[63]), .Z(n389) );
  ND2 U210 ( .A(n69), .B(n568), .Z(n65) );
  AO7 U211 ( .A(n569), .B(n570), .C(n68), .Z(n568) );
  ND2 U212 ( .A(n431), .B(n432), .Z(n406) );
  IVP U213 ( .A(B[53]), .Z(n431) );
  IVP U214 ( .A(A[53]), .Z(n432) );
  ND2 U215 ( .A(n120), .B(n121), .Z(n116) );
  ND2 U216 ( .A(n122), .B(n123), .Z(n121) );
  ND4 U217 ( .A(n457), .B(n458), .C(n459), .D(n460), .Z(n443) );
  NR2 U218 ( .A(n473), .B(n474), .Z(n458) );
  AO3 U219 ( .A(n479), .B(n24), .C(n480), .D(n481), .Z(n457) );
  AN3 U220 ( .A(A[52]), .B(B[52]), .C(n406), .Z(n423) );
  ND3 U221 ( .A(n284), .B(n285), .C(n283), .Z(n281) );
  ND2 U222 ( .A(B[31]), .B(A[31]), .Z(n283) );
  ND2 U223 ( .A(B[30]), .B(A[30]), .Z(n284) );
  ND3 U224 ( .A(A[29]), .B(B[29]), .C(n286), .Z(n285) );
  ND3 U225 ( .A(A[64]), .B(B[64]), .C(n456), .Z(n451) );
  ND2 U226 ( .A(n287), .B(n288), .Z(n286) );
  IVP U227 ( .A(B[30]), .Z(n287) );
  IVP U228 ( .A(A[30]), .Z(n288) );
  ND2 U229 ( .A(n454), .B(n455), .Z(n511) );
  ND2 U230 ( .A(n421), .B(n422), .Z(n392) );
  ND2 U231 ( .A(B[55]), .B(A[55]), .Z(n421) );
  AO3 U232 ( .A(n423), .B(n424), .C(n405), .D(n404), .Z(n422) );
  ND2 U233 ( .A(n429), .B(n430), .Z(n424) );
  EO U234 ( .A(n66), .B(n67), .Z(SUM[91]) );
  AO7 U235 ( .A(n70), .B(n71), .C(n72), .Z(n66) );
  EN U236 ( .A(n25), .B(n26), .Z(SUM[99]) );
  ND2 U237 ( .A(n27), .B(n28), .Z(n26) );
  ND2 U238 ( .A(n29), .B(n30), .Z(n25) );
  ND2 U239 ( .A(n31), .B(n32), .Z(n30) );
  EO U240 ( .A(n204), .B(n205), .Z(SUM[107]) );
  AO7 U241 ( .A(n200), .B(n208), .C(n196), .Z(n204) );
  EN U242 ( .A(n109), .B(n8), .Z(SUM[115]) );
  ND2 U243 ( .A(n110), .B(n107), .Z(n8) );
  ND2 U244 ( .A(n109), .B(n110), .Z(n108) );
  ND4 U245 ( .A(n68), .B(n74), .C(n79), .D(n83), .Z(n63) );
  ND4 U246 ( .A(n61), .B(n56), .C(n50), .D(n46), .Z(n523) );
  ND3 U247 ( .A(n96), .B(n103), .C(n102), .Z(n89) );
  AO7 U248 ( .A(n555), .B(n101), .C(n96), .Z(n91) );
  AO7 U249 ( .A(n436), .B(n437), .C(n438), .Z(n433) );
  ND2 U250 ( .A(B[58]), .B(A[58]), .Z(n438) );
  AO2 U251 ( .A(B[57]), .B(A[57]), .C(B[56]), .D(A[56]), .Z(n436) );
  ND2 U252 ( .A(n397), .B(n398), .Z(n437) );
  AO7 U253 ( .A(A[48]), .B(B[48]), .C(n364), .Z(n363) );
  NR2 U254 ( .A(A[34]), .B(B[34]), .Z(n328) );
  ND2 U255 ( .A(n439), .B(n440), .Z(n398) );
  IVP U256 ( .A(B[57]), .Z(n439) );
  IVP U257 ( .A(A[57]), .Z(n440) );
  ND2 U258 ( .A(n441), .B(n442), .Z(n397) );
  IVP U259 ( .A(B[58]), .Z(n441) );
  IVP U260 ( .A(A[58]), .Z(n442) );
  IVP U261 ( .A(n104), .Z(n88) );
  ND2 U262 ( .A(B[35]), .B(A[35]), .Z(n334) );
  ND2 U263 ( .A(B[34]), .B(A[34]), .Z(n333) );
  ND2 U264 ( .A(B[42]), .B(A[42]), .Z(n322) );
  ND2 U265 ( .A(B[38]), .B(A[38]), .Z(n348) );
  ND2 U266 ( .A(B[51]), .B(A[51]), .Z(n411) );
  ND2 U267 ( .A(A[50]), .B(B[50]), .Z(n410) );
  ND2 U268 ( .A(B[53]), .B(A[53]), .Z(n430) );
  ND2 U269 ( .A(B[54]), .B(A[54]), .Z(n429) );
  EN U270 ( .A(n73), .B(n9), .Z(SUM[90]) );
  ND2 U271 ( .A(n74), .B(n72), .Z(n9) );
  EN U272 ( .A(n55), .B(n10), .Z(SUM[93]) );
  ND2 U273 ( .A(n56), .B(n54), .Z(n10) );
  EN U274 ( .A(n32), .B(n11), .Z(SUM[98]) );
  ND2 U275 ( .A(n31), .B(n29), .Z(n11) );
  EN U276 ( .A(n248), .B(n12), .Z(SUM[101]) );
  ND2 U277 ( .A(n236), .B(n234), .Z(n12) );
  EN U278 ( .A(n209), .B(n13), .Z(SUM[106]) );
  ND2 U279 ( .A(n201), .B(n196), .Z(n13) );
  EN U280 ( .A(n181), .B(n14), .Z(SUM[109]) );
  ND2 U281 ( .A(n165), .B(n153), .Z(n14) );
  EN U282 ( .A(n116), .B(n15), .Z(SUM[114]) );
  ND2 U283 ( .A(n117), .B(n115), .Z(n15) );
  IVP U284 ( .A(n472), .Z(n469) );
  ND4 U285 ( .A(n27), .B(n41), .C(n37), .D(n31), .Z(n169) );
  ND4 U286 ( .A(n233), .B(n232), .C(n236), .D(n237), .Z(n163) );
  AO7 U287 ( .A(n140), .B(n141), .C(n142), .Z(n129) );
  AO6 U288 ( .A(n159), .B(n160), .C(n161), .Z(n140) );
  AO6 U289 ( .A(n143), .B(n144), .C(n145), .Z(n142) );
  AO3 U290 ( .A(n54), .B(n534), .C(n535), .D(n47), .Z(n533) );
  ND2 U291 ( .A(n50), .B(n46), .Z(n534) );
  ND2 U292 ( .A(n536), .B(n46), .Z(n535) );
  AO7 U293 ( .A(n226), .B(n163), .C(n227), .Z(n225) );
  AO6 U294 ( .A(n104), .B(n87), .C(n93), .Z(n98) );
  ND2 U295 ( .A(n191), .B(n192), .Z(n144) );
  AO7 U296 ( .A(n193), .B(n194), .C(n195), .Z(n192) );
  ND2 U297 ( .A(B[43]), .B(A[43]), .Z(n315) );
  EN U298 ( .A(n94), .B(n95), .Z(SUM[87]) );
  ND2 U299 ( .A(n96), .B(n97), .Z(n95) );
  AO7 U300 ( .A(n98), .B(n99), .C(n100), .Z(n94) );
  ND2 U301 ( .A(n102), .B(n103), .Z(n99) );
  EN U302 ( .A(n78), .B(n16), .Z(SUM[89]) );
  ND2 U303 ( .A(n79), .B(n77), .Z(n16) );
  EN U304 ( .A(n60), .B(n17), .Z(SUM[92]) );
  ND2 U305 ( .A(n61), .B(n59), .Z(n17) );
  EN U306 ( .A(n36), .B(n18), .Z(SUM[97]) );
  ND2 U307 ( .A(n37), .B(n35), .Z(n18) );
  EN U308 ( .A(n255), .B(n254), .Z(SUM[100]) );
  ND2 U309 ( .A(n253), .B(n237), .Z(n255) );
  EN U310 ( .A(n213), .B(n19), .Z(SUM[105]) );
  ND2 U311 ( .A(n202), .B(n198), .Z(n19) );
  EN U312 ( .A(n186), .B(n20), .Z(SUM[108]) );
  ND2 U313 ( .A(n164), .B(n147), .Z(n20) );
  EO U314 ( .A(n135), .B(n136), .Z(SUM[112]) );
  AO7 U315 ( .A(n126), .B(n134), .C(n139), .Z(n135) );
  EN U316 ( .A(n122), .B(n21), .Z(SUM[113]) );
  ND2 U317 ( .A(n123), .B(n120), .Z(n21) );
  ND4 U318 ( .A(n164), .B(n165), .C(n150), .D(n151), .Z(n146) );
  AO3 U319 ( .A(n146), .B(n147), .C(n148), .D(n149), .Z(n145) );
  ND3 U320 ( .A(n150), .B(n151), .C(n152), .Z(n149) );
  AO6 U321 ( .A(n154), .B(n151), .C(n155), .Z(n148) );
  EN U322 ( .A(n82), .B(n22), .Z(SUM[88]) );
  ND2 U323 ( .A(n81), .B(n83), .Z(n22) );
  EN U324 ( .A(n42), .B(n43), .Z(SUM[96]) );
  ND2 U325 ( .A(n40), .B(n41), .Z(n42) );
  EN U326 ( .A(n217), .B(n23), .Z(SUM[104]) );
  ND2 U327 ( .A(n197), .B(n203), .Z(n23) );
  ND4 U328 ( .A(n195), .B(n201), .C(n202), .D(n203), .Z(n158) );
  IVP U329 ( .A(n101), .Z(n100) );
  ND2 U330 ( .A(n489), .B(n481), .Z(n446) );
  NR2 U331 ( .A(n494), .B(n495), .Z(n489) );
  ND2 U332 ( .A(n485), .B(n486), .Z(n495) );
  AO7 U333 ( .A(A[72]), .B(B[72]), .C(n480), .Z(n494) );
  AO3 U334 ( .A(A[76]), .B(B[76]), .C(n463), .D(n464), .Z(n477) );
  ND2 U335 ( .A(n492), .B(n493), .Z(n463) );
  IVP U336 ( .A(B[78]), .Z(n492) );
  IVP U337 ( .A(A[78]), .Z(n493) );
  ND2 U338 ( .A(n498), .B(n499), .Z(n485) );
  IVP U339 ( .A(B[73]), .Z(n498) );
  IVP U340 ( .A(A[73]), .Z(n499) );
  ND2 U341 ( .A(n496), .B(n497), .Z(n486) );
  IVP U342 ( .A(B[74]), .Z(n496) );
  IVP U343 ( .A(A[74]), .Z(n497) );
  ND2 U344 ( .A(n490), .B(n491), .Z(n464) );
  IVP U345 ( .A(B[77]), .Z(n490) );
  IVP U346 ( .A(A[77]), .Z(n491) );
  ND2 U347 ( .A(n500), .B(n501), .Z(n480) );
  IVP U348 ( .A(B[75]), .Z(n500) );
  IVP U349 ( .A(A[75]), .Z(n501) );
  ND2 U350 ( .A(n509), .B(n510), .Z(n502) );
  IVP U351 ( .A(B[68]), .Z(n509) );
  IVP U352 ( .A(A[68]), .Z(n510) );
  NR3 U353 ( .A(n482), .B(n483), .C(n484), .Z(n479) );
  AO2 U354 ( .A(B[73]), .B(A[73]), .C(B[72]), .D(A[72]), .Z(n483) );
  IVP U355 ( .A(n486), .Z(n482) );
  IVP U356 ( .A(n485), .Z(n484) );
  AO2 U357 ( .A(B[66]), .B(A[66]), .C(B[65]), .D(A[65]), .Z(n450) );
  IVP U358 ( .A(n455), .Z(n452) );
  IVP U359 ( .A(n454), .Z(n453) );
  ND2 U360 ( .A(n519), .B(n520), .Z(n454) );
  IVP U361 ( .A(B[66]), .Z(n519) );
  IVP U362 ( .A(A[66]), .Z(n520) );
  ND2 U363 ( .A(n517), .B(n518), .Z(n455) );
  IVP U364 ( .A(B[67]), .Z(n517) );
  IVP U365 ( .A(A[67]), .Z(n518) );
  ND2 U366 ( .A(n503), .B(n504), .Z(n472) );
  IVP U367 ( .A(B[69]), .Z(n503) );
  IVP U368 ( .A(A[69]), .Z(n504) );
  ND2 U369 ( .A(n573), .B(n574), .Z(n74) );
  IVP U370 ( .A(B[90]), .Z(n573) );
  IVP U371 ( .A(A[90]), .Z(n574) );
  ND2 U372 ( .A(n575), .B(n576), .Z(n79) );
  IVP U373 ( .A(B[89]), .Z(n575) );
  IVP U374 ( .A(A[89]), .Z(n576) );
  AO7 U375 ( .A(n446), .B(n447), .C(n448), .Z(n444) );
  AO7 U376 ( .A(n449), .B(n4), .C(n1), .Z(n447) );
  ND3 U377 ( .A(A[71]), .B(B[71]), .C(n488), .Z(n448) );
  ND2 U378 ( .A(n505), .B(n506), .Z(n465) );
  IVP U379 ( .A(B[70]), .Z(n505) );
  IVP U380 ( .A(A[70]), .Z(n506) );
  ND2 U381 ( .A(n507), .B(n508), .Z(n467) );
  IVP U382 ( .A(B[71]), .Z(n507) );
  IVP U383 ( .A(A[71]), .Z(n508) );
  ND2 U384 ( .A(n515), .B(n516), .Z(n445) );
  IVP U385 ( .A(B[79]), .Z(n515) );
  IVP U386 ( .A(A[79]), .Z(n516) );
  ND4 U387 ( .A(n465), .B(n466), .C(n467), .D(n488), .Z(n459) );
  AO3 U388 ( .A(n468), .B(n469), .C(n470), .D(n471), .Z(n466) );
  ND2 U389 ( .A(A[68]), .B(B[68]), .Z(n468) );
  AO7 U390 ( .A(n537), .B(n558), .C(n559), .Z(n101) );
  ND2 U391 ( .A(A[84]), .B(B[84]), .Z(n558) );
  AO2 U392 ( .A(B[86]), .B(A[86]), .C(n560), .D(n561), .Z(n559) );
  NR2 U393 ( .A(n524), .B(n525), .Z(n104) );
  ND2 U394 ( .A(n527), .B(n528), .Z(n524) );
  AO7 U395 ( .A(A[80]), .B(B[80]), .C(n526), .Z(n525) );
  ND2 U396 ( .A(n577), .B(n578), .Z(n46) );
  IVP U397 ( .A(B[95]), .Z(n577) );
  IVP U398 ( .A(A[95]), .Z(n578) );
  AO7 U399 ( .A(A[85]), .B(B[85]), .C(n561), .Z(n537) );
  NR3 U400 ( .A(n546), .B(n547), .C(n548), .Z(n542) );
  AO2 U401 ( .A(B[80]), .B(A[80]), .C(B[81]), .D(A[81]), .Z(n546) );
  ND2 U402 ( .A(n556), .B(n557), .Z(n96) );
  IVP U403 ( .A(B[87]), .Z(n556) );
  IVP U404 ( .A(A[87]), .Z(n557) );
  ND2 U405 ( .A(n540), .B(n541), .Z(n93) );
  ND2 U406 ( .A(B[83]), .B(A[83]), .Z(n540) );
  AO7 U407 ( .A(n542), .B(n543), .C(n526), .Z(n541) );
  ND2 U408 ( .A(B[89]), .B(A[89]), .Z(n77) );
  ND2 U409 ( .A(B[88]), .B(A[88]), .Z(n81) );
  ND2 U410 ( .A(n571), .B(n572), .Z(n68) );
  IVP U411 ( .A(B[91]), .Z(n571) );
  IVP U412 ( .A(A[91]), .Z(n572) );
  ND2 U413 ( .A(n581), .B(n582), .Z(n56) );
  IVP U414 ( .A(B[93]), .Z(n581) );
  IVP U415 ( .A(A[93]), .Z(n582) );
  ND2 U416 ( .A(n583), .B(n584), .Z(n61) );
  IVP U417 ( .A(B[92]), .Z(n583) );
  IVP U418 ( .A(A[92]), .Z(n584) );
  ND2 U419 ( .A(n564), .B(n565), .Z(n83) );
  IVP U420 ( .A(B[88]), .Z(n564) );
  IVP U421 ( .A(A[88]), .Z(n565) );
  NR2 U422 ( .A(n477), .B(n478), .Z(n473) );
  ND2 U423 ( .A(A[75]), .B(B[75]), .Z(n478) );
  ND2 U424 ( .A(n562), .B(n563), .Z(n561) );
  IVP U425 ( .A(B[86]), .Z(n562) );
  IVP U426 ( .A(A[86]), .Z(n563) );
  ND2 U427 ( .A(n544), .B(n545), .Z(n526) );
  IVP U428 ( .A(B[83]), .Z(n544) );
  IVP U429 ( .A(A[83]), .Z(n545) );
  ND2 U430 ( .A(n551), .B(n552), .Z(n528) );
  IVP U431 ( .A(B[81]), .Z(n551) );
  IVP U432 ( .A(A[81]), .Z(n552) );
  ND2 U433 ( .A(n549), .B(n550), .Z(n527) );
  IVP U434 ( .A(B[82]), .Z(n549) );
  IVP U435 ( .A(A[82]), .Z(n550) );
  ND4 U436 ( .A(B[76]), .B(A[76]), .C(n463), .D(n464), .Z(n462) );
  ND2 U437 ( .A(n579), .B(n580), .Z(n50) );
  IVP U438 ( .A(B[94]), .Z(n579) );
  IVP U439 ( .A(A[94]), .Z(n580) );
  ND3 U440 ( .A(A[77]), .B(B[77]), .C(n463), .Z(n461) );
  ND2 U441 ( .A(n259), .B(n260), .Z(n31) );
  IVP U442 ( .A(B[98]), .Z(n259) );
  IVP U443 ( .A(A[98]), .Z(n260) );
  ND2 U444 ( .A(n244), .B(n245), .Z(n232) );
  IVP U445 ( .A(B[102]), .Z(n244) );
  IVP U446 ( .A(A[102]), .Z(n245) );
  ND2 U447 ( .A(n263), .B(n264), .Z(n27) );
  IVP U448 ( .A(B[99]), .Z(n263) );
  IVP U449 ( .A(A[99]), .Z(n264) );
  ND2 U450 ( .A(n240), .B(n241), .Z(n233) );
  IVP U451 ( .A(B[103]), .Z(n240) );
  IVP U452 ( .A(A[103]), .Z(n241) );
  ND2 U453 ( .A(n261), .B(n262), .Z(n37) );
  IVP U454 ( .A(B[97]), .Z(n261) );
  IVP U455 ( .A(A[97]), .Z(n262) );
  ND2 U456 ( .A(n249), .B(n250), .Z(n236) );
  IVP U457 ( .A(B[101]), .Z(n249) );
  IVP U458 ( .A(A[101]), .Z(n250) );
  ND2 U459 ( .A(n214), .B(n215), .Z(n202) );
  IVP U460 ( .A(B[105]), .Z(n214) );
  IVP U461 ( .A(A[105]), .Z(n215) );
  ND2 U462 ( .A(n210), .B(n211), .Z(n201) );
  IVP U463 ( .A(B[106]), .Z(n210) );
  IVP U464 ( .A(A[106]), .Z(n211) );
  ND2 U465 ( .A(n538), .B(n539), .Z(n103) );
  IVP U466 ( .A(B[84]), .Z(n538) );
  IVP U467 ( .A(A[84]), .Z(n539) );
  ND2 U468 ( .A(n28), .B(n256), .Z(n160) );
  AO3 U469 ( .A(n257), .B(n258), .C(n31), .D(n27), .Z(n256) );
  ND2 U470 ( .A(n35), .B(n29), .Z(n258) );
  AN3 U471 ( .A(A[96]), .B(B[96]), .C(n37), .Z(n257) );
  ND2 U472 ( .A(n228), .B(n229), .Z(n161) );
  AO3 U473 ( .A(n230), .B(n231), .C(n232), .D(n233), .Z(n229) );
  ND2 U474 ( .A(n234), .B(n235), .Z(n231) );
  AN3 U475 ( .A(A[100]), .B(B[100]), .C(n236), .Z(n230) );
  ND2 U476 ( .A(B[69]), .B(A[69]), .Z(n471) );
  ND2 U477 ( .A(B[70]), .B(A[70]), .Z(n470) );
  ND2 U478 ( .A(n475), .B(n476), .Z(n474) );
  ND2 U479 ( .A(B[78]), .B(A[78]), .Z(n475) );
  ND2 U480 ( .A(B[79]), .B(A[79]), .Z(n476) );
  AN2P U481 ( .A(B[74]), .B(A[74]), .Z(n24) );
  ND2 U482 ( .A(n173), .B(n174), .Z(n151) );
  IVP U483 ( .A(B[111]), .Z(n173) );
  IVP U484 ( .A(A[111]), .Z(n174) );
  ND2 U485 ( .A(B[93]), .B(A[93]), .Z(n54) );
  ND2 U486 ( .A(B[98]), .B(A[98]), .Z(n29) );
  ND2 U487 ( .A(B[97]), .B(A[97]), .Z(n35) );
  ND2 U488 ( .A(B[104]), .B(A[104]), .Z(n197) );
  ND2 U489 ( .A(B[101]), .B(A[101]), .Z(n234) );
  ND2 U490 ( .A(B[105]), .B(A[105]), .Z(n198) );
  ND2 U491 ( .A(B[102]), .B(A[102]), .Z(n235) );
  ND2 U492 ( .A(B[90]), .B(A[90]), .Z(n72) );
  ND2 U493 ( .A(B[94]), .B(A[94]), .Z(n48) );
  ND2 U494 ( .A(B[110]), .B(A[110]), .Z(n157) );
  ND2 U495 ( .A(B[95]), .B(A[95]), .Z(n47) );
  ND2 U496 ( .A(B[87]), .B(A[87]), .Z(n97) );
  ND2 U497 ( .A(B[111]), .B(A[111]), .Z(n156) );
  ND2 U498 ( .A(B[91]), .B(A[91]), .Z(n69) );
  ND2 U499 ( .A(n177), .B(n178), .Z(n150) );
  IVP U500 ( .A(B[110]), .Z(n177) );
  IVP U501 ( .A(A[110]), .Z(n178) );
  ND2 U502 ( .A(n206), .B(n207), .Z(n195) );
  IVP U503 ( .A(B[107]), .Z(n206) );
  IVP U504 ( .A(A[107]), .Z(n207) );
  ND2 U505 ( .A(B[92]), .B(A[92]), .Z(n59) );
  ND2 U506 ( .A(n218), .B(n219), .Z(n203) );
  IVP U507 ( .A(B[104]), .Z(n218) );
  IVP U508 ( .A(A[104]), .Z(n219) );
  ND2 U509 ( .A(n182), .B(n183), .Z(n165) );
  IVP U510 ( .A(B[109]), .Z(n182) );
  IVP U511 ( .A(A[109]), .Z(n183) );
  ND2 U512 ( .A(n187), .B(n188), .Z(n164) );
  IVP U513 ( .A(B[108]), .Z(n187) );
  IVP U514 ( .A(A[108]), .Z(n188) );
  ND2 U515 ( .A(B[109]), .B(A[109]), .Z(n153) );
  ND2 U516 ( .A(B[106]), .B(A[106]), .Z(n196) );
  ND2 U517 ( .A(B[99]), .B(A[99]), .Z(n28) );
  ND2 U518 ( .A(B[103]), .B(A[103]), .Z(n228) );
  ND2 U519 ( .A(B[108]), .B(A[108]), .Z(n147) );
  ND2 U520 ( .A(B[107]), .B(A[107]), .Z(n191) );
  ND2 U521 ( .A(n137), .B(n138), .Z(n130) );
  IVP U522 ( .A(B[112]), .Z(n137) );
  IVP U523 ( .A(A[112]), .Z(n138) );
  ND2 U524 ( .A(B[112]), .B(A[112]), .Z(n132) );
  ND2 U525 ( .A(B[96]), .B(A[96]), .Z(n40) );
  ND2 U526 ( .A(B[100]), .B(A[100]), .Z(n253) );
  ND2 U527 ( .A(n124), .B(n125), .Z(n123) );
  IVP U528 ( .A(B[113]), .Z(n124) );
  IVP U529 ( .A(A[113]), .Z(n125) );
  ND2 U530 ( .A(B[113]), .B(A[113]), .Z(n120) );
  ND2 U531 ( .A(n118), .B(n119), .Z(n117) );
  IVP U532 ( .A(B[114]), .Z(n118) );
  IVP U533 ( .A(A[114]), .Z(n119) );
  ND2 U534 ( .A(B[114]), .B(A[114]), .Z(n115) );
  ND2 U535 ( .A(n111), .B(n112), .Z(n110) );
  IVP U536 ( .A(B[115]), .Z(n111) );
  IVP U537 ( .A(A[115]), .Z(n112) );
  ND2 U538 ( .A(B[115]), .B(A[115]), .Z(n107) );
  EO U539 ( .A(n105), .B(n106), .Z(SUM[116]) );
  EO U540 ( .A(B[116]), .B(A[116]), .Z(n106) );
  IVA U541 ( .A(n36), .Z(n34) );
  IVA U542 ( .A(n37), .Z(n33) );
  IVA U543 ( .A(n41), .Z(n39) );
  IVA U544 ( .A(n55), .Z(n53) );
  IVA U545 ( .A(n56), .Z(n52) );
  IVA U546 ( .A(n60), .Z(n58) );
  IVA U547 ( .A(n61), .Z(n57) );
  IVA U548 ( .A(n65), .Z(n64) );
  AN2P U549 ( .A(n68), .B(n69), .Z(n67) );
  IVA U550 ( .A(n73), .Z(n71) );
  IVA U551 ( .A(n78), .Z(n76) );
  IVA U552 ( .A(n82), .Z(n62) );
  IVA U553 ( .A(n83), .Z(n80) );
  AN2P U554 ( .A(n90), .B(n91), .Z(n84) );
  IVA U555 ( .A(n89), .Z(n92) );
  ND2 U556 ( .A(n107), .B(n108), .Z(n105) );
  IVA U557 ( .A(n116), .Z(n114) );
  IVA U558 ( .A(n117), .Z(n113) );
  IVA U559 ( .A(n132), .Z(n131) );
  ND2 U560 ( .A(n133), .B(n130), .Z(n127) );
  IVA U561 ( .A(n134), .Z(n133) );
  AN2P U562 ( .A(n130), .B(n132), .Z(n136) );
  IVA U563 ( .A(n129), .Z(n139) );
  IVA U564 ( .A(n153), .Z(n152) );
  IVA U565 ( .A(n156), .Z(n155) );
  IVA U566 ( .A(n157), .Z(n154) );
  IVA U567 ( .A(n146), .Z(n143) );
  OR2 U568 ( .A(n158), .B(n146), .Z(n141) );
  IVA U569 ( .A(n163), .Z(n159) );
  IVA U570 ( .A(n181), .Z(n180) );
  IVA U571 ( .A(n165), .Z(n179) );
  IVA U572 ( .A(n186), .Z(n185) );
  IVA U573 ( .A(n164), .Z(n184) );
  IVA U574 ( .A(n144), .Z(n190) );
  IVA U575 ( .A(n196), .Z(n194) );
  AO1P U576 ( .A(n197), .B(n198), .C(n199), .D(n200), .Z(n193) );
  AN2P U577 ( .A(n195), .B(n191), .Z(n205) );
  IVA U578 ( .A(n209), .Z(n208) );
  IVA U579 ( .A(n201), .Z(n200) );
  IVA U580 ( .A(n213), .Z(n212) );
  IVA U581 ( .A(n202), .Z(n199) );
  IVA U582 ( .A(n217), .Z(n189) );
  IVA U583 ( .A(n203), .Z(n216) );
  OR2 U584 ( .A(n169), .B(n163), .Z(n223) );
  IVA U585 ( .A(n161), .Z(n227) );
  IVA U586 ( .A(n248), .Z(n247) );
  IVA U587 ( .A(n236), .Z(n246) );
  IVA U588 ( .A(n254), .Z(n252) );
  IVA U589 ( .A(n237), .Z(n251) );
  IVA U590 ( .A(n160), .Z(n226) );
  OR2 U591 ( .A(A[96]), .B(B[96]), .Z(n41) );
  IVA U592 ( .A(n43), .Z(n38) );
  AN2P U593 ( .A(n277), .B(n278), .Z(n276) );
  OR2 U594 ( .A(A[34]), .B(B[34]), .Z(n292) );
  AO1P U595 ( .A(n373), .B(n374), .C(n375), .D(n376), .Z(n372) );
  AO1P U596 ( .A(n450), .B(n451), .C(n452), .D(n453), .Z(n449) );
  AN2P U597 ( .A(n461), .B(n462), .Z(n460) );
  IVA U598 ( .A(n477), .Z(n481) );
  IVA U599 ( .A(n170), .Z(n267) );
  IVA U600 ( .A(n167), .Z(n265) );
  IVA U601 ( .A(n48), .Z(n536) );
  IVA U602 ( .A(n537), .Z(n102) );
  AN2P U603 ( .A(B[82]), .B(A[82]), .Z(n543) );
  IVA U604 ( .A(n527), .Z(n548) );
  IVA U605 ( .A(n528), .Z(n547) );
  IVA U606 ( .A(n91), .Z(n554) );
  AN2P U607 ( .A(A[85]), .B(B[85]), .Z(n560) );
  IVA U608 ( .A(n97), .Z(n555) );
  IVA U609 ( .A(n59), .Z(n567) );
  IVA U610 ( .A(n72), .Z(n570) );
  AO1P U611 ( .A(n81), .B(n77), .C(n75), .D(n70), .Z(n569) );
  IVA U612 ( .A(n74), .Z(n70) );
  IVA U613 ( .A(n79), .Z(n75) );
  IVA U614 ( .A(n523), .Z(n566) );
  OR2 U615 ( .A(A[100]), .B(B[100]), .Z(n237) );
endmodule


module LOG_POLY_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [29:0] A;
  input [95:0] B;
  output [125:0] PRODUCT;
  input TC;
  wire   \ab[29][95] , \ab[29][94] , \ab[29][93] , \ab[29][92] , \ab[29][91] ,
         \ab[29][90] , \ab[29][89] , \ab[29][88] , \ab[29][87] , \ab[29][86] ,
         \ab[29][85] , \ab[29][84] , \ab[29][83] , \ab[29][82] , \ab[29][81] ,
         \ab[29][80] , \ab[29][79] , \ab[29][78] , \ab[29][77] , \ab[29][76] ,
         \ab[29][75] , \ab[29][74] , \ab[29][73] , \ab[29][72] , \ab[29][71] ,
         \ab[29][70] , \ab[29][69] , \ab[29][68] , \ab[29][67] , \ab[29][66] ,
         \ab[29][65] , \ab[29][64] , \ab[29][63] , \ab[29][62] , \ab[29][61] ,
         \ab[29][60] , \ab[29][59] , \ab[29][58] , \ab[29][57] , \ab[29][56] ,
         \ab[29][55] , \ab[29][54] , \ab[29][53] , \ab[29][52] , \ab[29][51] ,
         \ab[29][50] , \ab[29][49] , \ab[29][48] , \ab[29][47] , \ab[29][46] ,
         \ab[29][45] , \ab[29][44] , \ab[29][43] , \ab[29][42] , \ab[29][41] ,
         \ab[29][40] , \ab[29][39] , \ab[29][38] , \ab[29][37] , \ab[29][36] ,
         \ab[29][35] , \ab[29][34] , \ab[29][33] , \ab[29][32] , \ab[29][31] ,
         \ab[29][30] , \ab[29][29] , \ab[29][28] , \ab[29][27] , \ab[29][26] ,
         \ab[29][25] , \ab[29][24] , \ab[29][23] , \ab[29][22] , \ab[29][21] ,
         \ab[29][20] , \ab[29][19] , \ab[29][18] , \ab[29][17] , \ab[29][16] ,
         \ab[29][15] , \ab[29][14] , \ab[29][13] , \ab[29][12] , \ab[29][11] ,
         \ab[29][10] , \ab[29][9] , \ab[29][8] , \ab[29][7] , \ab[29][6] ,
         \ab[29][5] , \ab[29][4] , \ab[29][3] , \ab[29][2] , \ab[29][1] ,
         \ab[29][0] , \ab[28][95] , \ab[28][94] , \ab[28][93] , \ab[28][92] ,
         \ab[28][91] , \ab[28][90] , \ab[28][89] , \ab[28][88] , \ab[28][87] ,
         \ab[28][86] , \ab[28][85] , \ab[28][84] , \ab[28][83] , \ab[28][82] ,
         \ab[28][81] , \ab[28][80] , \ab[28][79] , \ab[28][78] , \ab[28][77] ,
         \ab[28][76] , \ab[28][75] , \ab[28][74] , \ab[28][73] , \ab[28][72] ,
         \ab[28][71] , \ab[28][70] , \ab[28][69] , \ab[28][68] , \ab[28][67] ,
         \ab[28][66] , \ab[28][65] , \ab[28][64] , \ab[28][63] , \ab[28][62] ,
         \ab[28][61] , \ab[28][60] , \ab[28][59] , \ab[28][58] , \ab[28][57] ,
         \ab[28][56] , \ab[28][55] , \ab[28][54] , \ab[28][53] , \ab[28][52] ,
         \ab[28][51] , \ab[28][50] , \ab[28][49] , \ab[28][48] , \ab[28][47] ,
         \ab[28][46] , \ab[28][45] , \ab[28][44] , \ab[28][43] , \ab[28][42] ,
         \ab[28][41] , \ab[28][40] , \ab[28][39] , \ab[28][38] , \ab[28][37] ,
         \ab[28][36] , \ab[28][35] , \ab[28][34] , \ab[28][33] , \ab[28][32] ,
         \ab[28][31] , \ab[28][30] , \ab[28][29] , \ab[28][28] , \ab[28][27] ,
         \ab[28][26] , \ab[28][25] , \ab[28][24] , \ab[28][23] , \ab[28][22] ,
         \ab[28][21] , \ab[28][20] , \ab[28][19] , \ab[28][18] , \ab[28][17] ,
         \ab[28][16] , \ab[28][15] , \ab[28][14] , \ab[28][13] , \ab[28][12] ,
         \ab[28][11] , \ab[28][10] , \ab[28][9] , \ab[28][8] , \ab[28][7] ,
         \ab[28][6] , \ab[28][5] , \ab[28][4] , \ab[28][3] , \ab[28][2] ,
         \ab[28][1] , \ab[28][0] , \ab[27][95] , \ab[27][94] , \ab[27][93] ,
         \ab[27][92] , \ab[27][91] , \ab[27][90] , \ab[27][89] , \ab[27][88] ,
         \ab[27][87] , \ab[27][86] , \ab[27][85] , \ab[27][84] , \ab[27][83] ,
         \ab[27][82] , \ab[27][81] , \ab[27][80] , \ab[27][79] , \ab[27][78] ,
         \ab[27][77] , \ab[27][76] , \ab[27][75] , \ab[27][74] , \ab[27][73] ,
         \ab[27][72] , \ab[27][71] , \ab[27][70] , \ab[27][69] , \ab[27][68] ,
         \ab[27][67] , \ab[27][66] , \ab[27][65] , \ab[27][64] , \ab[27][63] ,
         \ab[27][62] , \ab[27][61] , \ab[27][60] , \ab[27][59] , \ab[27][58] ,
         \ab[27][57] , \ab[27][56] , \ab[27][55] , \ab[27][54] , \ab[27][53] ,
         \ab[27][52] , \ab[27][51] , \ab[27][50] , \ab[27][49] , \ab[27][48] ,
         \ab[27][47] , \ab[27][46] , \ab[27][45] , \ab[27][44] , \ab[27][43] ,
         \ab[27][42] , \ab[27][41] , \ab[27][40] , \ab[27][39] , \ab[27][38] ,
         \ab[27][37] , \ab[27][36] , \ab[27][35] , \ab[27][34] , \ab[27][33] ,
         \ab[27][32] , \ab[27][31] , \ab[27][30] , \ab[27][29] , \ab[27][28] ,
         \ab[27][27] , \ab[27][26] , \ab[27][25] , \ab[27][24] , \ab[27][23] ,
         \ab[27][22] , \ab[27][21] , \ab[27][20] , \ab[27][19] , \ab[27][18] ,
         \ab[27][17] , \ab[27][16] , \ab[27][15] , \ab[27][14] , \ab[27][13] ,
         \ab[27][12] , \ab[27][11] , \ab[27][10] , \ab[27][9] , \ab[27][8] ,
         \ab[27][7] , \ab[27][6] , \ab[27][5] , \ab[27][4] , \ab[27][3] ,
         \ab[27][2] , \ab[27][1] , \ab[27][0] , \ab[26][95] , \ab[26][94] ,
         \ab[26][93] , \ab[26][92] , \ab[26][91] , \ab[26][90] , \ab[26][89] ,
         \ab[26][88] , \ab[26][87] , \ab[26][86] , \ab[26][85] , \ab[26][84] ,
         \ab[26][83] , \ab[26][82] , \ab[26][81] , \ab[26][80] , \ab[26][79] ,
         \ab[26][78] , \ab[26][77] , \ab[26][76] , \ab[26][75] , \ab[26][74] ,
         \ab[26][73] , \ab[26][72] , \ab[26][71] , \ab[26][70] , \ab[26][69] ,
         \ab[26][68] , \ab[26][67] , \ab[26][66] , \ab[26][65] , \ab[26][64] ,
         \ab[26][63] , \ab[26][62] , \ab[26][61] , \ab[26][60] , \ab[26][59] ,
         \ab[26][58] , \ab[26][57] , \ab[26][56] , \ab[26][55] , \ab[26][54] ,
         \ab[26][53] , \ab[26][52] , \ab[26][51] , \ab[26][50] , \ab[26][49] ,
         \ab[26][48] , \ab[26][47] , \ab[26][46] , \ab[26][45] , \ab[26][44] ,
         \ab[26][43] , \ab[26][42] , \ab[26][41] , \ab[26][40] , \ab[26][39] ,
         \ab[26][38] , \ab[26][37] , \ab[26][36] , \ab[26][35] , \ab[26][34] ,
         \ab[26][33] , \ab[26][32] , \ab[26][31] , \ab[26][30] , \ab[26][29] ,
         \ab[26][28] , \ab[26][27] , \ab[26][26] , \ab[26][25] , \ab[26][24] ,
         \ab[26][23] , \ab[26][22] , \ab[26][21] , \ab[26][20] , \ab[26][19] ,
         \ab[26][18] , \ab[26][17] , \ab[26][16] , \ab[26][15] , \ab[26][14] ,
         \ab[26][13] , \ab[26][12] , \ab[26][11] , \ab[26][10] , \ab[26][9] ,
         \ab[26][8] , \ab[26][7] , \ab[26][6] , \ab[26][5] , \ab[26][4] ,
         \ab[26][3] , \ab[26][2] , \ab[26][1] , \ab[26][0] , \ab[25][95] ,
         \ab[25][94] , \ab[25][93] , \ab[25][92] , \ab[25][91] , \ab[25][90] ,
         \ab[25][89] , \ab[25][88] , \ab[25][87] , \ab[25][86] , \ab[25][85] ,
         \ab[25][84] , \ab[25][83] , \ab[25][82] , \ab[25][81] , \ab[25][80] ,
         \ab[25][79] , \ab[25][78] , \ab[25][77] , \ab[25][76] , \ab[25][75] ,
         \ab[25][74] , \ab[25][73] , \ab[25][72] , \ab[25][71] , \ab[25][70] ,
         \ab[25][69] , \ab[25][68] , \ab[25][67] , \ab[25][66] , \ab[25][65] ,
         \ab[25][64] , \ab[25][63] , \ab[25][62] , \ab[25][61] , \ab[25][60] ,
         \ab[25][59] , \ab[25][58] , \ab[25][57] , \ab[25][56] , \ab[25][55] ,
         \ab[25][54] , \ab[25][53] , \ab[25][52] , \ab[25][51] , \ab[25][50] ,
         \ab[25][49] , \ab[25][48] , \ab[25][47] , \ab[25][46] , \ab[25][45] ,
         \ab[25][44] , \ab[25][43] , \ab[25][42] , \ab[25][41] , \ab[25][40] ,
         \ab[25][39] , \ab[25][38] , \ab[25][37] , \ab[25][36] , \ab[25][35] ,
         \ab[25][34] , \ab[25][33] , \ab[25][32] , \ab[25][31] , \ab[25][30] ,
         \ab[25][29] , \ab[25][28] , \ab[25][27] , \ab[25][26] , \ab[25][25] ,
         \ab[25][24] , \ab[25][23] , \ab[25][22] , \ab[25][21] , \ab[25][20] ,
         \ab[25][19] , \ab[25][18] , \ab[25][17] , \ab[25][16] , \ab[25][15] ,
         \ab[25][14] , \ab[25][13] , \ab[25][12] , \ab[25][11] , \ab[25][10] ,
         \ab[25][9] , \ab[25][8] , \ab[25][7] , \ab[25][6] , \ab[25][5] ,
         \ab[25][4] , \ab[25][3] , \ab[25][2] , \ab[25][1] , \ab[25][0] ,
         \ab[24][95] , \ab[24][94] , \ab[24][93] , \ab[24][92] , \ab[24][91] ,
         \ab[24][90] , \ab[24][89] , \ab[24][88] , \ab[24][87] , \ab[24][86] ,
         \ab[24][85] , \ab[24][84] , \ab[24][83] , \ab[24][82] , \ab[24][81] ,
         \ab[24][80] , \ab[24][79] , \ab[24][78] , \ab[24][77] , \ab[24][76] ,
         \ab[24][75] , \ab[24][74] , \ab[24][73] , \ab[24][72] , \ab[24][71] ,
         \ab[24][70] , \ab[24][69] , \ab[24][68] , \ab[24][67] , \ab[24][66] ,
         \ab[24][65] , \ab[24][64] , \ab[24][63] , \ab[24][62] , \ab[24][61] ,
         \ab[24][60] , \ab[24][59] , \ab[24][58] , \ab[24][57] , \ab[24][56] ,
         \ab[24][55] , \ab[24][54] , \ab[24][53] , \ab[24][52] , \ab[24][51] ,
         \ab[24][50] , \ab[24][49] , \ab[24][48] , \ab[24][47] , \ab[24][46] ,
         \ab[24][45] , \ab[24][44] , \ab[24][43] , \ab[24][42] , \ab[24][41] ,
         \ab[24][40] , \ab[24][39] , \ab[24][38] , \ab[24][37] , \ab[24][36] ,
         \ab[24][35] , \ab[24][34] , \ab[24][33] , \ab[24][32] , \ab[24][31] ,
         \ab[24][30] , \ab[24][29] , \ab[24][28] , \ab[24][27] , \ab[24][26] ,
         \ab[24][25] , \ab[24][24] , \ab[24][23] , \ab[24][22] , \ab[24][21] ,
         \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] , \ab[24][16] ,
         \ab[24][15] , \ab[24][14] , \ab[24][13] , \ab[24][12] , \ab[24][11] ,
         \ab[24][10] , \ab[24][9] , \ab[24][8] , \ab[24][7] , \ab[24][6] ,
         \ab[24][5] , \ab[24][4] , \ab[24][3] , \ab[24][2] , \ab[24][1] ,
         \ab[24][0] , \ab[23][95] , \ab[23][94] , \ab[23][93] , \ab[23][92] ,
         \ab[23][91] , \ab[23][90] , \ab[23][89] , \ab[23][88] , \ab[23][87] ,
         \ab[23][86] , \ab[23][85] , \ab[23][84] , \ab[23][83] , \ab[23][82] ,
         \ab[23][81] , \ab[23][80] , \ab[23][79] , \ab[23][78] , \ab[23][77] ,
         \ab[23][76] , \ab[23][75] , \ab[23][74] , \ab[23][73] , \ab[23][72] ,
         \ab[23][71] , \ab[23][70] , \ab[23][69] , \ab[23][68] , \ab[23][67] ,
         \ab[23][66] , \ab[23][65] , \ab[23][64] , \ab[23][63] , \ab[23][62] ,
         \ab[23][61] , \ab[23][60] , \ab[23][59] , \ab[23][58] , \ab[23][57] ,
         \ab[23][56] , \ab[23][55] , \ab[23][54] , \ab[23][53] , \ab[23][52] ,
         \ab[23][51] , \ab[23][50] , \ab[23][49] , \ab[23][48] , \ab[23][47] ,
         \ab[23][46] , \ab[23][45] , \ab[23][44] , \ab[23][43] , \ab[23][42] ,
         \ab[23][41] , \ab[23][40] , \ab[23][39] , \ab[23][38] , \ab[23][37] ,
         \ab[23][36] , \ab[23][35] , \ab[23][34] , \ab[23][33] , \ab[23][32] ,
         \ab[23][31] , \ab[23][30] , \ab[23][29] , \ab[23][28] , \ab[23][27] ,
         \ab[23][26] , \ab[23][25] , \ab[23][24] , \ab[23][23] , \ab[23][22] ,
         \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] , \ab[23][17] ,
         \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] , \ab[23][12] ,
         \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] , \ab[23][7] ,
         \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] , \ab[23][2] ,
         \ab[23][1] , \ab[23][0] , \ab[22][95] , \ab[22][94] , \ab[22][93] ,
         \ab[22][92] , \ab[22][91] , \ab[22][90] , \ab[22][89] , \ab[22][88] ,
         \ab[22][87] , \ab[22][86] , \ab[22][85] , \ab[22][84] , \ab[22][83] ,
         \ab[22][82] , \ab[22][81] , \ab[22][80] , \ab[22][79] , \ab[22][78] ,
         \ab[22][77] , \ab[22][76] , \ab[22][75] , \ab[22][74] , \ab[22][73] ,
         \ab[22][72] , \ab[22][71] , \ab[22][70] , \ab[22][69] , \ab[22][68] ,
         \ab[22][67] , \ab[22][66] , \ab[22][65] , \ab[22][64] , \ab[22][63] ,
         \ab[22][62] , \ab[22][61] , \ab[22][60] , \ab[22][59] , \ab[22][58] ,
         \ab[22][57] , \ab[22][56] , \ab[22][55] , \ab[22][54] , \ab[22][53] ,
         \ab[22][52] , \ab[22][51] , \ab[22][50] , \ab[22][49] , \ab[22][48] ,
         \ab[22][47] , \ab[22][46] , \ab[22][45] , \ab[22][44] , \ab[22][43] ,
         \ab[22][42] , \ab[22][41] , \ab[22][40] , \ab[22][39] , \ab[22][38] ,
         \ab[22][37] , \ab[22][36] , \ab[22][35] , \ab[22][34] , \ab[22][33] ,
         \ab[22][32] , \ab[22][31] , \ab[22][30] , \ab[22][29] , \ab[22][28] ,
         \ab[22][27] , \ab[22][26] , \ab[22][25] , \ab[22][24] , \ab[22][23] ,
         \ab[22][22] , \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] ,
         \ab[22][17] , \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] ,
         \ab[22][12] , \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] ,
         \ab[22][7] , \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] ,
         \ab[22][2] , \ab[22][1] , \ab[22][0] , \ab[21][95] , \ab[21][94] ,
         \ab[21][93] , \ab[21][92] , \ab[21][91] , \ab[21][90] , \ab[21][89] ,
         \ab[21][88] , \ab[21][87] , \ab[21][86] , \ab[21][85] , \ab[21][84] ,
         \ab[21][83] , \ab[21][82] , \ab[21][81] , \ab[21][80] , \ab[21][79] ,
         \ab[21][78] , \ab[21][77] , \ab[21][76] , \ab[21][75] , \ab[21][74] ,
         \ab[21][73] , \ab[21][72] , \ab[21][71] , \ab[21][70] , \ab[21][69] ,
         \ab[21][68] , \ab[21][67] , \ab[21][66] , \ab[21][65] , \ab[21][64] ,
         \ab[21][63] , \ab[21][62] , \ab[21][61] , \ab[21][60] , \ab[21][59] ,
         \ab[21][58] , \ab[21][57] , \ab[21][56] , \ab[21][55] , \ab[21][54] ,
         \ab[21][53] , \ab[21][52] , \ab[21][51] , \ab[21][50] , \ab[21][49] ,
         \ab[21][48] , \ab[21][47] , \ab[21][46] , \ab[21][45] , \ab[21][44] ,
         \ab[21][43] , \ab[21][42] , \ab[21][41] , \ab[21][40] , \ab[21][39] ,
         \ab[21][38] , \ab[21][37] , \ab[21][36] , \ab[21][35] , \ab[21][34] ,
         \ab[21][33] , \ab[21][32] , \ab[21][31] , \ab[21][30] , \ab[21][29] ,
         \ab[21][28] , \ab[21][27] , \ab[21][26] , \ab[21][25] , \ab[21][24] ,
         \ab[21][23] , \ab[21][22] , \ab[21][21] , \ab[21][20] , \ab[21][19] ,
         \ab[21][18] , \ab[21][17] , \ab[21][16] , \ab[21][15] , \ab[21][14] ,
         \ab[21][13] , \ab[21][12] , \ab[21][11] , \ab[21][10] , \ab[21][9] ,
         \ab[21][8] , \ab[21][7] , \ab[21][6] , \ab[21][5] , \ab[21][4] ,
         \ab[21][3] , \ab[21][2] , \ab[21][1] , \ab[21][0] , \ab[20][95] ,
         \ab[20][94] , \ab[20][93] , \ab[20][92] , \ab[20][91] , \ab[20][90] ,
         \ab[20][89] , \ab[20][88] , \ab[20][87] , \ab[20][86] , \ab[20][85] ,
         \ab[20][84] , \ab[20][83] , \ab[20][82] , \ab[20][81] , \ab[20][80] ,
         \ab[20][79] , \ab[20][78] , \ab[20][77] , \ab[20][76] , \ab[20][75] ,
         \ab[20][74] , \ab[20][73] , \ab[20][72] , \ab[20][71] , \ab[20][70] ,
         \ab[20][69] , \ab[20][68] , \ab[20][67] , \ab[20][66] , \ab[20][65] ,
         \ab[20][64] , \ab[20][63] , \ab[20][62] , \ab[20][61] , \ab[20][60] ,
         \ab[20][59] , \ab[20][58] , \ab[20][57] , \ab[20][56] , \ab[20][55] ,
         \ab[20][54] , \ab[20][53] , \ab[20][52] , \ab[20][51] , \ab[20][50] ,
         \ab[20][49] , \ab[20][48] , \ab[20][47] , \ab[20][46] , \ab[20][45] ,
         \ab[20][44] , \ab[20][43] , \ab[20][42] , \ab[20][41] , \ab[20][40] ,
         \ab[20][39] , \ab[20][38] , \ab[20][37] , \ab[20][36] , \ab[20][35] ,
         \ab[20][34] , \ab[20][33] , \ab[20][32] , \ab[20][31] , \ab[20][30] ,
         \ab[20][29] , \ab[20][28] , \ab[20][27] , \ab[20][26] , \ab[20][25] ,
         \ab[20][24] , \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] ,
         \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] ,
         \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] ,
         \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] ,
         \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] ,
         \ab[19][95] , \ab[19][94] , \ab[19][93] , \ab[19][92] , \ab[19][91] ,
         \ab[19][90] , \ab[19][89] , \ab[19][88] , \ab[19][87] , \ab[19][86] ,
         \ab[19][85] , \ab[19][84] , \ab[19][83] , \ab[19][82] , \ab[19][81] ,
         \ab[19][80] , \ab[19][79] , \ab[19][78] , \ab[19][77] , \ab[19][76] ,
         \ab[19][75] , \ab[19][74] , \ab[19][73] , \ab[19][72] , \ab[19][71] ,
         \ab[19][70] , \ab[19][69] , \ab[19][68] , \ab[19][67] , \ab[19][66] ,
         \ab[19][65] , \ab[19][64] , \ab[19][63] , \ab[19][62] , \ab[19][61] ,
         \ab[19][60] , \ab[19][59] , \ab[19][58] , \ab[19][57] , \ab[19][56] ,
         \ab[19][55] , \ab[19][54] , \ab[19][53] , \ab[19][52] , \ab[19][51] ,
         \ab[19][50] , \ab[19][49] , \ab[19][48] , \ab[19][47] , \ab[19][46] ,
         \ab[19][45] , \ab[19][44] , \ab[19][43] , \ab[19][42] , \ab[19][41] ,
         \ab[19][40] , \ab[19][39] , \ab[19][38] , \ab[19][37] , \ab[19][36] ,
         \ab[19][35] , \ab[19][34] , \ab[19][33] , \ab[19][32] , \ab[19][31] ,
         \ab[19][30] , \ab[19][29] , \ab[19][28] , \ab[19][27] , \ab[19][26] ,
         \ab[19][25] , \ab[19][24] , \ab[19][23] , \ab[19][22] , \ab[19][21] ,
         \ab[19][20] , \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] ,
         \ab[19][15] , \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] ,
         \ab[19][10] , \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] ,
         \ab[19][5] , \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] ,
         \ab[19][0] , \ab[18][95] , \ab[18][94] , \ab[18][93] , \ab[18][92] ,
         \ab[18][91] , \ab[18][90] , \ab[18][89] , \ab[18][88] , \ab[18][87] ,
         \ab[18][86] , \ab[18][85] , \ab[18][84] , \ab[18][83] , \ab[18][82] ,
         \ab[18][81] , \ab[18][80] , \ab[18][79] , \ab[18][78] , \ab[18][77] ,
         \ab[18][76] , \ab[18][75] , \ab[18][74] , \ab[18][73] , \ab[18][72] ,
         \ab[18][71] , \ab[18][70] , \ab[18][69] , \ab[18][68] , \ab[18][67] ,
         \ab[18][66] , \ab[18][65] , \ab[18][64] , \ab[18][63] , \ab[18][62] ,
         \ab[18][61] , \ab[18][60] , \ab[18][59] , \ab[18][58] , \ab[18][57] ,
         \ab[18][56] , \ab[18][55] , \ab[18][54] , \ab[18][53] , \ab[18][52] ,
         \ab[18][51] , \ab[18][50] , \ab[18][49] , \ab[18][48] , \ab[18][47] ,
         \ab[18][46] , \ab[18][45] , \ab[18][44] , \ab[18][43] , \ab[18][42] ,
         \ab[18][41] , \ab[18][40] , \ab[18][39] , \ab[18][38] , \ab[18][37] ,
         \ab[18][36] , \ab[18][35] , \ab[18][34] , \ab[18][33] , \ab[18][32] ,
         \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] , \ab[18][27] ,
         \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] , \ab[18][22] ,
         \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] , \ab[18][17] ,
         \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] , \ab[18][12] ,
         \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] , \ab[18][7] ,
         \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] , \ab[18][2] ,
         \ab[18][1] , \ab[18][0] , \ab[17][95] , \ab[17][94] , \ab[17][93] ,
         \ab[17][92] , \ab[17][91] , \ab[17][90] , \ab[17][89] , \ab[17][88] ,
         \ab[17][87] , \ab[17][86] , \ab[17][85] , \ab[17][84] , \ab[17][83] ,
         \ab[17][82] , \ab[17][81] , \ab[17][80] , \ab[17][79] , \ab[17][78] ,
         \ab[17][77] , \ab[17][76] , \ab[17][75] , \ab[17][74] , \ab[17][73] ,
         \ab[17][72] , \ab[17][71] , \ab[17][70] , \ab[17][69] , \ab[17][68] ,
         \ab[17][67] , \ab[17][66] , \ab[17][65] , \ab[17][64] , \ab[17][63] ,
         \ab[17][62] , \ab[17][61] , \ab[17][60] , \ab[17][59] , \ab[17][58] ,
         \ab[17][57] , \ab[17][56] , \ab[17][55] , \ab[17][54] , \ab[17][53] ,
         \ab[17][52] , \ab[17][51] , \ab[17][50] , \ab[17][49] , \ab[17][48] ,
         \ab[17][47] , \ab[17][46] , \ab[17][45] , \ab[17][44] , \ab[17][43] ,
         \ab[17][42] , \ab[17][41] , \ab[17][40] , \ab[17][39] , \ab[17][38] ,
         \ab[17][37] , \ab[17][36] , \ab[17][35] , \ab[17][34] , \ab[17][33] ,
         \ab[17][32] , \ab[17][31] , \ab[17][30] , \ab[17][29] , \ab[17][28] ,
         \ab[17][27] , \ab[17][26] , \ab[17][25] , \ab[17][24] , \ab[17][23] ,
         \ab[17][22] , \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] ,
         \ab[17][17] , \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] ,
         \ab[17][12] , \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] ,
         \ab[17][7] , \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] ,
         \ab[17][2] , \ab[17][1] , \ab[17][0] , \ab[16][95] , \ab[16][94] ,
         \ab[16][93] , \ab[16][92] , \ab[16][91] , \ab[16][90] , \ab[16][89] ,
         \ab[16][88] , \ab[16][87] , \ab[16][86] , \ab[16][85] , \ab[16][84] ,
         \ab[16][83] , \ab[16][82] , \ab[16][81] , \ab[16][80] , \ab[16][79] ,
         \ab[16][78] , \ab[16][77] , \ab[16][76] , \ab[16][75] , \ab[16][74] ,
         \ab[16][73] , \ab[16][72] , \ab[16][71] , \ab[16][70] , \ab[16][69] ,
         \ab[16][68] , \ab[16][67] , \ab[16][66] , \ab[16][65] , \ab[16][64] ,
         \ab[16][63] , \ab[16][62] , \ab[16][61] , \ab[16][60] , \ab[16][59] ,
         \ab[16][58] , \ab[16][57] , \ab[16][56] , \ab[16][55] , \ab[16][54] ,
         \ab[16][53] , \ab[16][52] , \ab[16][51] , \ab[16][50] , \ab[16][49] ,
         \ab[16][48] , \ab[16][47] , \ab[16][46] , \ab[16][45] , \ab[16][44] ,
         \ab[16][43] , \ab[16][42] , \ab[16][41] , \ab[16][40] , \ab[16][39] ,
         \ab[16][38] , \ab[16][37] , \ab[16][36] , \ab[16][35] , \ab[16][34] ,
         \ab[16][33] , \ab[16][32] , \ab[16][31] , \ab[16][30] , \ab[16][29] ,
         \ab[16][28] , \ab[16][27] , \ab[16][26] , \ab[16][25] , \ab[16][24] ,
         \ab[16][23] , \ab[16][22] , \ab[16][21] , \ab[16][20] , \ab[16][19] ,
         \ab[16][18] , \ab[16][17] , \ab[16][16] , \ab[16][15] , \ab[16][14] ,
         \ab[16][13] , \ab[16][12] , \ab[16][11] , \ab[16][10] , \ab[16][9] ,
         \ab[16][8] , \ab[16][7] , \ab[16][6] , \ab[16][5] , \ab[16][4] ,
         \ab[16][3] , \ab[16][2] , \ab[16][1] , \ab[16][0] , \ab[15][95] ,
         \ab[15][94] , \ab[15][93] , \ab[15][92] , \ab[15][91] , \ab[15][90] ,
         \ab[15][89] , \ab[15][88] , \ab[15][87] , \ab[15][86] , \ab[15][85] ,
         \ab[15][84] , \ab[15][83] , \ab[15][82] , \ab[15][81] , \ab[15][80] ,
         \ab[15][79] , \ab[15][78] , \ab[15][77] , \ab[15][76] , \ab[15][75] ,
         \ab[15][74] , \ab[15][73] , \ab[15][72] , \ab[15][71] , \ab[15][70] ,
         \ab[15][69] , \ab[15][68] , \ab[15][67] , \ab[15][66] , \ab[15][65] ,
         \ab[15][64] , \ab[15][63] , \ab[15][62] , \ab[15][61] , \ab[15][60] ,
         \ab[15][59] , \ab[15][58] , \ab[15][57] , \ab[15][56] , \ab[15][55] ,
         \ab[15][54] , \ab[15][53] , \ab[15][52] , \ab[15][51] , \ab[15][50] ,
         \ab[15][49] , \ab[15][48] , \ab[15][47] , \ab[15][46] , \ab[15][45] ,
         \ab[15][44] , \ab[15][43] , \ab[15][42] , \ab[15][41] , \ab[15][40] ,
         \ab[15][39] , \ab[15][38] , \ab[15][37] , \ab[15][36] , \ab[15][35] ,
         \ab[15][34] , \ab[15][33] , \ab[15][32] , \ab[15][31] , \ab[15][30] ,
         \ab[15][29] , \ab[15][28] , \ab[15][27] , \ab[15][26] , \ab[15][25] ,
         \ab[15][24] , \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] ,
         \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] ,
         \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] ,
         \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] ,
         \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] ,
         \ab[14][95] , \ab[14][94] , \ab[14][93] , \ab[14][92] , \ab[14][91] ,
         \ab[14][90] , \ab[14][89] , \ab[14][88] , \ab[14][87] , \ab[14][86] ,
         \ab[14][85] , \ab[14][84] , \ab[14][83] , \ab[14][82] , \ab[14][81] ,
         \ab[14][80] , \ab[14][79] , \ab[14][78] , \ab[14][77] , \ab[14][76] ,
         \ab[14][75] , \ab[14][74] , \ab[14][73] , \ab[14][72] , \ab[14][71] ,
         \ab[14][70] , \ab[14][69] , \ab[14][68] , \ab[14][67] , \ab[14][66] ,
         \ab[14][65] , \ab[14][64] , \ab[14][63] , \ab[14][62] , \ab[14][61] ,
         \ab[14][60] , \ab[14][59] , \ab[14][58] , \ab[14][57] , \ab[14][56] ,
         \ab[14][55] , \ab[14][54] , \ab[14][53] , \ab[14][52] , \ab[14][51] ,
         \ab[14][50] , \ab[14][49] , \ab[14][48] , \ab[14][47] , \ab[14][46] ,
         \ab[14][45] , \ab[14][44] , \ab[14][43] , \ab[14][42] , \ab[14][41] ,
         \ab[14][40] , \ab[14][39] , \ab[14][38] , \ab[14][37] , \ab[14][36] ,
         \ab[14][35] , \ab[14][34] , \ab[14][33] , \ab[14][32] , \ab[14][31] ,
         \ab[14][30] , \ab[14][29] , \ab[14][28] , \ab[14][27] , \ab[14][26] ,
         \ab[14][25] , \ab[14][24] , \ab[14][23] , \ab[14][22] , \ab[14][21] ,
         \ab[14][20] , \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] ,
         \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] ,
         \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] ,
         \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] ,
         \ab[14][0] , \ab[13][95] , \ab[13][94] , \ab[13][93] , \ab[13][92] ,
         \ab[13][91] , \ab[13][90] , \ab[13][89] , \ab[13][88] , \ab[13][87] ,
         \ab[13][86] , \ab[13][85] , \ab[13][84] , \ab[13][83] , \ab[13][82] ,
         \ab[13][81] , \ab[13][80] , \ab[13][79] , \ab[13][78] , \ab[13][77] ,
         \ab[13][76] , \ab[13][75] , \ab[13][74] , \ab[13][73] , \ab[13][72] ,
         \ab[13][71] , \ab[13][70] , \ab[13][69] , \ab[13][68] , \ab[13][67] ,
         \ab[13][66] , \ab[13][65] , \ab[13][64] , \ab[13][63] , \ab[13][62] ,
         \ab[13][61] , \ab[13][60] , \ab[13][59] , \ab[13][58] , \ab[13][57] ,
         \ab[13][56] , \ab[13][55] , \ab[13][54] , \ab[13][53] , \ab[13][52] ,
         \ab[13][51] , \ab[13][50] , \ab[13][49] , \ab[13][48] , \ab[13][47] ,
         \ab[13][46] , \ab[13][45] , \ab[13][44] , \ab[13][43] , \ab[13][42] ,
         \ab[13][41] , \ab[13][40] , \ab[13][39] , \ab[13][38] , \ab[13][37] ,
         \ab[13][36] , \ab[13][35] , \ab[13][34] , \ab[13][33] , \ab[13][32] ,
         \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] , \ab[13][27] ,
         \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] , \ab[13][22] ,
         \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] , \ab[13][17] ,
         \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] , \ab[13][12] ,
         \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] , \ab[13][7] ,
         \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] , \ab[13][2] ,
         \ab[13][1] , \ab[13][0] , \ab[12][95] , \ab[12][94] , \ab[12][93] ,
         \ab[12][92] , \ab[12][91] , \ab[12][90] , \ab[12][89] , \ab[12][88] ,
         \ab[12][87] , \ab[12][86] , \ab[12][85] , \ab[12][84] , \ab[12][83] ,
         \ab[12][82] , \ab[12][81] , \ab[12][80] , \ab[12][79] , \ab[12][78] ,
         \ab[12][77] , \ab[12][76] , \ab[12][75] , \ab[12][74] , \ab[12][73] ,
         \ab[12][72] , \ab[12][71] , \ab[12][70] , \ab[12][69] , \ab[12][68] ,
         \ab[12][67] , \ab[12][66] , \ab[12][65] , \ab[12][64] , \ab[12][63] ,
         \ab[12][62] , \ab[12][61] , \ab[12][60] , \ab[12][59] , \ab[12][58] ,
         \ab[12][57] , \ab[12][56] , \ab[12][55] , \ab[12][54] , \ab[12][53] ,
         \ab[12][52] , \ab[12][51] , \ab[12][50] , \ab[12][49] , \ab[12][48] ,
         \ab[12][47] , \ab[12][46] , \ab[12][45] , \ab[12][44] , \ab[12][43] ,
         \ab[12][42] , \ab[12][41] , \ab[12][40] , \ab[12][39] , \ab[12][38] ,
         \ab[12][37] , \ab[12][36] , \ab[12][35] , \ab[12][34] , \ab[12][33] ,
         \ab[12][32] , \ab[12][31] , \ab[12][30] , \ab[12][29] , \ab[12][28] ,
         \ab[12][27] , \ab[12][26] , \ab[12][25] , \ab[12][24] , \ab[12][23] ,
         \ab[12][22] , \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] ,
         \ab[12][17] , \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] ,
         \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] ,
         \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] ,
         \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][95] , \ab[11][94] ,
         \ab[11][93] , \ab[11][92] , \ab[11][91] , \ab[11][90] , \ab[11][89] ,
         \ab[11][88] , \ab[11][87] , \ab[11][86] , \ab[11][85] , \ab[11][84] ,
         \ab[11][83] , \ab[11][82] , \ab[11][81] , \ab[11][80] , \ab[11][79] ,
         \ab[11][78] , \ab[11][77] , \ab[11][76] , \ab[11][75] , \ab[11][74] ,
         \ab[11][73] , \ab[11][72] , \ab[11][71] , \ab[11][70] , \ab[11][69] ,
         \ab[11][68] , \ab[11][67] , \ab[11][66] , \ab[11][65] , \ab[11][64] ,
         \ab[11][63] , \ab[11][62] , \ab[11][61] , \ab[11][60] , \ab[11][59] ,
         \ab[11][58] , \ab[11][57] , \ab[11][56] , \ab[11][55] , \ab[11][54] ,
         \ab[11][53] , \ab[11][52] , \ab[11][51] , \ab[11][50] , \ab[11][49] ,
         \ab[11][48] , \ab[11][47] , \ab[11][46] , \ab[11][45] , \ab[11][44] ,
         \ab[11][43] , \ab[11][42] , \ab[11][41] , \ab[11][40] , \ab[11][39] ,
         \ab[11][38] , \ab[11][37] , \ab[11][36] , \ab[11][35] , \ab[11][34] ,
         \ab[11][33] , \ab[11][32] , \ab[11][31] , \ab[11][30] , \ab[11][29] ,
         \ab[11][28] , \ab[11][27] , \ab[11][26] , \ab[11][25] , \ab[11][24] ,
         \ab[11][23] , \ab[11][22] , \ab[11][21] , \ab[11][20] , \ab[11][19] ,
         \ab[11][18] , \ab[11][17] , \ab[11][16] , \ab[11][15] , \ab[11][14] ,
         \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][95] ,
         \ab[10][94] , \ab[10][93] , \ab[10][92] , \ab[10][91] , \ab[10][90] ,
         \ab[10][89] , \ab[10][88] , \ab[10][87] , \ab[10][86] , \ab[10][85] ,
         \ab[10][84] , \ab[10][83] , \ab[10][82] , \ab[10][81] , \ab[10][80] ,
         \ab[10][79] , \ab[10][78] , \ab[10][77] , \ab[10][76] , \ab[10][75] ,
         \ab[10][74] , \ab[10][73] , \ab[10][72] , \ab[10][71] , \ab[10][70] ,
         \ab[10][69] , \ab[10][68] , \ab[10][67] , \ab[10][66] , \ab[10][65] ,
         \ab[10][64] , \ab[10][63] , \ab[10][62] , \ab[10][61] , \ab[10][60] ,
         \ab[10][59] , \ab[10][58] , \ab[10][57] , \ab[10][56] , \ab[10][55] ,
         \ab[10][54] , \ab[10][53] , \ab[10][52] , \ab[10][51] , \ab[10][50] ,
         \ab[10][49] , \ab[10][48] , \ab[10][47] , \ab[10][46] , \ab[10][45] ,
         \ab[10][44] , \ab[10][43] , \ab[10][42] , \ab[10][41] , \ab[10][40] ,
         \ab[10][39] , \ab[10][38] , \ab[10][37] , \ab[10][36] , \ab[10][35] ,
         \ab[10][34] , \ab[10][33] , \ab[10][32] , \ab[10][31] , \ab[10][30] ,
         \ab[10][29] , \ab[10][28] , \ab[10][27] , \ab[10][26] , \ab[10][25] ,
         \ab[10][24] , \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] ,
         \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][95] , \ab[9][94] , \ab[9][93] , \ab[9][92] , \ab[9][91] ,
         \ab[9][90] , \ab[9][89] , \ab[9][88] , \ab[9][87] , \ab[9][86] ,
         \ab[9][85] , \ab[9][84] , \ab[9][83] , \ab[9][82] , \ab[9][81] ,
         \ab[9][80] , \ab[9][79] , \ab[9][78] , \ab[9][77] , \ab[9][76] ,
         \ab[9][75] , \ab[9][74] , \ab[9][73] , \ab[9][72] , \ab[9][71] ,
         \ab[9][70] , \ab[9][69] , \ab[9][68] , \ab[9][67] , \ab[9][66] ,
         \ab[9][65] , \ab[9][64] , \ab[9][63] , \ab[9][62] , \ab[9][61] ,
         \ab[9][60] , \ab[9][59] , \ab[9][58] , \ab[9][57] , \ab[9][56] ,
         \ab[9][55] , \ab[9][54] , \ab[9][53] , \ab[9][52] , \ab[9][51] ,
         \ab[9][50] , \ab[9][49] , \ab[9][48] , \ab[9][47] , \ab[9][46] ,
         \ab[9][45] , \ab[9][44] , \ab[9][43] , \ab[9][42] , \ab[9][41] ,
         \ab[9][40] , \ab[9][39] , \ab[9][38] , \ab[9][37] , \ab[9][36] ,
         \ab[9][35] , \ab[9][34] , \ab[9][33] , \ab[9][32] , \ab[9][31] ,
         \ab[9][30] , \ab[9][29] , \ab[9][28] , \ab[9][27] , \ab[9][26] ,
         \ab[9][25] , \ab[9][24] , \ab[9][23] , \ab[9][22] , \ab[9][21] ,
         \ab[9][20] , \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] ,
         \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] ,
         \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] ,
         \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] ,
         \ab[9][0] , \ab[8][95] , \ab[8][94] , \ab[8][93] , \ab[8][92] ,
         \ab[8][91] , \ab[8][90] , \ab[8][89] , \ab[8][88] , \ab[8][87] ,
         \ab[8][86] , \ab[8][85] , \ab[8][84] , \ab[8][83] , \ab[8][82] ,
         \ab[8][81] , \ab[8][80] , \ab[8][79] , \ab[8][78] , \ab[8][77] ,
         \ab[8][76] , \ab[8][75] , \ab[8][74] , \ab[8][73] , \ab[8][72] ,
         \ab[8][71] , \ab[8][70] , \ab[8][69] , \ab[8][68] , \ab[8][67] ,
         \ab[8][66] , \ab[8][65] , \ab[8][64] , \ab[8][63] , \ab[8][62] ,
         \ab[8][61] , \ab[8][60] , \ab[8][59] , \ab[8][58] , \ab[8][57] ,
         \ab[8][56] , \ab[8][55] , \ab[8][54] , \ab[8][53] , \ab[8][52] ,
         \ab[8][51] , \ab[8][50] , \ab[8][49] , \ab[8][48] , \ab[8][47] ,
         \ab[8][46] , \ab[8][45] , \ab[8][44] , \ab[8][43] , \ab[8][42] ,
         \ab[8][41] , \ab[8][40] , \ab[8][39] , \ab[8][38] , \ab[8][37] ,
         \ab[8][36] , \ab[8][35] , \ab[8][34] , \ab[8][33] , \ab[8][32] ,
         \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] , \ab[8][27] ,
         \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] , \ab[8][22] ,
         \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] , \ab[8][17] ,
         \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] , \ab[8][12] ,
         \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] ,
         \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] ,
         \ab[8][1] , \ab[8][0] , \ab[7][95] , \ab[7][94] , \ab[7][93] ,
         \ab[7][92] , \ab[7][91] , \ab[7][90] , \ab[7][89] , \ab[7][88] ,
         \ab[7][87] , \ab[7][86] , \ab[7][85] , \ab[7][84] , \ab[7][83] ,
         \ab[7][82] , \ab[7][81] , \ab[7][80] , \ab[7][79] , \ab[7][78] ,
         \ab[7][77] , \ab[7][76] , \ab[7][75] , \ab[7][74] , \ab[7][73] ,
         \ab[7][72] , \ab[7][71] , \ab[7][70] , \ab[7][69] , \ab[7][68] ,
         \ab[7][67] , \ab[7][66] , \ab[7][65] , \ab[7][64] , \ab[7][63] ,
         \ab[7][62] , \ab[7][61] , \ab[7][60] , \ab[7][59] , \ab[7][58] ,
         \ab[7][57] , \ab[7][56] , \ab[7][55] , \ab[7][54] , \ab[7][53] ,
         \ab[7][52] , \ab[7][51] , \ab[7][50] , \ab[7][49] , \ab[7][48] ,
         \ab[7][47] , \ab[7][46] , \ab[7][45] , \ab[7][44] , \ab[7][43] ,
         \ab[7][42] , \ab[7][41] , \ab[7][40] , \ab[7][39] , \ab[7][38] ,
         \ab[7][37] , \ab[7][36] , \ab[7][35] , \ab[7][34] , \ab[7][33] ,
         \ab[7][32] , \ab[7][31] , \ab[7][30] , \ab[7][29] , \ab[7][28] ,
         \ab[7][27] , \ab[7][26] , \ab[7][25] , \ab[7][24] , \ab[7][23] ,
         \ab[7][22] , \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] ,
         \ab[7][17] , \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] ,
         \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] ,
         \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][95] , \ab[6][94] ,
         \ab[6][93] , \ab[6][92] , \ab[6][91] , \ab[6][90] , \ab[6][89] ,
         \ab[6][88] , \ab[6][87] , \ab[6][86] , \ab[6][85] , \ab[6][84] ,
         \ab[6][83] , \ab[6][82] , \ab[6][81] , \ab[6][80] , \ab[6][79] ,
         \ab[6][78] , \ab[6][77] , \ab[6][76] , \ab[6][75] , \ab[6][74] ,
         \ab[6][73] , \ab[6][72] , \ab[6][71] , \ab[6][70] , \ab[6][69] ,
         \ab[6][68] , \ab[6][67] , \ab[6][66] , \ab[6][65] , \ab[6][64] ,
         \ab[6][63] , \ab[6][62] , \ab[6][61] , \ab[6][60] , \ab[6][59] ,
         \ab[6][58] , \ab[6][57] , \ab[6][56] , \ab[6][55] , \ab[6][54] ,
         \ab[6][53] , \ab[6][52] , \ab[6][51] , \ab[6][50] , \ab[6][49] ,
         \ab[6][48] , \ab[6][47] , \ab[6][46] , \ab[6][45] , \ab[6][44] ,
         \ab[6][43] , \ab[6][42] , \ab[6][41] , \ab[6][40] , \ab[6][39] ,
         \ab[6][38] , \ab[6][37] , \ab[6][36] , \ab[6][35] , \ab[6][34] ,
         \ab[6][33] , \ab[6][32] , \ab[6][31] , \ab[6][30] , \ab[6][29] ,
         \ab[6][28] , \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] ,
         \ab[6][23] , \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] ,
         \ab[6][18] , \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][95] ,
         \ab[5][94] , \ab[5][93] , \ab[5][92] , \ab[5][91] , \ab[5][90] ,
         \ab[5][89] , \ab[5][88] , \ab[5][87] , \ab[5][86] , \ab[5][85] ,
         \ab[5][84] , \ab[5][83] , \ab[5][82] , \ab[5][81] , \ab[5][80] ,
         \ab[5][79] , \ab[5][78] , \ab[5][77] , \ab[5][76] , \ab[5][75] ,
         \ab[5][74] , \ab[5][73] , \ab[5][72] , \ab[5][71] , \ab[5][70] ,
         \ab[5][69] , \ab[5][68] , \ab[5][67] , \ab[5][66] , \ab[5][65] ,
         \ab[5][64] , \ab[5][63] , \ab[5][62] , \ab[5][61] , \ab[5][60] ,
         \ab[5][59] , \ab[5][58] , \ab[5][57] , \ab[5][56] , \ab[5][55] ,
         \ab[5][54] , \ab[5][53] , \ab[5][52] , \ab[5][51] , \ab[5][50] ,
         \ab[5][49] , \ab[5][48] , \ab[5][47] , \ab[5][46] , \ab[5][45] ,
         \ab[5][44] , \ab[5][43] , \ab[5][42] , \ab[5][41] , \ab[5][40] ,
         \ab[5][39] , \ab[5][38] , \ab[5][37] , \ab[5][36] , \ab[5][35] ,
         \ab[5][34] , \ab[5][33] , \ab[5][32] , \ab[5][31] , \ab[5][30] ,
         \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] , \ab[5][25] ,
         \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] ,
         \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][95] , \ab[4][94] , \ab[4][93] , \ab[4][92] , \ab[4][91] ,
         \ab[4][90] , \ab[4][89] , \ab[4][88] , \ab[4][87] , \ab[4][86] ,
         \ab[4][85] , \ab[4][84] , \ab[4][83] , \ab[4][82] , \ab[4][81] ,
         \ab[4][80] , \ab[4][79] , \ab[4][78] , \ab[4][77] , \ab[4][76] ,
         \ab[4][75] , \ab[4][74] , \ab[4][73] , \ab[4][72] , \ab[4][71] ,
         \ab[4][70] , \ab[4][69] , \ab[4][68] , \ab[4][67] , \ab[4][66] ,
         \ab[4][65] , \ab[4][64] , \ab[4][63] , \ab[4][62] , \ab[4][61] ,
         \ab[4][60] , \ab[4][59] , \ab[4][58] , \ab[4][57] , \ab[4][56] ,
         \ab[4][55] , \ab[4][54] , \ab[4][53] , \ab[4][52] , \ab[4][51] ,
         \ab[4][50] , \ab[4][49] , \ab[4][48] , \ab[4][47] , \ab[4][46] ,
         \ab[4][45] , \ab[4][44] , \ab[4][43] , \ab[4][42] , \ab[4][41] ,
         \ab[4][40] , \ab[4][39] , \ab[4][38] , \ab[4][37] , \ab[4][36] ,
         \ab[4][35] , \ab[4][34] , \ab[4][33] , \ab[4][32] , \ab[4][31] ,
         \ab[4][30] , \ab[4][29] , \ab[4][28] , \ab[4][27] , \ab[4][26] ,
         \ab[4][25] , \ab[4][24] , \ab[4][23] , \ab[4][22] , \ab[4][21] ,
         \ab[4][20] , \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] ,
         \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] ,
         \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] ,
         \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] ,
         \ab[4][0] , \ab[3][95] , \ab[3][94] , \ab[3][93] , \ab[3][92] ,
         \ab[3][91] , \ab[3][90] , \ab[3][89] , \ab[3][88] , \ab[3][87] ,
         \ab[3][86] , \ab[3][85] , \ab[3][84] , \ab[3][83] , \ab[3][82] ,
         \ab[3][81] , \ab[3][80] , \ab[3][79] , \ab[3][78] , \ab[3][77] ,
         \ab[3][76] , \ab[3][75] , \ab[3][74] , \ab[3][73] , \ab[3][72] ,
         \ab[3][71] , \ab[3][70] , \ab[3][69] , \ab[3][68] , \ab[3][67] ,
         \ab[3][66] , \ab[3][65] , \ab[3][64] , \ab[3][63] , \ab[3][62] ,
         \ab[3][61] , \ab[3][60] , \ab[3][59] , \ab[3][58] , \ab[3][57] ,
         \ab[3][56] , \ab[3][55] , \ab[3][54] , \ab[3][53] , \ab[3][52] ,
         \ab[3][51] , \ab[3][50] , \ab[3][49] , \ab[3][48] , \ab[3][47] ,
         \ab[3][46] , \ab[3][45] , \ab[3][44] , \ab[3][43] , \ab[3][42] ,
         \ab[3][41] , \ab[3][40] , \ab[3][39] , \ab[3][38] , \ab[3][37] ,
         \ab[3][36] , \ab[3][35] , \ab[3][34] , \ab[3][33] , \ab[3][32] ,
         \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] , \ab[3][27] ,
         \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] , \ab[3][22] ,
         \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] , \ab[3][17] ,
         \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] , \ab[3][12] ,
         \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] ,
         \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] ,
         \ab[3][1] , \ab[3][0] , \ab[2][95] , \ab[2][94] , \ab[2][93] ,
         \ab[2][92] , \ab[2][91] , \ab[2][90] , \ab[2][89] , \ab[2][88] ,
         \ab[2][87] , \ab[2][86] , \ab[2][85] , \ab[2][84] , \ab[2][83] ,
         \ab[2][82] , \ab[2][81] , \ab[2][80] , \ab[2][79] , \ab[2][78] ,
         \ab[2][77] , \ab[2][76] , \ab[2][75] , \ab[2][74] , \ab[2][73] ,
         \ab[2][72] , \ab[2][71] , \ab[2][70] , \ab[2][69] , \ab[2][68] ,
         \ab[2][67] , \ab[2][66] , \ab[2][65] , \ab[2][64] , \ab[2][63] ,
         \ab[2][62] , \ab[2][61] , \ab[2][60] , \ab[2][59] , \ab[2][58] ,
         \ab[2][57] , \ab[2][56] , \ab[2][55] , \ab[2][54] , \ab[2][53] ,
         \ab[2][52] , \ab[2][51] , \ab[2][50] , \ab[2][49] , \ab[2][48] ,
         \ab[2][47] , \ab[2][46] , \ab[2][45] , \ab[2][44] , \ab[2][43] ,
         \ab[2][42] , \ab[2][41] , \ab[2][40] , \ab[2][39] , \ab[2][38] ,
         \ab[2][37] , \ab[2][36] , \ab[2][35] , \ab[2][34] , \ab[2][33] ,
         \ab[2][32] , \ab[2][31] , \ab[2][30] , \ab[2][29] , \ab[2][28] ,
         \ab[2][27] , \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] ,
         \ab[2][22] , \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] ,
         \ab[2][17] , \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] ,
         \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][95] , \ab[1][94] ,
         \ab[1][93] , \ab[1][92] , \ab[1][91] , \ab[1][90] , \ab[1][89] ,
         \ab[1][88] , \ab[1][87] , \ab[1][86] , \ab[1][85] , \ab[1][84] ,
         \ab[1][83] , \ab[1][82] , \ab[1][81] , \ab[1][80] , \ab[1][79] ,
         \ab[1][78] , \ab[1][77] , \ab[1][76] , \ab[1][75] , \ab[1][74] ,
         \ab[1][73] , \ab[1][72] , \ab[1][71] , \ab[1][70] , \ab[1][69] ,
         \ab[1][68] , \ab[1][67] , \ab[1][66] , \ab[1][65] , \ab[1][64] ,
         \ab[1][63] , \ab[1][62] , \ab[1][61] , \ab[1][60] , \ab[1][59] ,
         \ab[1][58] , \ab[1][57] , \ab[1][56] , \ab[1][55] , \ab[1][54] ,
         \ab[1][53] , \ab[1][52] , \ab[1][51] , \ab[1][50] , \ab[1][49] ,
         \ab[1][48] , \ab[1][47] , \ab[1][46] , \ab[1][45] , \ab[1][44] ,
         \ab[1][43] , \ab[1][42] , \ab[1][41] , \ab[1][40] , \ab[1][39] ,
         \ab[1][38] , \ab[1][37] , \ab[1][36] , \ab[1][35] , \ab[1][34] ,
         \ab[1][33] , \ab[1][32] , \ab[1][31] , \ab[1][30] , \ab[1][29] ,
         \ab[1][28] , \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] ,
         \ab[1][23] , \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] ,
         \ab[1][18] , \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[0][95] , \ab[0][94] , \ab[0][93] ,
         \ab[0][92] , \ab[0][91] , \ab[0][90] , \ab[0][89] , \ab[0][88] ,
         \ab[0][87] , \ab[0][86] , \ab[0][85] , \ab[0][84] , \ab[0][83] ,
         \ab[0][82] , \ab[0][81] , \ab[0][80] , \ab[0][79] , \ab[0][78] ,
         \ab[0][77] , \ab[0][76] , \ab[0][75] , \ab[0][74] , \ab[0][73] ,
         \ab[0][72] , \ab[0][71] , \ab[0][70] , \ab[0][69] , \ab[0][68] ,
         \ab[0][67] , \ab[0][66] , \ab[0][65] , \ab[0][64] , \ab[0][63] ,
         \ab[0][62] , \ab[0][61] , \ab[0][60] , \ab[0][59] , \ab[0][58] ,
         \ab[0][57] , \ab[0][56] , \ab[0][55] , \ab[0][54] , \ab[0][53] ,
         \ab[0][52] , \ab[0][51] , \ab[0][50] , \ab[0][49] , \ab[0][48] ,
         \ab[0][47] , \ab[0][46] , \ab[0][45] , \ab[0][44] , \ab[0][43] ,
         \ab[0][42] , \ab[0][41] , \ab[0][40] , \ab[0][39] , \ab[0][38] ,
         \ab[0][37] , \ab[0][36] , \ab[0][35] , \ab[0][34] , \ab[0][33] ,
         \ab[0][32] , \ab[0][31] , \ab[0][30] , \ab[0][29] , \ab[0][28] ,
         \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] , \ab[0][23] ,
         \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] , \ab[0][18] ,
         \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] , \ab[0][13] ,
         \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] , \ab[0][8] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \CARRYB[3][31] , \CARRYB[3][30] , \CARRYB[3][29] ,
         \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] ,
         \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] ,
         \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] ,
         \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][94] , \CARRYB[2][93] , \CARRYB[2][92] ,
         \CARRYB[2][91] , \CARRYB[2][90] , \CARRYB[2][89] , \CARRYB[2][88] ,
         \CARRYB[2][87] , \CARRYB[2][86] , \CARRYB[2][85] , \CARRYB[2][84] ,
         \CARRYB[2][83] , \CARRYB[2][82] , \CARRYB[2][81] , \CARRYB[2][80] ,
         \CARRYB[2][79] , \CARRYB[2][78] , \CARRYB[2][77] , \CARRYB[2][76] ,
         \CARRYB[2][75] , \CARRYB[2][74] , \CARRYB[2][73] , \CARRYB[2][72] ,
         \CARRYB[2][71] , \CARRYB[2][70] , \CARRYB[2][69] , \CARRYB[2][68] ,
         \CARRYB[2][67] , \CARRYB[2][66] , \CARRYB[2][65] , \CARRYB[2][64] ,
         \CARRYB[2][63] , \CARRYB[2][62] , \CARRYB[2][61] , \CARRYB[2][60] ,
         \CARRYB[2][59] , \CARRYB[2][58] , \CARRYB[2][57] , \CARRYB[2][56] ,
         \CARRYB[2][55] , \CARRYB[2][54] , \CARRYB[2][53] , \CARRYB[2][52] ,
         \CARRYB[2][51] , \CARRYB[2][50] , \CARRYB[2][49] , \CARRYB[2][48] ,
         \CARRYB[2][47] , \CARRYB[2][46] , \CARRYB[2][45] , \CARRYB[2][44] ,
         \CARRYB[2][43] , \CARRYB[2][42] , \CARRYB[2][41] , \CARRYB[2][40] ,
         \CARRYB[2][39] , \CARRYB[2][38] , \CARRYB[2][37] , \CARRYB[2][36] ,
         \CARRYB[2][35] , \CARRYB[2][34] , \CARRYB[2][33] , \CARRYB[2][32] ,
         \CARRYB[2][31] , \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] ,
         \CARRYB[2][27] , \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] ,
         \CARRYB[2][23] , \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] ,
         \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] ,
         \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[1][94] , \CARRYB[1][93] , \CARRYB[1][92] , \CARRYB[1][91] ,
         \CARRYB[1][90] , \CARRYB[1][89] , \CARRYB[1][88] , \CARRYB[1][87] ,
         \CARRYB[1][86] , \CARRYB[1][85] , \CARRYB[1][84] , \CARRYB[1][83] ,
         \CARRYB[1][82] , \CARRYB[1][81] , \CARRYB[1][80] , \CARRYB[1][79] ,
         \CARRYB[1][78] , \CARRYB[1][77] , \CARRYB[1][76] , \CARRYB[1][75] ,
         \CARRYB[1][74] , \CARRYB[1][73] , \CARRYB[1][72] , \CARRYB[1][71] ,
         \CARRYB[1][70] , \CARRYB[1][69] , \CARRYB[1][68] , \CARRYB[1][67] ,
         \CARRYB[1][66] , \CARRYB[1][65] , \CARRYB[1][64] , \CARRYB[1][63] ,
         \CARRYB[1][62] , \CARRYB[1][61] , \CARRYB[1][60] , \CARRYB[1][59] ,
         \CARRYB[1][58] , \CARRYB[1][57] , \CARRYB[1][56] , \CARRYB[1][55] ,
         \CARRYB[1][54] , \CARRYB[1][53] , \CARRYB[1][52] , \CARRYB[1][51] ,
         \CARRYB[1][50] , \CARRYB[1][49] , \CARRYB[1][48] , \CARRYB[1][47] ,
         \CARRYB[1][46] , \CARRYB[1][45] , \CARRYB[1][44] , \CARRYB[1][43] ,
         \CARRYB[1][42] , \CARRYB[1][41] , \CARRYB[1][40] , \CARRYB[1][39] ,
         \CARRYB[1][38] , \CARRYB[1][37] , \CARRYB[1][36] , \CARRYB[1][35] ,
         \CARRYB[1][34] , \CARRYB[1][33] , \CARRYB[1][32] , \CARRYB[1][31] ,
         \CARRYB[1][30] , \CARRYB[1][29] , \CARRYB[1][28] , \CARRYB[1][27] ,
         \CARRYB[1][26] , \CARRYB[1][25] , \CARRYB[1][24] , \CARRYB[1][23] ,
         \CARRYB[1][22] , \CARRYB[1][21] , \CARRYB[1][20] , \CARRYB[1][19] ,
         \CARRYB[1][18] , \CARRYB[1][17] , \CARRYB[1][16] , \CARRYB[1][15] ,
         \CARRYB[1][14] , \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] ,
         \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] ,
         \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[3][31] ,
         \SUMB[3][30] , \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] ,
         \SUMB[3][26] , \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] ,
         \SUMB[3][22] , \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] ,
         \SUMB[3][18] , \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] ,
         \SUMB[3][14] , \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] ,
         \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \SUMB[2][94] , \SUMB[2][93] , \SUMB[2][92] , \SUMB[2][91] ,
         \SUMB[2][90] , \SUMB[2][89] , \SUMB[2][88] , \SUMB[2][87] ,
         \SUMB[2][86] , \SUMB[2][85] , \SUMB[2][84] , \SUMB[2][83] ,
         \SUMB[2][82] , \SUMB[2][81] , \SUMB[2][80] , \SUMB[2][79] ,
         \SUMB[2][78] , \SUMB[2][77] , \SUMB[2][76] , \SUMB[2][75] ,
         \SUMB[2][74] , \SUMB[2][73] , \SUMB[2][72] , \SUMB[2][71] ,
         \SUMB[2][70] , \SUMB[2][69] , \SUMB[2][68] , \SUMB[2][67] ,
         \SUMB[2][66] , \SUMB[2][65] , \SUMB[2][64] , \SUMB[2][63] ,
         \SUMB[2][62] , \SUMB[2][61] , \SUMB[2][60] , \SUMB[2][59] ,
         \SUMB[2][58] , \SUMB[2][57] , \SUMB[2][56] , \SUMB[2][55] ,
         \SUMB[2][54] , \SUMB[2][53] , \SUMB[2][52] , \SUMB[2][51] ,
         \SUMB[2][50] , \SUMB[2][49] , \SUMB[2][48] , \SUMB[2][47] ,
         \SUMB[2][46] , \SUMB[2][45] , \SUMB[2][44] , \SUMB[2][43] ,
         \SUMB[2][42] , \SUMB[2][41] , \SUMB[2][40] , \SUMB[2][39] ,
         \SUMB[2][38] , \SUMB[2][37] , \SUMB[2][36] , \SUMB[2][35] ,
         \SUMB[2][34] , \SUMB[2][33] , \SUMB[2][32] , \SUMB[2][31] ,
         \SUMB[2][30] , \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] ,
         \SUMB[2][26] , \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] ,
         \SUMB[2][22] , \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] ,
         \SUMB[2][18] , \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][94] , \SUMB[1][93] , \SUMB[1][92] , \SUMB[1][91] ,
         \SUMB[1][90] , \SUMB[1][89] , \SUMB[1][88] , \SUMB[1][87] ,
         \SUMB[1][86] , \SUMB[1][85] , \SUMB[1][84] , \SUMB[1][83] ,
         \SUMB[1][82] , \SUMB[1][81] , \SUMB[1][80] , \SUMB[1][79] ,
         \SUMB[1][78] , \SUMB[1][77] , \SUMB[1][76] , \SUMB[1][75] ,
         \SUMB[1][74] , \SUMB[1][73] , \SUMB[1][72] , \SUMB[1][71] ,
         \SUMB[1][70] , \SUMB[1][69] , \SUMB[1][68] , \SUMB[1][67] ,
         \SUMB[1][66] , \SUMB[1][65] , \SUMB[1][64] , \SUMB[1][63] ,
         \SUMB[1][62] , \SUMB[1][61] , \SUMB[1][60] , \SUMB[1][59] ,
         \SUMB[1][58] , \SUMB[1][57] , \SUMB[1][56] , \SUMB[1][55] ,
         \SUMB[1][54] , \SUMB[1][53] , \SUMB[1][52] , \SUMB[1][51] ,
         \SUMB[1][50] , \SUMB[1][49] , \SUMB[1][48] , \SUMB[1][47] ,
         \SUMB[1][46] , \SUMB[1][45] , \SUMB[1][44] , \SUMB[1][43] ,
         \SUMB[1][42] , \SUMB[1][41] , \SUMB[1][40] , \SUMB[1][39] ,
         \SUMB[1][38] , \SUMB[1][37] , \SUMB[1][36] , \SUMB[1][35] ,
         \SUMB[1][34] , \SUMB[1][33] , \SUMB[1][32] , \SUMB[1][31] ,
         \SUMB[1][30] , \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] ,
         \SUMB[1][26] , \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] ,
         \SUMB[1][22] , \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] ,
         \SUMB[1][18] , \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] ,
         \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[8][63] , \CARRYB[8][62] , \CARRYB[8][61] , \CARRYB[8][60] ,
         \CARRYB[8][59] , \CARRYB[8][58] , \CARRYB[8][57] , \CARRYB[8][56] ,
         \CARRYB[8][55] , \CARRYB[8][54] , \CARRYB[8][53] , \CARRYB[8][52] ,
         \CARRYB[8][51] , \CARRYB[8][50] , \CARRYB[8][49] , \CARRYB[8][48] ,
         \CARRYB[8][47] , \CARRYB[8][46] , \CARRYB[8][45] , \CARRYB[8][44] ,
         \CARRYB[8][43] , \CARRYB[8][42] , \CARRYB[8][41] , \CARRYB[8][40] ,
         \CARRYB[8][39] , \CARRYB[8][38] , \CARRYB[8][37] , \CARRYB[8][36] ,
         \CARRYB[8][35] , \CARRYB[8][34] , \CARRYB[8][33] , \CARRYB[8][32] ,
         \CARRYB[8][31] , \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] ,
         \CARRYB[8][27] , \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] ,
         \CARRYB[8][23] , \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] ,
         \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] ,
         \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][94] , \CARRYB[7][93] , \CARRYB[7][92] , \CARRYB[7][91] ,
         \CARRYB[7][90] , \CARRYB[7][89] , \CARRYB[7][88] , \CARRYB[7][87] ,
         \CARRYB[7][86] , \CARRYB[7][85] , \CARRYB[7][84] , \CARRYB[7][83] ,
         \CARRYB[7][82] , \CARRYB[7][81] , \CARRYB[7][80] , \CARRYB[7][79] ,
         \CARRYB[7][78] , \CARRYB[7][77] , \CARRYB[7][76] , \CARRYB[7][75] ,
         \CARRYB[7][74] , \CARRYB[7][73] , \CARRYB[7][72] , \CARRYB[7][71] ,
         \CARRYB[7][70] , \CARRYB[7][69] , \CARRYB[7][68] , \CARRYB[7][67] ,
         \CARRYB[7][66] , \CARRYB[7][65] , \CARRYB[7][64] , \CARRYB[7][63] ,
         \CARRYB[7][62] , \CARRYB[7][61] , \CARRYB[7][60] , \CARRYB[7][59] ,
         \CARRYB[7][58] , \CARRYB[7][57] , \CARRYB[7][56] , \CARRYB[7][55] ,
         \CARRYB[7][54] , \CARRYB[7][53] , \CARRYB[7][52] , \CARRYB[7][51] ,
         \CARRYB[7][50] , \CARRYB[7][49] , \CARRYB[7][48] , \CARRYB[7][47] ,
         \CARRYB[7][46] , \CARRYB[7][45] , \CARRYB[7][44] , \CARRYB[7][43] ,
         \CARRYB[7][42] , \CARRYB[7][41] , \CARRYB[7][40] , \CARRYB[7][39] ,
         \CARRYB[7][38] , \CARRYB[7][37] , \CARRYB[7][36] , \CARRYB[7][35] ,
         \CARRYB[7][34] , \CARRYB[7][33] , \CARRYB[7][32] , \CARRYB[7][31] ,
         \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] ,
         \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] ,
         \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] ,
         \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] ,
         \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] ,
         \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] ,
         \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] ,
         \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][94] ,
         \CARRYB[6][93] , \CARRYB[6][92] , \CARRYB[6][91] , \CARRYB[6][90] ,
         \CARRYB[6][89] , \CARRYB[6][88] , \CARRYB[6][87] , \CARRYB[6][86] ,
         \CARRYB[6][85] , \CARRYB[6][84] , \CARRYB[6][83] , \CARRYB[6][82] ,
         \CARRYB[6][81] , \CARRYB[6][80] , \CARRYB[6][79] , \CARRYB[6][78] ,
         \CARRYB[6][77] , \CARRYB[6][76] , \CARRYB[6][75] , \CARRYB[6][74] ,
         \CARRYB[6][73] , \CARRYB[6][72] , \CARRYB[6][71] , \CARRYB[6][70] ,
         \CARRYB[6][69] , \CARRYB[6][68] , \CARRYB[6][67] , \CARRYB[6][66] ,
         \CARRYB[6][65] , \CARRYB[6][64] , \CARRYB[6][63] , \CARRYB[6][62] ,
         \CARRYB[6][61] , \CARRYB[6][60] , \CARRYB[6][59] , \CARRYB[6][58] ,
         \CARRYB[6][57] , \CARRYB[6][56] , \CARRYB[6][55] , \CARRYB[6][54] ,
         \CARRYB[6][53] , \CARRYB[6][52] , \CARRYB[6][51] , \CARRYB[6][50] ,
         \CARRYB[6][49] , \CARRYB[6][48] , \CARRYB[6][47] , \CARRYB[6][46] ,
         \CARRYB[6][45] , \CARRYB[6][44] , \CARRYB[6][43] , \CARRYB[6][42] ,
         \CARRYB[6][41] , \CARRYB[6][40] , \CARRYB[6][39] , \CARRYB[6][38] ,
         \CARRYB[6][37] , \CARRYB[6][36] , \CARRYB[6][35] , \CARRYB[6][34] ,
         \CARRYB[6][33] , \CARRYB[6][32] , \CARRYB[6][31] , \CARRYB[6][30] ,
         \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] ,
         \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] ,
         \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] ,
         \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] ,
         \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] ,
         \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][94] , \CARRYB[5][93] ,
         \CARRYB[5][92] , \CARRYB[5][91] , \CARRYB[5][90] , \CARRYB[5][89] ,
         \CARRYB[5][88] , \CARRYB[5][87] , \CARRYB[5][86] , \CARRYB[5][85] ,
         \CARRYB[5][84] , \CARRYB[5][83] , \CARRYB[5][82] , \CARRYB[5][81] ,
         \CARRYB[5][80] , \CARRYB[5][79] , \CARRYB[5][78] , \CARRYB[5][77] ,
         \CARRYB[5][76] , \CARRYB[5][75] , \CARRYB[5][74] , \CARRYB[5][73] ,
         \CARRYB[5][72] , \CARRYB[5][71] , \CARRYB[5][70] , \CARRYB[5][69] ,
         \CARRYB[5][68] , \CARRYB[5][67] , \CARRYB[5][66] , \CARRYB[5][65] ,
         \CARRYB[5][64] , \CARRYB[5][63] , \CARRYB[5][62] , \CARRYB[5][61] ,
         \CARRYB[5][60] , \CARRYB[5][59] , \CARRYB[5][58] , \CARRYB[5][57] ,
         \CARRYB[5][56] , \CARRYB[5][55] , \CARRYB[5][54] , \CARRYB[5][53] ,
         \CARRYB[5][52] , \CARRYB[5][51] , \CARRYB[5][50] , \CARRYB[5][49] ,
         \CARRYB[5][48] , \CARRYB[5][47] , \CARRYB[5][46] , \CARRYB[5][45] ,
         \CARRYB[5][44] , \CARRYB[5][43] , \CARRYB[5][42] , \CARRYB[5][41] ,
         \CARRYB[5][40] , \CARRYB[5][39] , \CARRYB[5][38] , \CARRYB[5][37] ,
         \CARRYB[5][36] , \CARRYB[5][35] , \CARRYB[5][34] , \CARRYB[5][33] ,
         \CARRYB[5][32] , \CARRYB[5][31] , \CARRYB[5][30] , \CARRYB[5][29] ,
         \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] ,
         \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] ,
         \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] ,
         \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][94] , \CARRYB[4][93] , \CARRYB[4][92] ,
         \CARRYB[4][91] , \CARRYB[4][90] , \CARRYB[4][89] , \CARRYB[4][88] ,
         \CARRYB[4][87] , \CARRYB[4][86] , \CARRYB[4][85] , \CARRYB[4][84] ,
         \CARRYB[4][83] , \CARRYB[4][82] , \CARRYB[4][81] , \CARRYB[4][80] ,
         \CARRYB[4][79] , \CARRYB[4][78] , \CARRYB[4][77] , \CARRYB[4][76] ,
         \CARRYB[4][75] , \CARRYB[4][74] , \CARRYB[4][73] , \CARRYB[4][72] ,
         \CARRYB[4][71] , \CARRYB[4][70] , \CARRYB[4][69] , \CARRYB[4][68] ,
         \CARRYB[4][67] , \CARRYB[4][66] , \CARRYB[4][65] , \CARRYB[4][64] ,
         \CARRYB[4][63] , \CARRYB[4][62] , \CARRYB[4][61] , \CARRYB[4][60] ,
         \CARRYB[4][59] , \CARRYB[4][58] , \CARRYB[4][57] , \CARRYB[4][56] ,
         \CARRYB[4][55] , \CARRYB[4][54] , \CARRYB[4][53] , \CARRYB[4][52] ,
         \CARRYB[4][51] , \CARRYB[4][50] , \CARRYB[4][49] , \CARRYB[4][48] ,
         \CARRYB[4][47] , \CARRYB[4][46] , \CARRYB[4][45] , \CARRYB[4][44] ,
         \CARRYB[4][43] , \CARRYB[4][42] , \CARRYB[4][41] , \CARRYB[4][40] ,
         \CARRYB[4][39] , \CARRYB[4][38] , \CARRYB[4][37] , \CARRYB[4][36] ,
         \CARRYB[4][35] , \CARRYB[4][34] , \CARRYB[4][33] , \CARRYB[4][32] ,
         \CARRYB[4][31] , \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] ,
         \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] ,
         \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] ,
         \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] ,
         \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][94] , \CARRYB[3][93] , \CARRYB[3][92] , \CARRYB[3][91] ,
         \CARRYB[3][90] , \CARRYB[3][89] , \CARRYB[3][88] , \CARRYB[3][87] ,
         \CARRYB[3][86] , \CARRYB[3][85] , \CARRYB[3][84] , \CARRYB[3][83] ,
         \CARRYB[3][82] , \CARRYB[3][81] , \CARRYB[3][80] , \CARRYB[3][79] ,
         \CARRYB[3][78] , \CARRYB[3][77] , \CARRYB[3][76] , \CARRYB[3][75] ,
         \CARRYB[3][74] , \CARRYB[3][73] , \CARRYB[3][72] , \CARRYB[3][71] ,
         \CARRYB[3][70] , \CARRYB[3][69] , \CARRYB[3][68] , \CARRYB[3][67] ,
         \CARRYB[3][66] , \CARRYB[3][65] , \CARRYB[3][64] , \CARRYB[3][63] ,
         \CARRYB[3][62] , \CARRYB[3][61] , \CARRYB[3][60] , \CARRYB[3][59] ,
         \CARRYB[3][58] , \CARRYB[3][57] , \CARRYB[3][56] , \CARRYB[3][55] ,
         \CARRYB[3][54] , \CARRYB[3][53] , \CARRYB[3][52] , \CARRYB[3][51] ,
         \CARRYB[3][50] , \CARRYB[3][49] , \CARRYB[3][48] , \CARRYB[3][47] ,
         \CARRYB[3][46] , \CARRYB[3][45] , \CARRYB[3][44] , \CARRYB[3][43] ,
         \CARRYB[3][42] , \CARRYB[3][41] , \CARRYB[3][40] , \CARRYB[3][39] ,
         \CARRYB[3][38] , \CARRYB[3][37] , \CARRYB[3][36] , \CARRYB[3][35] ,
         \CARRYB[3][34] , \CARRYB[3][33] , \CARRYB[3][32] , \SUMB[8][63] ,
         \SUMB[8][62] , \SUMB[8][61] , \SUMB[8][60] , \SUMB[8][59] ,
         \SUMB[8][58] , \SUMB[8][57] , \SUMB[8][56] , \SUMB[8][55] ,
         \SUMB[8][54] , \SUMB[8][53] , \SUMB[8][52] , \SUMB[8][51] ,
         \SUMB[8][50] , \SUMB[8][49] , \SUMB[8][48] , \SUMB[8][47] ,
         \SUMB[8][46] , \SUMB[8][45] , \SUMB[8][44] , \SUMB[8][43] ,
         \SUMB[8][42] , \SUMB[8][41] , \SUMB[8][40] , \SUMB[8][39] ,
         \SUMB[8][38] , \SUMB[8][37] , \SUMB[8][36] , \SUMB[8][35] ,
         \SUMB[8][34] , \SUMB[8][33] , \SUMB[8][32] , \SUMB[8][31] ,
         \SUMB[8][30] , \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] ,
         \SUMB[8][26] , \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] ,
         \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][94] , \SUMB[7][93] , \SUMB[7][92] , \SUMB[7][91] ,
         \SUMB[7][90] , \SUMB[7][89] , \SUMB[7][88] , \SUMB[7][87] ,
         \SUMB[7][86] , \SUMB[7][85] , \SUMB[7][84] , \SUMB[7][83] ,
         \SUMB[7][82] , \SUMB[7][81] , \SUMB[7][80] , \SUMB[7][79] ,
         \SUMB[7][78] , \SUMB[7][77] , \SUMB[7][76] , \SUMB[7][75] ,
         \SUMB[7][74] , \SUMB[7][73] , \SUMB[7][72] , \SUMB[7][71] ,
         \SUMB[7][70] , \SUMB[7][69] , \SUMB[7][68] , \SUMB[7][67] ,
         \SUMB[7][66] , \SUMB[7][65] , \SUMB[7][64] , \SUMB[7][63] ,
         \SUMB[7][62] , \SUMB[7][61] , \SUMB[7][60] , \SUMB[7][59] ,
         \SUMB[7][58] , \SUMB[7][57] , \SUMB[7][56] , \SUMB[7][55] ,
         \SUMB[7][54] , \SUMB[7][53] , \SUMB[7][52] , \SUMB[7][51] ,
         \SUMB[7][50] , \SUMB[7][49] , \SUMB[7][48] , \SUMB[7][47] ,
         \SUMB[7][46] , \SUMB[7][45] , \SUMB[7][44] , \SUMB[7][43] ,
         \SUMB[7][42] , \SUMB[7][41] , \SUMB[7][40] , \SUMB[7][39] ,
         \SUMB[7][38] , \SUMB[7][37] , \SUMB[7][36] , \SUMB[7][35] ,
         \SUMB[7][34] , \SUMB[7][33] , \SUMB[7][32] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][94] , \SUMB[6][93] , \SUMB[6][92] , \SUMB[6][91] ,
         \SUMB[6][90] , \SUMB[6][89] , \SUMB[6][88] , \SUMB[6][87] ,
         \SUMB[6][86] , \SUMB[6][85] , \SUMB[6][84] , \SUMB[6][83] ,
         \SUMB[6][82] , \SUMB[6][81] , \SUMB[6][80] , \SUMB[6][79] ,
         \SUMB[6][78] , \SUMB[6][77] , \SUMB[6][76] , \SUMB[6][75] ,
         \SUMB[6][74] , \SUMB[6][73] , \SUMB[6][72] , \SUMB[6][71] ,
         \SUMB[6][70] , \SUMB[6][69] , \SUMB[6][68] , \SUMB[6][67] ,
         \SUMB[6][66] , \SUMB[6][65] , \SUMB[6][64] , \SUMB[6][63] ,
         \SUMB[6][62] , \SUMB[6][61] , \SUMB[6][60] , \SUMB[6][59] ,
         \SUMB[6][58] , \SUMB[6][57] , \SUMB[6][56] , \SUMB[6][55] ,
         \SUMB[6][54] , \SUMB[6][53] , \SUMB[6][52] , \SUMB[6][51] ,
         \SUMB[6][50] , \SUMB[6][49] , \SUMB[6][48] , \SUMB[6][47] ,
         \SUMB[6][46] , \SUMB[6][45] , \SUMB[6][44] , \SUMB[6][43] ,
         \SUMB[6][42] , \SUMB[6][41] , \SUMB[6][40] , \SUMB[6][39] ,
         \SUMB[6][38] , \SUMB[6][37] , \SUMB[6][36] , \SUMB[6][35] ,
         \SUMB[6][34] , \SUMB[6][33] , \SUMB[6][32] , \SUMB[6][31] ,
         \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] ,
         \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] ,
         \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] ,
         \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][94] , \SUMB[5][93] , \SUMB[5][92] , \SUMB[5][91] ,
         \SUMB[5][90] , \SUMB[5][89] , \SUMB[5][88] , \SUMB[5][87] ,
         \SUMB[5][86] , \SUMB[5][85] , \SUMB[5][84] , \SUMB[5][83] ,
         \SUMB[5][82] , \SUMB[5][81] , \SUMB[5][80] , \SUMB[5][79] ,
         \SUMB[5][78] , \SUMB[5][77] , \SUMB[5][76] , \SUMB[5][75] ,
         \SUMB[5][74] , \SUMB[5][73] , \SUMB[5][72] , \SUMB[5][71] ,
         \SUMB[5][70] , \SUMB[5][69] , \SUMB[5][68] , \SUMB[5][67] ,
         \SUMB[5][66] , \SUMB[5][65] , \SUMB[5][64] , \SUMB[5][63] ,
         \SUMB[5][62] , \SUMB[5][61] , \SUMB[5][60] , \SUMB[5][59] ,
         \SUMB[5][58] , \SUMB[5][57] , \SUMB[5][56] , \SUMB[5][55] ,
         \SUMB[5][54] , \SUMB[5][53] , \SUMB[5][52] , \SUMB[5][51] ,
         \SUMB[5][50] , \SUMB[5][49] , \SUMB[5][48] , \SUMB[5][47] ,
         \SUMB[5][46] , \SUMB[5][45] , \SUMB[5][44] , \SUMB[5][43] ,
         \SUMB[5][42] , \SUMB[5][41] , \SUMB[5][40] , \SUMB[5][39] ,
         \SUMB[5][38] , \SUMB[5][37] , \SUMB[5][36] , \SUMB[5][35] ,
         \SUMB[5][34] , \SUMB[5][33] , \SUMB[5][32] , \SUMB[5][31] ,
         \SUMB[5][30] , \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] ,
         \SUMB[5][26] , \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] ,
         \SUMB[5][22] , \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] ,
         \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][94] , \SUMB[4][93] , \SUMB[4][92] , \SUMB[4][91] ,
         \SUMB[4][90] , \SUMB[4][89] , \SUMB[4][88] , \SUMB[4][87] ,
         \SUMB[4][86] , \SUMB[4][85] , \SUMB[4][84] , \SUMB[4][83] ,
         \SUMB[4][82] , \SUMB[4][81] , \SUMB[4][80] , \SUMB[4][79] ,
         \SUMB[4][78] , \SUMB[4][77] , \SUMB[4][76] , \SUMB[4][75] ,
         \SUMB[4][74] , \SUMB[4][73] , \SUMB[4][72] , \SUMB[4][71] ,
         \SUMB[4][70] , \SUMB[4][69] , \SUMB[4][68] , \SUMB[4][67] ,
         \SUMB[4][66] , \SUMB[4][65] , \SUMB[4][64] , \SUMB[4][63] ,
         \SUMB[4][62] , \SUMB[4][61] , \SUMB[4][60] , \SUMB[4][59] ,
         \SUMB[4][58] , \SUMB[4][57] , \SUMB[4][56] , \SUMB[4][55] ,
         \SUMB[4][54] , \SUMB[4][53] , \SUMB[4][52] , \SUMB[4][51] ,
         \SUMB[4][50] , \SUMB[4][49] , \SUMB[4][48] , \SUMB[4][47] ,
         \SUMB[4][46] , \SUMB[4][45] , \SUMB[4][44] , \SUMB[4][43] ,
         \SUMB[4][42] , \SUMB[4][41] , \SUMB[4][40] , \SUMB[4][39] ,
         \SUMB[4][38] , \SUMB[4][37] , \SUMB[4][36] , \SUMB[4][35] ,
         \SUMB[4][34] , \SUMB[4][33] , \SUMB[4][32] , \SUMB[4][31] ,
         \SUMB[4][30] , \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] ,
         \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][94] , \SUMB[3][93] , \SUMB[3][92] , \SUMB[3][91] ,
         \SUMB[3][90] , \SUMB[3][89] , \SUMB[3][88] , \SUMB[3][87] ,
         \SUMB[3][86] , \SUMB[3][85] , \SUMB[3][84] , \SUMB[3][83] ,
         \SUMB[3][82] , \SUMB[3][81] , \SUMB[3][80] , \SUMB[3][79] ,
         \SUMB[3][78] , \SUMB[3][77] , \SUMB[3][76] , \SUMB[3][75] ,
         \SUMB[3][74] , \SUMB[3][73] , \SUMB[3][72] , \SUMB[3][71] ,
         \SUMB[3][70] , \SUMB[3][69] , \SUMB[3][68] , \SUMB[3][67] ,
         \SUMB[3][66] , \SUMB[3][65] , \SUMB[3][64] , \SUMB[3][63] ,
         \SUMB[3][62] , \SUMB[3][61] , \SUMB[3][60] , \SUMB[3][59] ,
         \SUMB[3][58] , \SUMB[3][57] , \SUMB[3][56] , \SUMB[3][55] ,
         \SUMB[3][54] , \SUMB[3][53] , \SUMB[3][52] , \SUMB[3][51] ,
         \SUMB[3][50] , \SUMB[3][49] , \SUMB[3][48] , \SUMB[3][47] ,
         \SUMB[3][46] , \SUMB[3][45] , \SUMB[3][44] , \SUMB[3][43] ,
         \SUMB[3][42] , \SUMB[3][41] , \SUMB[3][40] , \SUMB[3][39] ,
         \SUMB[3][38] , \SUMB[3][37] , \SUMB[3][36] , \SUMB[3][35] ,
         \SUMB[3][34] , \SUMB[3][33] , \SUMB[3][32] , \CARRYB[13][94] ,
         \CARRYB[13][93] , \CARRYB[13][92] , \CARRYB[13][91] ,
         \CARRYB[13][90] , \CARRYB[13][89] , \CARRYB[13][88] ,
         \CARRYB[13][87] , \CARRYB[13][86] , \CARRYB[13][85] ,
         \CARRYB[13][84] , \CARRYB[13][83] , \CARRYB[13][82] ,
         \CARRYB[13][81] , \CARRYB[13][80] , \CARRYB[13][79] ,
         \CARRYB[13][78] , \CARRYB[13][77] , \CARRYB[13][76] ,
         \CARRYB[13][75] , \CARRYB[13][74] , \CARRYB[13][73] ,
         \CARRYB[13][72] , \CARRYB[13][71] , \CARRYB[13][70] ,
         \CARRYB[13][69] , \CARRYB[13][68] , \CARRYB[13][67] ,
         \CARRYB[13][66] , \CARRYB[13][65] , \CARRYB[13][64] ,
         \CARRYB[13][63] , \CARRYB[13][62] , \CARRYB[13][61] ,
         \CARRYB[13][60] , \CARRYB[13][59] , \CARRYB[13][58] ,
         \CARRYB[13][57] , \CARRYB[13][56] , \CARRYB[13][55] ,
         \CARRYB[13][54] , \CARRYB[13][53] , \CARRYB[13][52] ,
         \CARRYB[13][51] , \CARRYB[13][50] , \CARRYB[13][49] ,
         \CARRYB[13][48] , \CARRYB[13][47] , \CARRYB[13][46] ,
         \CARRYB[13][45] , \CARRYB[13][44] , \CARRYB[13][43] ,
         \CARRYB[13][42] , \CARRYB[13][41] , \CARRYB[13][40] ,
         \CARRYB[13][39] , \CARRYB[13][38] , \CARRYB[13][37] ,
         \CARRYB[13][36] , \CARRYB[13][35] , \CARRYB[13][34] ,
         \CARRYB[13][33] , \CARRYB[13][32] , \CARRYB[13][31] ,
         \CARRYB[13][30] , \CARRYB[13][29] , \CARRYB[13][28] ,
         \CARRYB[13][27] , \CARRYB[13][26] , \CARRYB[13][25] ,
         \CARRYB[13][24] , \CARRYB[13][23] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][94] , \CARRYB[12][93] , \CARRYB[12][92] ,
         \CARRYB[12][91] , \CARRYB[12][90] , \CARRYB[12][89] ,
         \CARRYB[12][88] , \CARRYB[12][87] , \CARRYB[12][86] ,
         \CARRYB[12][85] , \CARRYB[12][84] , \CARRYB[12][83] ,
         \CARRYB[12][82] , \CARRYB[12][81] , \CARRYB[12][80] ,
         \CARRYB[12][79] , \CARRYB[12][78] , \CARRYB[12][77] ,
         \CARRYB[12][76] , \CARRYB[12][75] , \CARRYB[12][74] ,
         \CARRYB[12][73] , \CARRYB[12][72] , \CARRYB[12][71] ,
         \CARRYB[12][70] , \CARRYB[12][69] , \CARRYB[12][68] ,
         \CARRYB[12][67] , \CARRYB[12][66] , \CARRYB[12][65] ,
         \CARRYB[12][64] , \CARRYB[12][63] , \CARRYB[12][62] ,
         \CARRYB[12][61] , \CARRYB[12][60] , \CARRYB[12][59] ,
         \CARRYB[12][58] , \CARRYB[12][57] , \CARRYB[12][56] ,
         \CARRYB[12][55] , \CARRYB[12][54] , \CARRYB[12][53] ,
         \CARRYB[12][52] , \CARRYB[12][51] , \CARRYB[12][50] ,
         \CARRYB[12][49] , \CARRYB[12][48] , \CARRYB[12][47] ,
         \CARRYB[12][46] , \CARRYB[12][45] , \CARRYB[12][44] ,
         \CARRYB[12][43] , \CARRYB[12][42] , \CARRYB[12][41] ,
         \CARRYB[12][40] , \CARRYB[12][39] , \CARRYB[12][38] ,
         \CARRYB[12][37] , \CARRYB[12][36] , \CARRYB[12][35] ,
         \CARRYB[12][34] , \CARRYB[12][33] , \CARRYB[12][32] ,
         \CARRYB[12][31] , \CARRYB[12][30] , \CARRYB[12][29] ,
         \CARRYB[12][28] , \CARRYB[12][27] , \CARRYB[12][26] ,
         \CARRYB[12][25] , \CARRYB[12][24] , \CARRYB[12][23] ,
         \CARRYB[12][22] , \CARRYB[12][21] , \CARRYB[12][20] ,
         \CARRYB[12][19] , \CARRYB[12][18] , \CARRYB[12][17] ,
         \CARRYB[12][16] , \CARRYB[12][15] , \CARRYB[12][14] ,
         \CARRYB[12][13] , \CARRYB[12][12] , \CARRYB[12][11] ,
         \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] , \CARRYB[12][7] ,
         \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] , \CARRYB[11][94] ,
         \CARRYB[11][93] , \CARRYB[11][92] , \CARRYB[11][91] ,
         \CARRYB[11][90] , \CARRYB[11][89] , \CARRYB[11][88] ,
         \CARRYB[11][87] , \CARRYB[11][86] , \CARRYB[11][85] ,
         \CARRYB[11][84] , \CARRYB[11][83] , \CARRYB[11][82] ,
         \CARRYB[11][81] , \CARRYB[11][80] , \CARRYB[11][79] ,
         \CARRYB[11][78] , \CARRYB[11][77] , \CARRYB[11][76] ,
         \CARRYB[11][75] , \CARRYB[11][74] , \CARRYB[11][73] ,
         \CARRYB[11][72] , \CARRYB[11][71] , \CARRYB[11][70] ,
         \CARRYB[11][69] , \CARRYB[11][68] , \CARRYB[11][67] ,
         \CARRYB[11][66] , \CARRYB[11][65] , \CARRYB[11][64] ,
         \CARRYB[11][63] , \CARRYB[11][62] , \CARRYB[11][61] ,
         \CARRYB[11][60] , \CARRYB[11][59] , \CARRYB[11][58] ,
         \CARRYB[11][57] , \CARRYB[11][56] , \CARRYB[11][55] ,
         \CARRYB[11][54] , \CARRYB[11][53] , \CARRYB[11][52] ,
         \CARRYB[11][51] , \CARRYB[11][50] , \CARRYB[11][49] ,
         \CARRYB[11][48] , \CARRYB[11][47] , \CARRYB[11][46] ,
         \CARRYB[11][45] , \CARRYB[11][44] , \CARRYB[11][43] ,
         \CARRYB[11][42] , \CARRYB[11][41] , \CARRYB[11][40] ,
         \CARRYB[11][39] , \CARRYB[11][38] , \CARRYB[11][37] ,
         \CARRYB[11][36] , \CARRYB[11][35] , \CARRYB[11][34] ,
         \CARRYB[11][33] , \CARRYB[11][32] , \CARRYB[11][31] ,
         \CARRYB[11][30] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][23] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][94] , \CARRYB[10][93] , \CARRYB[10][92] ,
         \CARRYB[10][91] , \CARRYB[10][90] , \CARRYB[10][89] ,
         \CARRYB[10][88] , \CARRYB[10][87] , \CARRYB[10][86] ,
         \CARRYB[10][85] , \CARRYB[10][84] , \CARRYB[10][83] ,
         \CARRYB[10][82] , \CARRYB[10][81] , \CARRYB[10][80] ,
         \CARRYB[10][79] , \CARRYB[10][78] , \CARRYB[10][77] ,
         \CARRYB[10][76] , \CARRYB[10][75] , \CARRYB[10][74] ,
         \CARRYB[10][73] , \CARRYB[10][72] , \CARRYB[10][71] ,
         \CARRYB[10][70] , \CARRYB[10][69] , \CARRYB[10][68] ,
         \CARRYB[10][67] , \CARRYB[10][66] , \CARRYB[10][65] ,
         \CARRYB[10][64] , \CARRYB[10][63] , \CARRYB[10][62] ,
         \CARRYB[10][61] , \CARRYB[10][60] , \CARRYB[10][59] ,
         \CARRYB[10][58] , \CARRYB[10][57] , \CARRYB[10][56] ,
         \CARRYB[10][55] , \CARRYB[10][54] , \CARRYB[10][53] ,
         \CARRYB[10][52] , \CARRYB[10][51] , \CARRYB[10][50] ,
         \CARRYB[10][49] , \CARRYB[10][48] , \CARRYB[10][47] ,
         \CARRYB[10][46] , \CARRYB[10][45] , \CARRYB[10][44] ,
         \CARRYB[10][43] , \CARRYB[10][42] , \CARRYB[10][41] ,
         \CARRYB[10][40] , \CARRYB[10][39] , \CARRYB[10][38] ,
         \CARRYB[10][37] , \CARRYB[10][36] , \CARRYB[10][35] ,
         \CARRYB[10][34] , \CARRYB[10][33] , \CARRYB[10][32] ,
         \CARRYB[10][31] , \CARRYB[10][30] , \CARRYB[10][29] ,
         \CARRYB[10][28] , \CARRYB[10][27] , \CARRYB[10][26] ,
         \CARRYB[10][25] , \CARRYB[10][24] , \CARRYB[10][23] ,
         \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][94] ,
         \CARRYB[9][93] , \CARRYB[9][92] , \CARRYB[9][91] , \CARRYB[9][90] ,
         \CARRYB[9][89] , \CARRYB[9][88] , \CARRYB[9][87] , \CARRYB[9][86] ,
         \CARRYB[9][85] , \CARRYB[9][84] , \CARRYB[9][83] , \CARRYB[9][82] ,
         \CARRYB[9][81] , \CARRYB[9][80] , \CARRYB[9][79] , \CARRYB[9][78] ,
         \CARRYB[9][77] , \CARRYB[9][76] , \CARRYB[9][75] , \CARRYB[9][74] ,
         \CARRYB[9][73] , \CARRYB[9][72] , \CARRYB[9][71] , \CARRYB[9][70] ,
         \CARRYB[9][69] , \CARRYB[9][68] , \CARRYB[9][67] , \CARRYB[9][66] ,
         \CARRYB[9][65] , \CARRYB[9][64] , \CARRYB[9][63] , \CARRYB[9][62] ,
         \CARRYB[9][61] , \CARRYB[9][60] , \CARRYB[9][59] , \CARRYB[9][58] ,
         \CARRYB[9][57] , \CARRYB[9][56] , \CARRYB[9][55] , \CARRYB[9][54] ,
         \CARRYB[9][53] , \CARRYB[9][52] , \CARRYB[9][51] , \CARRYB[9][50] ,
         \CARRYB[9][49] , \CARRYB[9][48] , \CARRYB[9][47] , \CARRYB[9][46] ,
         \CARRYB[9][45] , \CARRYB[9][44] , \CARRYB[9][43] , \CARRYB[9][42] ,
         \CARRYB[9][41] , \CARRYB[9][40] , \CARRYB[9][39] , \CARRYB[9][38] ,
         \CARRYB[9][37] , \CARRYB[9][36] , \CARRYB[9][35] , \CARRYB[9][34] ,
         \CARRYB[9][33] , \CARRYB[9][32] , \CARRYB[9][31] , \CARRYB[9][30] ,
         \CARRYB[9][29] , \CARRYB[9][28] , \CARRYB[9][27] , \CARRYB[9][26] ,
         \CARRYB[9][25] , \CARRYB[9][24] , \CARRYB[9][23] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][94] , \CARRYB[8][93] ,
         \CARRYB[8][92] , \CARRYB[8][91] , \CARRYB[8][90] , \CARRYB[8][89] ,
         \CARRYB[8][88] , \CARRYB[8][87] , \CARRYB[8][86] , \CARRYB[8][85] ,
         \CARRYB[8][84] , \CARRYB[8][83] , \CARRYB[8][82] , \CARRYB[8][81] ,
         \CARRYB[8][80] , \CARRYB[8][79] , \CARRYB[8][78] , \CARRYB[8][77] ,
         \CARRYB[8][76] , \CARRYB[8][75] , \CARRYB[8][74] , \CARRYB[8][73] ,
         \CARRYB[8][72] , \CARRYB[8][71] , \CARRYB[8][70] , \CARRYB[8][69] ,
         \CARRYB[8][68] , \CARRYB[8][67] , \CARRYB[8][66] , \CARRYB[8][65] ,
         \CARRYB[8][64] , \SUMB[13][94] , \SUMB[13][93] , \SUMB[13][92] ,
         \SUMB[13][91] , \SUMB[13][90] , \SUMB[13][89] , \SUMB[13][88] ,
         \SUMB[13][87] , \SUMB[13][86] , \SUMB[13][85] , \SUMB[13][84] ,
         \SUMB[13][83] , \SUMB[13][82] , \SUMB[13][81] , \SUMB[13][80] ,
         \SUMB[13][79] , \SUMB[13][78] , \SUMB[13][77] , \SUMB[13][76] ,
         \SUMB[13][75] , \SUMB[13][74] , \SUMB[13][73] , \SUMB[13][72] ,
         \SUMB[13][71] , \SUMB[13][70] , \SUMB[13][69] , \SUMB[13][68] ,
         \SUMB[13][67] , \SUMB[13][66] , \SUMB[13][65] , \SUMB[13][64] ,
         \SUMB[13][63] , \SUMB[13][62] , \SUMB[13][61] , \SUMB[13][60] ,
         \SUMB[13][59] , \SUMB[13][58] , \SUMB[13][57] , \SUMB[13][56] ,
         \SUMB[13][55] , \SUMB[13][54] , \SUMB[13][53] , \SUMB[13][52] ,
         \SUMB[13][51] , \SUMB[13][50] , \SUMB[13][49] , \SUMB[13][48] ,
         \SUMB[13][47] , \SUMB[13][46] , \SUMB[13][45] , \SUMB[13][44] ,
         \SUMB[13][43] , \SUMB[13][42] , \SUMB[13][41] , \SUMB[13][40] ,
         \SUMB[13][39] , \SUMB[13][38] , \SUMB[13][37] , \SUMB[13][36] ,
         \SUMB[13][35] , \SUMB[13][34] , \SUMB[13][33] , \SUMB[13][32] ,
         \SUMB[13][31] , \SUMB[13][30] , \SUMB[13][29] , \SUMB[13][28] ,
         \SUMB[13][27] , \SUMB[13][26] , \SUMB[13][25] , \SUMB[13][24] ,
         \SUMB[13][23] , \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] ,
         \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] ,
         \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][94] ,
         \SUMB[12][93] , \SUMB[12][92] , \SUMB[12][91] , \SUMB[12][90] ,
         \SUMB[12][89] , \SUMB[12][88] , \SUMB[12][87] , \SUMB[12][86] ,
         \SUMB[12][85] , \SUMB[12][84] , \SUMB[12][83] , \SUMB[12][82] ,
         \SUMB[12][81] , \SUMB[12][80] , \SUMB[12][79] , \SUMB[12][78] ,
         \SUMB[12][77] , \SUMB[12][76] , \SUMB[12][75] , \SUMB[12][74] ,
         \SUMB[12][73] , \SUMB[12][72] , \SUMB[12][71] , \SUMB[12][70] ,
         \SUMB[12][69] , \SUMB[12][68] , \SUMB[12][67] , \SUMB[12][66] ,
         \SUMB[12][65] , \SUMB[12][64] , \SUMB[12][63] , \SUMB[12][62] ,
         \SUMB[12][61] , \SUMB[12][60] , \SUMB[12][59] , \SUMB[12][58] ,
         \SUMB[12][57] , \SUMB[12][56] , \SUMB[12][55] , \SUMB[12][54] ,
         \SUMB[12][53] , \SUMB[12][52] , \SUMB[12][51] , \SUMB[12][50] ,
         \SUMB[12][49] , \SUMB[12][48] , \SUMB[12][47] , \SUMB[12][46] ,
         \SUMB[12][45] , \SUMB[12][44] , \SUMB[12][43] , \SUMB[12][42] ,
         \SUMB[12][41] , \SUMB[12][40] , \SUMB[12][39] , \SUMB[12][38] ,
         \SUMB[12][37] , \SUMB[12][36] , \SUMB[12][35] , \SUMB[12][34] ,
         \SUMB[12][33] , \SUMB[12][32] , \SUMB[12][31] , \SUMB[12][30] ,
         \SUMB[12][29] , \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] ,
         \SUMB[12][25] , \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] ,
         \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] ,
         \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][94] , \SUMB[11][93] , \SUMB[11][92] ,
         \SUMB[11][91] , \SUMB[11][90] , \SUMB[11][89] , \SUMB[11][88] ,
         \SUMB[11][87] , \SUMB[11][86] , \SUMB[11][85] , \SUMB[11][84] ,
         \SUMB[11][83] , \SUMB[11][82] , \SUMB[11][81] , \SUMB[11][80] ,
         \SUMB[11][79] , \SUMB[11][78] , \SUMB[11][77] , \SUMB[11][76] ,
         \SUMB[11][75] , \SUMB[11][74] , \SUMB[11][73] , \SUMB[11][72] ,
         \SUMB[11][71] , \SUMB[11][70] , \SUMB[11][69] , \SUMB[11][68] ,
         \SUMB[11][67] , \SUMB[11][66] , \SUMB[11][65] , \SUMB[11][64] ,
         \SUMB[11][63] , \SUMB[11][62] , \SUMB[11][61] , \SUMB[11][60] ,
         \SUMB[11][59] , \SUMB[11][58] , \SUMB[11][57] , \SUMB[11][56] ,
         \SUMB[11][55] , \SUMB[11][54] , \SUMB[11][53] , \SUMB[11][52] ,
         \SUMB[11][51] , \SUMB[11][50] , \SUMB[11][49] , \SUMB[11][48] ,
         \SUMB[11][47] , \SUMB[11][46] , \SUMB[11][45] , \SUMB[11][44] ,
         \SUMB[11][43] , \SUMB[11][42] , \SUMB[11][41] , \SUMB[11][40] ,
         \SUMB[11][39] , \SUMB[11][38] , \SUMB[11][37] , \SUMB[11][36] ,
         \SUMB[11][35] , \SUMB[11][34] , \SUMB[11][33] , \SUMB[11][32] ,
         \SUMB[11][31] , \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] ,
         \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] ,
         \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][94] ,
         \SUMB[10][93] , \SUMB[10][92] , \SUMB[10][91] , \SUMB[10][90] ,
         \SUMB[10][89] , \SUMB[10][88] , \SUMB[10][87] , \SUMB[10][86] ,
         \SUMB[10][85] , \SUMB[10][84] , \SUMB[10][83] , \SUMB[10][82] ,
         \SUMB[10][81] , \SUMB[10][80] , \SUMB[10][79] , \SUMB[10][78] ,
         \SUMB[10][77] , \SUMB[10][76] , \SUMB[10][75] , \SUMB[10][74] ,
         \SUMB[10][73] , \SUMB[10][72] , \SUMB[10][71] , \SUMB[10][70] ,
         \SUMB[10][69] , \SUMB[10][68] , \SUMB[10][67] , \SUMB[10][66] ,
         \SUMB[10][65] , \SUMB[10][64] , \SUMB[10][63] , \SUMB[10][62] ,
         \SUMB[10][61] , \SUMB[10][60] , \SUMB[10][59] , \SUMB[10][58] ,
         \SUMB[10][57] , \SUMB[10][56] , \SUMB[10][55] , \SUMB[10][54] ,
         \SUMB[10][53] , \SUMB[10][52] , \SUMB[10][51] , \SUMB[10][50] ,
         \SUMB[10][49] , \SUMB[10][48] , \SUMB[10][47] , \SUMB[10][46] ,
         \SUMB[10][45] , \SUMB[10][44] , \SUMB[10][43] , \SUMB[10][42] ,
         \SUMB[10][41] , \SUMB[10][40] , \SUMB[10][39] , \SUMB[10][38] ,
         \SUMB[10][37] , \SUMB[10][36] , \SUMB[10][35] , \SUMB[10][34] ,
         \SUMB[10][33] , \SUMB[10][32] , \SUMB[10][31] , \SUMB[10][30] ,
         \SUMB[10][29] , \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] ,
         \SUMB[10][25] , \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] ,
         \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] ,
         \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][94] , \SUMB[9][93] , \SUMB[9][92] ,
         \SUMB[9][91] , \SUMB[9][90] , \SUMB[9][89] , \SUMB[9][88] ,
         \SUMB[9][87] , \SUMB[9][86] , \SUMB[9][85] , \SUMB[9][84] ,
         \SUMB[9][83] , \SUMB[9][82] , \SUMB[9][81] , \SUMB[9][80] ,
         \SUMB[9][79] , \SUMB[9][78] , \SUMB[9][77] , \SUMB[9][76] ,
         \SUMB[9][75] , \SUMB[9][74] , \SUMB[9][73] , \SUMB[9][72] ,
         \SUMB[9][71] , \SUMB[9][70] , \SUMB[9][69] , \SUMB[9][68] ,
         \SUMB[9][67] , \SUMB[9][66] , \SUMB[9][65] , \SUMB[9][64] ,
         \SUMB[9][63] , \SUMB[9][62] , \SUMB[9][61] , \SUMB[9][60] ,
         \SUMB[9][59] , \SUMB[9][58] , \SUMB[9][57] , \SUMB[9][56] ,
         \SUMB[9][55] , \SUMB[9][54] , \SUMB[9][53] , \SUMB[9][52] ,
         \SUMB[9][51] , \SUMB[9][50] , \SUMB[9][49] , \SUMB[9][48] ,
         \SUMB[9][47] , \SUMB[9][46] , \SUMB[9][45] , \SUMB[9][44] ,
         \SUMB[9][43] , \SUMB[9][42] , \SUMB[9][41] , \SUMB[9][40] ,
         \SUMB[9][39] , \SUMB[9][38] , \SUMB[9][37] , \SUMB[9][36] ,
         \SUMB[9][35] , \SUMB[9][34] , \SUMB[9][33] , \SUMB[9][32] ,
         \SUMB[9][31] , \SUMB[9][30] , \SUMB[9][29] , \SUMB[9][28] ,
         \SUMB[9][27] , \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] ,
         \SUMB[9][23] , \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] ,
         \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] ,
         \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][94] , \SUMB[8][93] ,
         \SUMB[8][92] , \SUMB[8][91] , \SUMB[8][90] , \SUMB[8][89] ,
         \SUMB[8][88] , \SUMB[8][87] , \SUMB[8][86] , \SUMB[8][85] ,
         \SUMB[8][84] , \SUMB[8][83] , \SUMB[8][82] , \SUMB[8][81] ,
         \SUMB[8][80] , \SUMB[8][79] , \SUMB[8][78] , \SUMB[8][77] ,
         \SUMB[8][76] , \SUMB[8][75] , \SUMB[8][74] , \SUMB[8][73] ,
         \SUMB[8][72] , \SUMB[8][71] , \SUMB[8][70] , \SUMB[8][69] ,
         \SUMB[8][68] , \SUMB[8][67] , \SUMB[8][66] , \SUMB[8][65] ,
         \SUMB[8][64] , \CARRYB[19][31] , \CARRYB[19][30] , \CARRYB[19][29] ,
         \CARRYB[19][28] , \CARRYB[19][27] , \CARRYB[19][26] ,
         \CARRYB[19][25] , \CARRYB[19][24] , \CARRYB[19][23] ,
         \CARRYB[19][22] , \CARRYB[19][21] , \CARRYB[19][20] ,
         \CARRYB[19][19] , \CARRYB[19][18] , \CARRYB[19][17] ,
         \CARRYB[19][16] , \CARRYB[19][15] , \CARRYB[19][14] ,
         \CARRYB[19][13] , \CARRYB[19][12] , \CARRYB[19][11] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][94] ,
         \CARRYB[18][93] , \CARRYB[18][92] , \CARRYB[18][91] ,
         \CARRYB[18][90] , \CARRYB[18][89] , \CARRYB[18][88] ,
         \CARRYB[18][87] , \CARRYB[18][86] , \CARRYB[18][85] ,
         \CARRYB[18][84] , \CARRYB[18][83] , \CARRYB[18][82] ,
         \CARRYB[18][81] , \CARRYB[18][80] , \CARRYB[18][79] ,
         \CARRYB[18][78] , \CARRYB[18][77] , \CARRYB[18][76] ,
         \CARRYB[18][75] , \CARRYB[18][74] , \CARRYB[18][73] ,
         \CARRYB[18][72] , \CARRYB[18][71] , \CARRYB[18][70] ,
         \CARRYB[18][69] , \CARRYB[18][68] , \CARRYB[18][67] ,
         \CARRYB[18][66] , \CARRYB[18][65] , \CARRYB[18][64] ,
         \CARRYB[18][63] , \CARRYB[18][62] , \CARRYB[18][61] ,
         \CARRYB[18][60] , \CARRYB[18][59] , \CARRYB[18][58] ,
         \CARRYB[18][57] , \CARRYB[18][56] , \CARRYB[18][55] ,
         \CARRYB[18][54] , \CARRYB[18][53] , \CARRYB[18][52] ,
         \CARRYB[18][51] , \CARRYB[18][50] , \CARRYB[18][49] ,
         \CARRYB[18][48] , \CARRYB[18][47] , \CARRYB[18][46] ,
         \CARRYB[18][45] , \CARRYB[18][44] , \CARRYB[18][43] ,
         \CARRYB[18][42] , \CARRYB[18][41] , \CARRYB[18][40] ,
         \CARRYB[18][39] , \CARRYB[18][38] , \CARRYB[18][37] ,
         \CARRYB[18][36] , \CARRYB[18][35] , \CARRYB[18][34] ,
         \CARRYB[18][33] , \CARRYB[18][32] , \CARRYB[18][31] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][94] , \CARRYB[17][93] , \CARRYB[17][92] ,
         \CARRYB[17][91] , \CARRYB[17][90] , \CARRYB[17][89] ,
         \CARRYB[17][88] , \CARRYB[17][87] , \CARRYB[17][86] ,
         \CARRYB[17][85] , \CARRYB[17][84] , \CARRYB[17][83] ,
         \CARRYB[17][82] , \CARRYB[17][81] , \CARRYB[17][80] ,
         \CARRYB[17][79] , \CARRYB[17][78] , \CARRYB[17][77] ,
         \CARRYB[17][76] , \CARRYB[17][75] , \CARRYB[17][74] ,
         \CARRYB[17][73] , \CARRYB[17][72] , \CARRYB[17][71] ,
         \CARRYB[17][70] , \CARRYB[17][69] , \CARRYB[17][68] ,
         \CARRYB[17][67] , \CARRYB[17][66] , \CARRYB[17][65] ,
         \CARRYB[17][64] , \CARRYB[17][63] , \CARRYB[17][62] ,
         \CARRYB[17][61] , \CARRYB[17][60] , \CARRYB[17][59] ,
         \CARRYB[17][58] , \CARRYB[17][57] , \CARRYB[17][56] ,
         \CARRYB[17][55] , \CARRYB[17][54] , \CARRYB[17][53] ,
         \CARRYB[17][52] , \CARRYB[17][51] , \CARRYB[17][50] ,
         \CARRYB[17][49] , \CARRYB[17][48] , \CARRYB[17][47] ,
         \CARRYB[17][46] , \CARRYB[17][45] , \CARRYB[17][44] ,
         \CARRYB[17][43] , \CARRYB[17][42] , \CARRYB[17][41] ,
         \CARRYB[17][40] , \CARRYB[17][39] , \CARRYB[17][38] ,
         \CARRYB[17][37] , \CARRYB[17][36] , \CARRYB[17][35] ,
         \CARRYB[17][34] , \CARRYB[17][33] , \CARRYB[17][32] ,
         \CARRYB[17][31] , \CARRYB[17][30] , \CARRYB[17][29] ,
         \CARRYB[17][28] , \CARRYB[17][27] , \CARRYB[17][26] ,
         \CARRYB[17][25] , \CARRYB[17][24] , \CARRYB[17][23] ,
         \CARRYB[17][22] , \CARRYB[17][21] , \CARRYB[17][20] ,
         \CARRYB[17][19] , \CARRYB[17][18] , \CARRYB[17][17] ,
         \CARRYB[17][16] , \CARRYB[17][15] , \CARRYB[17][14] ,
         \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][94] ,
         \CARRYB[16][93] , \CARRYB[16][92] , \CARRYB[16][91] ,
         \CARRYB[16][90] , \CARRYB[16][89] , \CARRYB[16][88] ,
         \CARRYB[16][87] , \CARRYB[16][86] , \CARRYB[16][85] ,
         \CARRYB[16][84] , \CARRYB[16][83] , \CARRYB[16][82] ,
         \CARRYB[16][81] , \CARRYB[16][80] , \CARRYB[16][79] ,
         \CARRYB[16][78] , \CARRYB[16][77] , \CARRYB[16][76] ,
         \CARRYB[16][75] , \CARRYB[16][74] , \CARRYB[16][73] ,
         \CARRYB[16][72] , \CARRYB[16][71] , \CARRYB[16][70] ,
         \CARRYB[16][69] , \CARRYB[16][68] , \CARRYB[16][67] ,
         \CARRYB[16][66] , \CARRYB[16][65] , \CARRYB[16][64] ,
         \CARRYB[16][63] , \CARRYB[16][62] , \CARRYB[16][61] ,
         \CARRYB[16][60] , \CARRYB[16][59] , \CARRYB[16][58] ,
         \CARRYB[16][57] , \CARRYB[16][56] , \CARRYB[16][55] ,
         \CARRYB[16][54] , \CARRYB[16][53] , \CARRYB[16][52] ,
         \CARRYB[16][51] , \CARRYB[16][50] , \CARRYB[16][49] ,
         \CARRYB[16][48] , \CARRYB[16][47] , \CARRYB[16][46] ,
         \CARRYB[16][45] , \CARRYB[16][44] , \CARRYB[16][43] ,
         \CARRYB[16][42] , \CARRYB[16][41] , \CARRYB[16][40] ,
         \CARRYB[16][39] , \CARRYB[16][38] , \CARRYB[16][37] ,
         \CARRYB[16][36] , \CARRYB[16][35] , \CARRYB[16][34] ,
         \CARRYB[16][33] , \CARRYB[16][32] , \CARRYB[16][31] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \CARRYB[15][94] , \CARRYB[15][93] , \CARRYB[15][92] ,
         \CARRYB[15][91] , \CARRYB[15][90] , \CARRYB[15][89] ,
         \CARRYB[15][88] , \CARRYB[15][87] , \CARRYB[15][86] ,
         \CARRYB[15][85] , \CARRYB[15][84] , \CARRYB[15][83] ,
         \CARRYB[15][82] , \CARRYB[15][81] , \CARRYB[15][80] ,
         \CARRYB[15][79] , \CARRYB[15][78] , \CARRYB[15][77] ,
         \CARRYB[15][76] , \CARRYB[15][75] , \CARRYB[15][74] ,
         \CARRYB[15][73] , \CARRYB[15][72] , \CARRYB[15][71] ,
         \CARRYB[15][70] , \CARRYB[15][69] , \CARRYB[15][68] ,
         \CARRYB[15][67] , \CARRYB[15][66] , \CARRYB[15][65] ,
         \CARRYB[15][64] , \CARRYB[15][63] , \CARRYB[15][62] ,
         \CARRYB[15][61] , \CARRYB[15][60] , \CARRYB[15][59] ,
         \CARRYB[15][58] , \CARRYB[15][57] , \CARRYB[15][56] ,
         \CARRYB[15][55] , \CARRYB[15][54] , \CARRYB[15][53] ,
         \CARRYB[15][52] , \CARRYB[15][51] , \CARRYB[15][50] ,
         \CARRYB[15][49] , \CARRYB[15][48] , \CARRYB[15][47] ,
         \CARRYB[15][46] , \CARRYB[15][45] , \CARRYB[15][44] ,
         \CARRYB[15][43] , \CARRYB[15][42] , \CARRYB[15][41] ,
         \CARRYB[15][40] , \CARRYB[15][39] , \CARRYB[15][38] ,
         \CARRYB[15][37] , \CARRYB[15][36] , \CARRYB[15][35] ,
         \CARRYB[15][34] , \CARRYB[15][33] , \CARRYB[15][32] ,
         \CARRYB[15][31] , \CARRYB[15][30] , \CARRYB[15][29] ,
         \CARRYB[15][28] , \CARRYB[15][27] , \CARRYB[15][26] ,
         \CARRYB[15][25] , \CARRYB[15][24] , \CARRYB[15][23] ,
         \CARRYB[15][22] , \CARRYB[15][21] , \CARRYB[15][20] ,
         \CARRYB[15][19] , \CARRYB[15][18] , \CARRYB[15][17] ,
         \CARRYB[15][16] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][94] ,
         \CARRYB[14][93] , \CARRYB[14][92] , \CARRYB[14][91] ,
         \CARRYB[14][90] , \CARRYB[14][89] , \CARRYB[14][88] ,
         \CARRYB[14][87] , \CARRYB[14][86] , \CARRYB[14][85] ,
         \CARRYB[14][84] , \CARRYB[14][83] , \CARRYB[14][82] ,
         \CARRYB[14][81] , \CARRYB[14][80] , \CARRYB[14][79] ,
         \CARRYB[14][78] , \CARRYB[14][77] , \CARRYB[14][76] ,
         \CARRYB[14][75] , \CARRYB[14][74] , \CARRYB[14][73] ,
         \CARRYB[14][72] , \CARRYB[14][71] , \CARRYB[14][70] ,
         \CARRYB[14][69] , \CARRYB[14][68] , \CARRYB[14][67] ,
         \CARRYB[14][66] , \CARRYB[14][65] , \CARRYB[14][64] ,
         \CARRYB[14][63] , \CARRYB[14][62] , \CARRYB[14][61] ,
         \CARRYB[14][60] , \CARRYB[14][59] , \CARRYB[14][58] ,
         \CARRYB[14][57] , \CARRYB[14][56] , \CARRYB[14][55] ,
         \CARRYB[14][54] , \CARRYB[14][53] , \CARRYB[14][52] ,
         \CARRYB[14][51] , \CARRYB[14][50] , \CARRYB[14][49] ,
         \CARRYB[14][48] , \CARRYB[14][47] , \CARRYB[14][46] ,
         \CARRYB[14][45] , \CARRYB[14][44] , \CARRYB[14][43] ,
         \CARRYB[14][42] , \CARRYB[14][41] , \CARRYB[14][40] ,
         \CARRYB[14][39] , \CARRYB[14][38] , \CARRYB[14][37] ,
         \CARRYB[14][36] , \CARRYB[14][35] , \CARRYB[14][34] ,
         \CARRYB[14][33] , \CARRYB[14][32] , \CARRYB[14][31] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \SUMB[19][31] , \SUMB[19][30] , \SUMB[19][29] ,
         \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] , \SUMB[19][25] ,
         \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] , \SUMB[19][21] ,
         \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] ,
         \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] ,
         \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] ,
         \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] ,
         \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] ,
         \SUMB[18][94] , \SUMB[18][93] , \SUMB[18][92] , \SUMB[18][91] ,
         \SUMB[18][90] , \SUMB[18][89] , \SUMB[18][88] , \SUMB[18][87] ,
         \SUMB[18][86] , \SUMB[18][85] , \SUMB[18][84] , \SUMB[18][83] ,
         \SUMB[18][82] , \SUMB[18][81] , \SUMB[18][80] , \SUMB[18][79] ,
         \SUMB[18][78] , \SUMB[18][77] , \SUMB[18][76] , \SUMB[18][75] ,
         \SUMB[18][74] , \SUMB[18][73] , \SUMB[18][72] , \SUMB[18][71] ,
         \SUMB[18][70] , \SUMB[18][69] , \SUMB[18][68] , \SUMB[18][67] ,
         \SUMB[18][66] , \SUMB[18][65] , \SUMB[18][64] , \SUMB[18][63] ,
         \SUMB[18][62] , \SUMB[18][61] , \SUMB[18][60] , \SUMB[18][59] ,
         \SUMB[18][58] , \SUMB[18][57] , \SUMB[18][56] , \SUMB[18][55] ,
         \SUMB[18][54] , \SUMB[18][53] , \SUMB[18][52] , \SUMB[18][51] ,
         \SUMB[18][50] , \SUMB[18][49] , \SUMB[18][48] , \SUMB[18][47] ,
         \SUMB[18][46] , \SUMB[18][45] , \SUMB[18][44] , \SUMB[18][43] ,
         \SUMB[18][42] , \SUMB[18][41] , \SUMB[18][40] , \SUMB[18][39] ,
         \SUMB[18][38] , \SUMB[18][37] , \SUMB[18][36] , \SUMB[18][35] ,
         \SUMB[18][34] , \SUMB[18][33] , \SUMB[18][32] , \SUMB[18][31] ,
         \SUMB[18][30] , \SUMB[18][29] , \SUMB[18][28] , \SUMB[18][27] ,
         \SUMB[18][26] , \SUMB[18][25] , \SUMB[18][24] , \SUMB[18][23] ,
         \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] ,
         \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] ,
         \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] ,
         \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] ,
         \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][94] , \SUMB[17][93] ,
         \SUMB[17][92] , \SUMB[17][91] , \SUMB[17][90] , \SUMB[17][89] ,
         \SUMB[17][88] , \SUMB[17][87] , \SUMB[17][86] , \SUMB[17][85] ,
         \SUMB[17][84] , \SUMB[17][83] , \SUMB[17][82] , \SUMB[17][81] ,
         \SUMB[17][80] , \SUMB[17][79] , \SUMB[17][78] , \SUMB[17][77] ,
         \SUMB[17][76] , \SUMB[17][75] , \SUMB[17][74] , \SUMB[17][73] ,
         \SUMB[17][72] , \SUMB[17][71] , \SUMB[17][70] , \SUMB[17][69] ,
         \SUMB[17][68] , \SUMB[17][67] , \SUMB[17][66] , \SUMB[17][65] ,
         \SUMB[17][64] , \SUMB[17][63] , \SUMB[17][62] , \SUMB[17][61] ,
         \SUMB[17][60] , \SUMB[17][59] , \SUMB[17][58] , \SUMB[17][57] ,
         \SUMB[17][56] , \SUMB[17][55] , \SUMB[17][54] , \SUMB[17][53] ,
         \SUMB[17][52] , \SUMB[17][51] , \SUMB[17][50] , \SUMB[17][49] ,
         \SUMB[17][48] , \SUMB[17][47] , \SUMB[17][46] , \SUMB[17][45] ,
         \SUMB[17][44] , \SUMB[17][43] , \SUMB[17][42] , \SUMB[17][41] ,
         \SUMB[17][40] , \SUMB[17][39] , \SUMB[17][38] , \SUMB[17][37] ,
         \SUMB[17][36] , \SUMB[17][35] , \SUMB[17][34] , \SUMB[17][33] ,
         \SUMB[17][32] , \SUMB[17][31] , \SUMB[17][30] , \SUMB[17][29] ,
         \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] , \SUMB[17][25] ,
         \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] , \SUMB[17][21] ,
         \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] ,
         \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][94] , \SUMB[16][93] , \SUMB[16][92] , \SUMB[16][91] ,
         \SUMB[16][90] , \SUMB[16][89] , \SUMB[16][88] , \SUMB[16][87] ,
         \SUMB[16][86] , \SUMB[16][85] , \SUMB[16][84] , \SUMB[16][83] ,
         \SUMB[16][82] , \SUMB[16][81] , \SUMB[16][80] , \SUMB[16][79] ,
         \SUMB[16][78] , \SUMB[16][77] , \SUMB[16][76] , \SUMB[16][75] ,
         \SUMB[16][74] , \SUMB[16][73] , \SUMB[16][72] , \SUMB[16][71] ,
         \SUMB[16][70] , \SUMB[16][69] , \SUMB[16][68] , \SUMB[16][67] ,
         \SUMB[16][66] , \SUMB[16][65] , \SUMB[16][64] , \SUMB[16][63] ,
         \SUMB[16][62] , \SUMB[16][61] , \SUMB[16][60] , \SUMB[16][59] ,
         \SUMB[16][58] , \SUMB[16][57] , \SUMB[16][56] , \SUMB[16][55] ,
         \SUMB[16][54] , \SUMB[16][53] , \SUMB[16][52] , \SUMB[16][51] ,
         \SUMB[16][50] , \SUMB[16][49] , \SUMB[16][48] , \SUMB[16][47] ,
         \SUMB[16][46] , \SUMB[16][45] , \SUMB[16][44] , \SUMB[16][43] ,
         \SUMB[16][42] , \SUMB[16][41] , \SUMB[16][40] , \SUMB[16][39] ,
         \SUMB[16][38] , \SUMB[16][37] , \SUMB[16][36] , \SUMB[16][35] ,
         \SUMB[16][34] , \SUMB[16][33] , \SUMB[16][32] , \SUMB[16][31] ,
         \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] , \SUMB[16][27] ,
         \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] , \SUMB[16][23] ,
         \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][19] ,
         \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] , \SUMB[16][15] ,
         \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] ,
         \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] ,
         \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] ,
         \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][94] , \SUMB[15][93] ,
         \SUMB[15][92] , \SUMB[15][91] , \SUMB[15][90] , \SUMB[15][89] ,
         \SUMB[15][88] , \SUMB[15][87] , \SUMB[15][86] , \SUMB[15][85] ,
         \SUMB[15][84] , \SUMB[15][83] , \SUMB[15][82] , \SUMB[15][81] ,
         \SUMB[15][80] , \SUMB[15][79] , \SUMB[15][78] , \SUMB[15][77] ,
         \SUMB[15][76] , \SUMB[15][75] , \SUMB[15][74] , \SUMB[15][73] ,
         \SUMB[15][72] , \SUMB[15][71] , \SUMB[15][70] , \SUMB[15][69] ,
         \SUMB[15][68] , \SUMB[15][67] , \SUMB[15][66] , \SUMB[15][65] ,
         \SUMB[15][64] , \SUMB[15][63] , \SUMB[15][62] , \SUMB[15][61] ,
         \SUMB[15][60] , \SUMB[15][59] , \SUMB[15][58] , \SUMB[15][57] ,
         \SUMB[15][56] , \SUMB[15][55] , \SUMB[15][54] , \SUMB[15][53] ,
         \SUMB[15][52] , \SUMB[15][51] , \SUMB[15][50] , \SUMB[15][49] ,
         \SUMB[15][48] , \SUMB[15][47] , \SUMB[15][46] , \SUMB[15][45] ,
         \SUMB[15][44] , \SUMB[15][43] , \SUMB[15][42] , \SUMB[15][41] ,
         \SUMB[15][40] , \SUMB[15][39] , \SUMB[15][38] , \SUMB[15][37] ,
         \SUMB[15][36] , \SUMB[15][35] , \SUMB[15][34] , \SUMB[15][33] ,
         \SUMB[15][32] , \SUMB[15][31] , \SUMB[15][30] , \SUMB[15][29] ,
         \SUMB[15][28] , \SUMB[15][27] , \SUMB[15][26] , \SUMB[15][25] ,
         \SUMB[15][24] , \SUMB[15][23] , \SUMB[15][22] , \SUMB[15][21] ,
         \SUMB[15][20] , \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] ,
         \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][94] , \SUMB[14][93] , \SUMB[14][92] , \SUMB[14][91] ,
         \SUMB[14][90] , \SUMB[14][89] , \SUMB[14][88] , \SUMB[14][87] ,
         \SUMB[14][86] , \SUMB[14][85] , \SUMB[14][84] , \SUMB[14][83] ,
         \SUMB[14][82] , \SUMB[14][81] , \SUMB[14][80] , \SUMB[14][79] ,
         \SUMB[14][78] , \SUMB[14][77] , \SUMB[14][76] , \SUMB[14][75] ,
         \SUMB[14][74] , \SUMB[14][73] , \SUMB[14][72] , \SUMB[14][71] ,
         \SUMB[14][70] , \SUMB[14][69] , \SUMB[14][68] , \SUMB[14][67] ,
         \SUMB[14][66] , \SUMB[14][65] , \SUMB[14][64] , \SUMB[14][63] ,
         \SUMB[14][62] , \SUMB[14][61] , \SUMB[14][60] , \SUMB[14][59] ,
         \SUMB[14][58] , \SUMB[14][57] , \SUMB[14][56] , \SUMB[14][55] ,
         \SUMB[14][54] , \SUMB[14][53] , \SUMB[14][52] , \SUMB[14][51] ,
         \SUMB[14][50] , \SUMB[14][49] , \SUMB[14][48] , \SUMB[14][47] ,
         \SUMB[14][46] , \SUMB[14][45] , \SUMB[14][44] , \SUMB[14][43] ,
         \SUMB[14][42] , \SUMB[14][41] , \SUMB[14][40] , \SUMB[14][39] ,
         \SUMB[14][38] , \SUMB[14][37] , \SUMB[14][36] , \SUMB[14][35] ,
         \SUMB[14][34] , \SUMB[14][33] , \SUMB[14][32] , \SUMB[14][31] ,
         \SUMB[14][30] , \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] ,
         \SUMB[14][26] , \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] ,
         \SUMB[14][22] , \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] ,
         \SUMB[14][18] , \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] ,
         \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] ,
         \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] ,
         \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] ,
         \SUMB[14][2] , \SUMB[14][1] , \CARRYB[24][63] , \CARRYB[24][62] ,
         \CARRYB[24][61] , \CARRYB[24][60] , \CARRYB[24][59] ,
         \CARRYB[24][58] , \CARRYB[24][57] , \CARRYB[24][56] ,
         \CARRYB[24][55] , \CARRYB[24][54] , \CARRYB[24][53] ,
         \CARRYB[24][52] , \CARRYB[24][51] , \CARRYB[24][50] ,
         \CARRYB[24][49] , \CARRYB[24][48] , \CARRYB[24][47] ,
         \CARRYB[24][46] , \CARRYB[24][45] , \CARRYB[24][44] ,
         \CARRYB[24][43] , \CARRYB[24][42] , \CARRYB[24][41] ,
         \CARRYB[24][40] , \CARRYB[24][39] , \CARRYB[24][38] ,
         \CARRYB[24][37] , \CARRYB[24][36] , \CARRYB[24][35] ,
         \CARRYB[24][34] , \CARRYB[24][33] , \CARRYB[24][32] ,
         \CARRYB[24][31] , \CARRYB[24][30] , \CARRYB[24][29] ,
         \CARRYB[24][28] , \CARRYB[24][27] , \CARRYB[24][26] ,
         \CARRYB[24][25] , \CARRYB[24][24] , \CARRYB[24][23] ,
         \CARRYB[24][22] , \CARRYB[24][21] , \CARRYB[24][20] ,
         \CARRYB[24][19] , \CARRYB[24][18] , \CARRYB[24][17] ,
         \CARRYB[24][16] , \CARRYB[24][15] , \CARRYB[24][14] ,
         \CARRYB[24][13] , \CARRYB[24][12] , \CARRYB[24][11] ,
         \CARRYB[24][10] , \CARRYB[24][9] , \CARRYB[24][8] , \CARRYB[24][7] ,
         \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][3] ,
         \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] , \CARRYB[23][94] ,
         \CARRYB[23][93] , \CARRYB[23][92] , \CARRYB[23][91] ,
         \CARRYB[23][90] , \CARRYB[23][89] , \CARRYB[23][88] ,
         \CARRYB[23][87] , \CARRYB[23][86] , \CARRYB[23][85] ,
         \CARRYB[23][84] , \CARRYB[23][83] , \CARRYB[23][82] ,
         \CARRYB[23][81] , \CARRYB[23][80] , \CARRYB[23][79] ,
         \CARRYB[23][78] , \CARRYB[23][77] , \CARRYB[23][76] ,
         \CARRYB[23][75] , \CARRYB[23][74] , \CARRYB[23][73] ,
         \CARRYB[23][72] , \CARRYB[23][71] , \CARRYB[23][70] ,
         \CARRYB[23][69] , \CARRYB[23][68] , \CARRYB[23][67] ,
         \CARRYB[23][66] , \CARRYB[23][65] , \CARRYB[23][64] ,
         \CARRYB[23][63] , \CARRYB[23][62] , \CARRYB[23][61] ,
         \CARRYB[23][60] , \CARRYB[23][59] , \CARRYB[23][58] ,
         \CARRYB[23][57] , \CARRYB[23][56] , \CARRYB[23][55] ,
         \CARRYB[23][54] , \CARRYB[23][53] , \CARRYB[23][52] ,
         \CARRYB[23][51] , \CARRYB[23][50] , \CARRYB[23][49] ,
         \CARRYB[23][48] , \CARRYB[23][47] , \CARRYB[23][46] ,
         \CARRYB[23][45] , \CARRYB[23][44] , \CARRYB[23][43] ,
         \CARRYB[23][42] , \CARRYB[23][41] , \CARRYB[23][40] ,
         \CARRYB[23][39] , \CARRYB[23][38] , \CARRYB[23][37] ,
         \CARRYB[23][36] , \CARRYB[23][35] , \CARRYB[23][34] ,
         \CARRYB[23][33] , \CARRYB[23][32] , \CARRYB[23][31] ,
         \CARRYB[23][30] , \CARRYB[23][29] , \CARRYB[23][28] ,
         \CARRYB[23][27] , \CARRYB[23][26] , \CARRYB[23][25] ,
         \CARRYB[23][24] , \CARRYB[23][23] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][94] , \CARRYB[22][93] , \CARRYB[22][92] ,
         \CARRYB[22][91] , \CARRYB[22][90] , \CARRYB[22][89] ,
         \CARRYB[22][88] , \CARRYB[22][87] , \CARRYB[22][86] ,
         \CARRYB[22][85] , \CARRYB[22][84] , \CARRYB[22][83] ,
         \CARRYB[22][82] , \CARRYB[22][81] , \CARRYB[22][80] ,
         \CARRYB[22][79] , \CARRYB[22][78] , \CARRYB[22][77] ,
         \CARRYB[22][76] , \CARRYB[22][75] , \CARRYB[22][74] ,
         \CARRYB[22][73] , \CARRYB[22][72] , \CARRYB[22][71] ,
         \CARRYB[22][70] , \CARRYB[22][69] , \CARRYB[22][68] ,
         \CARRYB[22][67] , \CARRYB[22][66] , \CARRYB[22][65] ,
         \CARRYB[22][64] , \CARRYB[22][63] , \CARRYB[22][62] ,
         \CARRYB[22][61] , \CARRYB[22][60] , \CARRYB[22][59] ,
         \CARRYB[22][58] , \CARRYB[22][57] , \CARRYB[22][56] ,
         \CARRYB[22][55] , \CARRYB[22][54] , \CARRYB[22][53] ,
         \CARRYB[22][52] , \CARRYB[22][51] , \CARRYB[22][50] ,
         \CARRYB[22][49] , \CARRYB[22][48] , \CARRYB[22][47] ,
         \CARRYB[22][46] , \CARRYB[22][45] , \CARRYB[22][44] ,
         \CARRYB[22][43] , \CARRYB[22][42] , \CARRYB[22][41] ,
         \CARRYB[22][40] , \CARRYB[22][39] , \CARRYB[22][38] ,
         \CARRYB[22][37] , \CARRYB[22][36] , \CARRYB[22][35] ,
         \CARRYB[22][34] , \CARRYB[22][33] , \CARRYB[22][32] ,
         \CARRYB[22][31] , \CARRYB[22][30] , \CARRYB[22][29] ,
         \CARRYB[22][28] , \CARRYB[22][27] , \CARRYB[22][26] ,
         \CARRYB[22][25] , \CARRYB[22][24] , \CARRYB[22][23] ,
         \CARRYB[22][22] , \CARRYB[22][21] , \CARRYB[22][20] ,
         \CARRYB[22][19] , \CARRYB[22][18] , \CARRYB[22][17] ,
         \CARRYB[22][16] , \CARRYB[22][15] , \CARRYB[22][14] ,
         \CARRYB[22][13] , \CARRYB[22][12] , \CARRYB[22][11] ,
         \CARRYB[22][10] , \CARRYB[22][9] , \CARRYB[22][8] , \CARRYB[22][7] ,
         \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][94] ,
         \CARRYB[21][93] , \CARRYB[21][92] , \CARRYB[21][91] ,
         \CARRYB[21][90] , \CARRYB[21][89] , \CARRYB[21][88] ,
         \CARRYB[21][87] , \CARRYB[21][86] , \CARRYB[21][85] ,
         \CARRYB[21][84] , \CARRYB[21][83] , \CARRYB[21][82] ,
         \CARRYB[21][81] , \CARRYB[21][80] , \CARRYB[21][79] ,
         \CARRYB[21][78] , \CARRYB[21][77] , \CARRYB[21][76] ,
         \CARRYB[21][75] , \CARRYB[21][74] , \CARRYB[21][73] ,
         \CARRYB[21][72] , \CARRYB[21][71] , \CARRYB[21][70] ,
         \CARRYB[21][69] , \CARRYB[21][68] , \CARRYB[21][67] ,
         \CARRYB[21][66] , \CARRYB[21][65] , \CARRYB[21][64] ,
         \CARRYB[21][63] , \CARRYB[21][62] , \CARRYB[21][61] ,
         \CARRYB[21][60] , \CARRYB[21][59] , \CARRYB[21][58] ,
         \CARRYB[21][57] , \CARRYB[21][56] , \CARRYB[21][55] ,
         \CARRYB[21][54] , \CARRYB[21][53] , \CARRYB[21][52] ,
         \CARRYB[21][51] , \CARRYB[21][50] , \CARRYB[21][49] ,
         \CARRYB[21][48] , \CARRYB[21][47] , \CARRYB[21][46] ,
         \CARRYB[21][45] , \CARRYB[21][44] , \CARRYB[21][43] ,
         \CARRYB[21][42] , \CARRYB[21][41] , \CARRYB[21][40] ,
         \CARRYB[21][39] , \CARRYB[21][38] , \CARRYB[21][37] ,
         \CARRYB[21][36] , \CARRYB[21][35] , \CARRYB[21][34] ,
         \CARRYB[21][33] , \CARRYB[21][32] , \CARRYB[21][31] ,
         \CARRYB[21][30] , \CARRYB[21][29] , \CARRYB[21][28] ,
         \CARRYB[21][27] , \CARRYB[21][26] , \CARRYB[21][25] ,
         \CARRYB[21][24] , \CARRYB[21][23] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][94] , \CARRYB[20][93] , \CARRYB[20][92] ,
         \CARRYB[20][91] , \CARRYB[20][90] , \CARRYB[20][89] ,
         \CARRYB[20][88] , \CARRYB[20][87] , \CARRYB[20][86] ,
         \CARRYB[20][85] , \CARRYB[20][84] , \CARRYB[20][83] ,
         \CARRYB[20][82] , \CARRYB[20][81] , \CARRYB[20][80] ,
         \CARRYB[20][79] , \CARRYB[20][78] , \CARRYB[20][77] ,
         \CARRYB[20][76] , \CARRYB[20][75] , \CARRYB[20][74] ,
         \CARRYB[20][73] , \CARRYB[20][72] , \CARRYB[20][71] ,
         \CARRYB[20][70] , \CARRYB[20][69] , \CARRYB[20][68] ,
         \CARRYB[20][67] , \CARRYB[20][66] , \CARRYB[20][65] ,
         \CARRYB[20][64] , \CARRYB[20][63] , \CARRYB[20][62] ,
         \CARRYB[20][61] , \CARRYB[20][60] , \CARRYB[20][59] ,
         \CARRYB[20][58] , \CARRYB[20][57] , \CARRYB[20][56] ,
         \CARRYB[20][55] , \CARRYB[20][54] , \CARRYB[20][53] ,
         \CARRYB[20][52] , \CARRYB[20][51] , \CARRYB[20][50] ,
         \CARRYB[20][49] , \CARRYB[20][48] , \CARRYB[20][47] ,
         \CARRYB[20][46] , \CARRYB[20][45] , \CARRYB[20][44] ,
         \CARRYB[20][43] , \CARRYB[20][42] , \CARRYB[20][41] ,
         \CARRYB[20][40] , \CARRYB[20][39] , \CARRYB[20][38] ,
         \CARRYB[20][37] , \CARRYB[20][36] , \CARRYB[20][35] ,
         \CARRYB[20][34] , \CARRYB[20][33] , \CARRYB[20][32] ,
         \CARRYB[20][31] , \CARRYB[20][30] , \CARRYB[20][29] ,
         \CARRYB[20][28] , \CARRYB[20][27] , \CARRYB[20][26] ,
         \CARRYB[20][25] , \CARRYB[20][24] , \CARRYB[20][23] ,
         \CARRYB[20][22] , \CARRYB[20][21] , \CARRYB[20][20] ,
         \CARRYB[20][19] , \CARRYB[20][18] , \CARRYB[20][17] ,
         \CARRYB[20][16] , \CARRYB[20][15] , \CARRYB[20][14] ,
         \CARRYB[20][13] , \CARRYB[20][12] , \CARRYB[20][11] ,
         \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] , \CARRYB[20][7] ,
         \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] , \CARRYB[20][3] ,
         \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] , \CARRYB[19][94] ,
         \CARRYB[19][93] , \CARRYB[19][92] , \CARRYB[19][91] ,
         \CARRYB[19][90] , \CARRYB[19][89] , \CARRYB[19][88] ,
         \CARRYB[19][87] , \CARRYB[19][86] , \CARRYB[19][85] ,
         \CARRYB[19][84] , \CARRYB[19][83] , \CARRYB[19][82] ,
         \CARRYB[19][81] , \CARRYB[19][80] , \CARRYB[19][79] ,
         \CARRYB[19][78] , \CARRYB[19][77] , \CARRYB[19][76] ,
         \CARRYB[19][75] , \CARRYB[19][74] , \CARRYB[19][73] ,
         \CARRYB[19][72] , \CARRYB[19][71] , \CARRYB[19][70] ,
         \CARRYB[19][69] , \CARRYB[19][68] , \CARRYB[19][67] ,
         \CARRYB[19][66] , \CARRYB[19][65] , \CARRYB[19][64] ,
         \CARRYB[19][63] , \CARRYB[19][62] , \CARRYB[19][61] ,
         \CARRYB[19][60] , \CARRYB[19][59] , \CARRYB[19][58] ,
         \CARRYB[19][57] , \CARRYB[19][56] , \CARRYB[19][55] ,
         \CARRYB[19][54] , \CARRYB[19][53] , \CARRYB[19][52] ,
         \CARRYB[19][51] , \CARRYB[19][50] , \CARRYB[19][49] ,
         \CARRYB[19][48] , \CARRYB[19][47] , \CARRYB[19][46] ,
         \CARRYB[19][45] , \CARRYB[19][44] , \CARRYB[19][43] ,
         \CARRYB[19][42] , \CARRYB[19][41] , \CARRYB[19][40] ,
         \CARRYB[19][39] , \CARRYB[19][38] , \CARRYB[19][37] ,
         \CARRYB[19][36] , \CARRYB[19][35] , \CARRYB[19][34] ,
         \CARRYB[19][33] , \CARRYB[19][32] , \SUMB[24][63] , \SUMB[24][62] ,
         \SUMB[24][61] , \SUMB[24][60] , \SUMB[24][59] , \SUMB[24][58] ,
         \SUMB[24][57] , \SUMB[24][56] , \SUMB[24][55] , \SUMB[24][54] ,
         \SUMB[24][53] , \SUMB[24][52] , \SUMB[24][51] , \SUMB[24][50] ,
         \SUMB[24][49] , \SUMB[24][48] , \SUMB[24][47] , \SUMB[24][46] ,
         \SUMB[24][45] , \SUMB[24][44] , \SUMB[24][43] , \SUMB[24][42] ,
         \SUMB[24][41] , \SUMB[24][40] , \SUMB[24][39] , \SUMB[24][38] ,
         \SUMB[24][37] , \SUMB[24][36] , \SUMB[24][35] , \SUMB[24][34] ,
         \SUMB[24][33] , \SUMB[24][32] , \SUMB[24][31] , \SUMB[24][30] ,
         \SUMB[24][29] , \SUMB[24][28] , \SUMB[24][27] , \SUMB[24][26] ,
         \SUMB[24][25] , \SUMB[24][24] , \SUMB[24][23] , \SUMB[24][22] ,
         \SUMB[24][21] , \SUMB[24][20] , \SUMB[24][19] , \SUMB[24][18] ,
         \SUMB[24][17] , \SUMB[24][16] , \SUMB[24][15] , \SUMB[24][14] ,
         \SUMB[24][13] , \SUMB[24][12] , \SUMB[24][11] , \SUMB[24][10] ,
         \SUMB[24][9] , \SUMB[24][8] , \SUMB[24][7] , \SUMB[24][6] ,
         \SUMB[24][5] , \SUMB[24][4] , \SUMB[24][3] , \SUMB[24][2] ,
         \SUMB[24][1] , \SUMB[23][94] , \SUMB[23][93] , \SUMB[23][92] ,
         \SUMB[23][91] , \SUMB[23][90] , \SUMB[23][89] , \SUMB[23][88] ,
         \SUMB[23][87] , \SUMB[23][86] , \SUMB[23][85] , \SUMB[23][84] ,
         \SUMB[23][83] , \SUMB[23][82] , \SUMB[23][81] , \SUMB[23][80] ,
         \SUMB[23][79] , \SUMB[23][78] , \SUMB[23][77] , \SUMB[23][76] ,
         \SUMB[23][75] , \SUMB[23][74] , \SUMB[23][73] , \SUMB[23][72] ,
         \SUMB[23][71] , \SUMB[23][70] , \SUMB[23][69] , \SUMB[23][68] ,
         \SUMB[23][67] , \SUMB[23][66] , \SUMB[23][65] , \SUMB[23][64] ,
         \SUMB[23][63] , \SUMB[23][62] , \SUMB[23][61] , \SUMB[23][60] ,
         \SUMB[23][59] , \SUMB[23][58] , \SUMB[23][57] , \SUMB[23][56] ,
         \SUMB[23][55] , \SUMB[23][54] , \SUMB[23][53] , \SUMB[23][52] ,
         \SUMB[23][51] , \SUMB[23][50] , \SUMB[23][49] , \SUMB[23][48] ,
         \SUMB[23][47] , \SUMB[23][46] , \SUMB[23][45] , \SUMB[23][44] ,
         \SUMB[23][43] , \SUMB[23][42] , \SUMB[23][41] , \SUMB[23][40] ,
         \SUMB[23][39] , \SUMB[23][38] , \SUMB[23][37] , \SUMB[23][36] ,
         \SUMB[23][35] , \SUMB[23][34] , \SUMB[23][33] , \SUMB[23][32] ,
         \SUMB[23][31] , \SUMB[23][30] , \SUMB[23][29] , \SUMB[23][28] ,
         \SUMB[23][27] , \SUMB[23][26] , \SUMB[23][25] , \SUMB[23][24] ,
         \SUMB[23][23] , \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] ,
         \SUMB[23][19] , \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] ,
         \SUMB[23][15] , \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] ,
         \SUMB[23][11] , \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] ,
         \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] ,
         \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][94] ,
         \SUMB[22][93] , \SUMB[22][92] , \SUMB[22][91] , \SUMB[22][90] ,
         \SUMB[22][89] , \SUMB[22][88] , \SUMB[22][87] , \SUMB[22][86] ,
         \SUMB[22][85] , \SUMB[22][84] , \SUMB[22][83] , \SUMB[22][82] ,
         \SUMB[22][81] , \SUMB[22][80] , \SUMB[22][79] , \SUMB[22][78] ,
         \SUMB[22][77] , \SUMB[22][76] , \SUMB[22][75] , \SUMB[22][74] ,
         \SUMB[22][73] , \SUMB[22][72] , \SUMB[22][71] , \SUMB[22][70] ,
         \SUMB[22][69] , \SUMB[22][68] , \SUMB[22][67] , \SUMB[22][66] ,
         \SUMB[22][65] , \SUMB[22][64] , \SUMB[22][63] , \SUMB[22][62] ,
         \SUMB[22][61] , \SUMB[22][60] , \SUMB[22][59] , \SUMB[22][58] ,
         \SUMB[22][57] , \SUMB[22][56] , \SUMB[22][55] , \SUMB[22][54] ,
         \SUMB[22][53] , \SUMB[22][52] , \SUMB[22][51] , \SUMB[22][50] ,
         \SUMB[22][49] , \SUMB[22][48] , \SUMB[22][47] , \SUMB[22][46] ,
         \SUMB[22][45] , \SUMB[22][44] , \SUMB[22][43] , \SUMB[22][42] ,
         \SUMB[22][41] , \SUMB[22][40] , \SUMB[22][39] , \SUMB[22][38] ,
         \SUMB[22][37] , \SUMB[22][36] , \SUMB[22][35] , \SUMB[22][34] ,
         \SUMB[22][33] , \SUMB[22][32] , \SUMB[22][31] , \SUMB[22][30] ,
         \SUMB[22][29] , \SUMB[22][28] , \SUMB[22][27] , \SUMB[22][26] ,
         \SUMB[22][25] , \SUMB[22][24] , \SUMB[22][23] , \SUMB[22][22] ,
         \SUMB[22][21] , \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] ,
         \SUMB[22][17] , \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] ,
         \SUMB[22][13] , \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] ,
         \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] ,
         \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] ,
         \SUMB[22][1] , \SUMB[21][94] , \SUMB[21][93] , \SUMB[21][92] ,
         \SUMB[21][91] , \SUMB[21][90] , \SUMB[21][89] , \SUMB[21][88] ,
         \SUMB[21][87] , \SUMB[21][86] , \SUMB[21][85] , \SUMB[21][84] ,
         \SUMB[21][83] , \SUMB[21][82] , \SUMB[21][81] , \SUMB[21][80] ,
         \SUMB[21][79] , \SUMB[21][78] , \SUMB[21][77] , \SUMB[21][76] ,
         \SUMB[21][75] , \SUMB[21][74] , \SUMB[21][73] , \SUMB[21][72] ,
         \SUMB[21][71] , \SUMB[21][70] , \SUMB[21][69] , \SUMB[21][68] ,
         \SUMB[21][67] , \SUMB[21][66] , \SUMB[21][65] , \SUMB[21][64] ,
         \SUMB[21][63] , \SUMB[21][62] , \SUMB[21][61] , \SUMB[21][60] ,
         \SUMB[21][59] , \SUMB[21][58] , \SUMB[21][57] , \SUMB[21][56] ,
         \SUMB[21][55] , \SUMB[21][54] , \SUMB[21][53] , \SUMB[21][52] ,
         \SUMB[21][51] , \SUMB[21][50] , \SUMB[21][49] , \SUMB[21][48] ,
         \SUMB[21][47] , \SUMB[21][46] , \SUMB[21][45] , \SUMB[21][44] ,
         \SUMB[21][43] , \SUMB[21][42] , \SUMB[21][41] , \SUMB[21][40] ,
         \SUMB[21][39] , \SUMB[21][38] , \SUMB[21][37] , \SUMB[21][36] ,
         \SUMB[21][35] , \SUMB[21][34] , \SUMB[21][33] , \SUMB[21][32] ,
         \SUMB[21][31] , \SUMB[21][30] , \SUMB[21][29] , \SUMB[21][28] ,
         \SUMB[21][27] , \SUMB[21][26] , \SUMB[21][25] , \SUMB[21][24] ,
         \SUMB[21][23] , \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] ,
         \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] ,
         \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] ,
         \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] ,
         \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] ,
         \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][94] ,
         \SUMB[20][93] , \SUMB[20][92] , \SUMB[20][91] , \SUMB[20][90] ,
         \SUMB[20][89] , \SUMB[20][88] , \SUMB[20][87] , \SUMB[20][86] ,
         \SUMB[20][85] , \SUMB[20][84] , \SUMB[20][83] , \SUMB[20][82] ,
         \SUMB[20][81] , \SUMB[20][80] , \SUMB[20][79] , \SUMB[20][78] ,
         \SUMB[20][77] , \SUMB[20][76] , \SUMB[20][75] , \SUMB[20][74] ,
         \SUMB[20][73] , \SUMB[20][72] , \SUMB[20][71] , \SUMB[20][70] ,
         \SUMB[20][69] , \SUMB[20][68] , \SUMB[20][67] , \SUMB[20][66] ,
         \SUMB[20][65] , \SUMB[20][64] , \SUMB[20][63] , \SUMB[20][62] ,
         \SUMB[20][61] , \SUMB[20][60] , \SUMB[20][59] , \SUMB[20][58] ,
         \SUMB[20][57] , \SUMB[20][56] , \SUMB[20][55] , \SUMB[20][54] ,
         \SUMB[20][53] , \SUMB[20][52] , \SUMB[20][51] , \SUMB[20][50] ,
         \SUMB[20][49] , \SUMB[20][48] , \SUMB[20][47] , \SUMB[20][46] ,
         \SUMB[20][45] , \SUMB[20][44] , \SUMB[20][43] , \SUMB[20][42] ,
         \SUMB[20][41] , \SUMB[20][40] , \SUMB[20][39] , \SUMB[20][38] ,
         \SUMB[20][37] , \SUMB[20][36] , \SUMB[20][35] , \SUMB[20][34] ,
         \SUMB[20][33] , \SUMB[20][32] , \SUMB[20][31] , \SUMB[20][30] ,
         \SUMB[20][29] , \SUMB[20][28] , \SUMB[20][27] , \SUMB[20][26] ,
         \SUMB[20][25] , \SUMB[20][24] , \SUMB[20][23] , \SUMB[20][22] ,
         \SUMB[20][21] , \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] ,
         \SUMB[20][17] , \SUMB[20][16] , \SUMB[20][15] , \SUMB[20][14] ,
         \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] , \SUMB[20][10] ,
         \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] ,
         \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] ,
         \SUMB[20][1] , \SUMB[19][94] , \SUMB[19][93] , \SUMB[19][92] ,
         \SUMB[19][91] , \SUMB[19][90] , \SUMB[19][89] , \SUMB[19][88] ,
         \SUMB[19][87] , \SUMB[19][86] , \SUMB[19][85] , \SUMB[19][84] ,
         \SUMB[19][83] , \SUMB[19][82] , \SUMB[19][81] , \SUMB[19][80] ,
         \SUMB[19][79] , \SUMB[19][78] , \SUMB[19][77] , \SUMB[19][76] ,
         \SUMB[19][75] , \SUMB[19][74] , \SUMB[19][73] , \SUMB[19][72] ,
         \SUMB[19][71] , \SUMB[19][70] , \SUMB[19][69] , \SUMB[19][68] ,
         \SUMB[19][67] , \SUMB[19][66] , \SUMB[19][65] , \SUMB[19][64] ,
         \SUMB[19][63] , \SUMB[19][62] , \SUMB[19][61] , \SUMB[19][60] ,
         \SUMB[19][59] , \SUMB[19][58] , \SUMB[19][57] , \SUMB[19][56] ,
         \SUMB[19][55] , \SUMB[19][54] , \SUMB[19][53] , \SUMB[19][52] ,
         \SUMB[19][51] , \SUMB[19][50] , \SUMB[19][49] , \SUMB[19][48] ,
         \SUMB[19][47] , \SUMB[19][46] , \SUMB[19][45] , \SUMB[19][44] ,
         \SUMB[19][43] , \SUMB[19][42] , \SUMB[19][41] , \SUMB[19][40] ,
         \SUMB[19][39] , \SUMB[19][38] , \SUMB[19][37] , \SUMB[19][36] ,
         \SUMB[19][35] , \SUMB[19][34] , \SUMB[19][33] , \SUMB[19][32] ,
         \CARRYB[29][94] , \CARRYB[29][93] , \CARRYB[29][92] ,
         \CARRYB[29][91] , \CARRYB[29][90] , \CARRYB[29][89] ,
         \CARRYB[29][88] , \CARRYB[29][87] , \CARRYB[29][86] ,
         \CARRYB[29][85] , \CARRYB[29][84] , \CARRYB[29][83] ,
         \CARRYB[29][82] , \CARRYB[29][81] , \CARRYB[29][80] ,
         \CARRYB[29][79] , \CARRYB[29][78] , \CARRYB[29][77] ,
         \CARRYB[29][76] , \CARRYB[29][75] , \CARRYB[29][74] ,
         \CARRYB[29][73] , \CARRYB[29][72] , \CARRYB[29][71] ,
         \CARRYB[29][70] , \CARRYB[29][69] , \CARRYB[29][68] ,
         \CARRYB[29][67] , \CARRYB[29][66] , \CARRYB[29][65] ,
         \CARRYB[29][64] , \CARRYB[29][63] , \CARRYB[29][62] ,
         \CARRYB[29][61] , \CARRYB[29][60] , \CARRYB[29][59] ,
         \CARRYB[29][58] , \CARRYB[29][57] , \CARRYB[29][56] ,
         \CARRYB[29][55] , \CARRYB[29][54] , \CARRYB[29][53] ,
         \CARRYB[29][52] , \CARRYB[29][51] , \CARRYB[29][50] ,
         \CARRYB[29][49] , \CARRYB[29][48] , \CARRYB[29][47] ,
         \CARRYB[29][46] , \CARRYB[29][45] , \CARRYB[29][44] ,
         \CARRYB[29][43] , \CARRYB[29][42] , \CARRYB[29][41] ,
         \CARRYB[29][40] , \CARRYB[29][39] , \CARRYB[29][38] ,
         \CARRYB[29][37] , \CARRYB[29][36] , \CARRYB[29][35] ,
         \CARRYB[29][34] , \CARRYB[29][33] , \CARRYB[29][32] ,
         \CARRYB[29][31] , \CARRYB[29][30] , \CARRYB[29][29] ,
         \CARRYB[29][28] , \CARRYB[29][27] , \CARRYB[29][26] ,
         \CARRYB[29][25] , \CARRYB[29][24] , \CARRYB[29][23] ,
         \CARRYB[29][22] , \CARRYB[29][21] , \CARRYB[29][20] ,
         \CARRYB[29][19] , \CARRYB[29][18] , \CARRYB[29][17] ,
         \CARRYB[29][16] , \CARRYB[29][15] , \CARRYB[29][14] ,
         \CARRYB[29][13] , \CARRYB[29][12] , \CARRYB[29][11] ,
         \CARRYB[29][10] , \CARRYB[29][9] , \CARRYB[29][8] , \CARRYB[29][7] ,
         \CARRYB[29][6] , \CARRYB[29][5] , \CARRYB[29][4] , \CARRYB[29][3] ,
         \CARRYB[29][2] , \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][94] ,
         \CARRYB[28][93] , \CARRYB[28][92] , \CARRYB[28][91] ,
         \CARRYB[28][90] , \CARRYB[28][89] , \CARRYB[28][88] ,
         \CARRYB[28][87] , \CARRYB[28][86] , \CARRYB[28][85] ,
         \CARRYB[28][84] , \CARRYB[28][83] , \CARRYB[28][82] ,
         \CARRYB[28][81] , \CARRYB[28][80] , \CARRYB[28][79] ,
         \CARRYB[28][78] , \CARRYB[28][77] , \CARRYB[28][76] ,
         \CARRYB[28][75] , \CARRYB[28][74] , \CARRYB[28][73] ,
         \CARRYB[28][72] , \CARRYB[28][71] , \CARRYB[28][70] ,
         \CARRYB[28][69] , \CARRYB[28][68] , \CARRYB[28][67] ,
         \CARRYB[28][66] , \CARRYB[28][65] , \CARRYB[28][64] ,
         \CARRYB[28][63] , \CARRYB[28][62] , \CARRYB[28][61] ,
         \CARRYB[28][60] , \CARRYB[28][59] , \CARRYB[28][58] ,
         \CARRYB[28][57] , \CARRYB[28][56] , \CARRYB[28][55] ,
         \CARRYB[28][54] , \CARRYB[28][53] , \CARRYB[28][52] ,
         \CARRYB[28][51] , \CARRYB[28][50] , \CARRYB[28][49] ,
         \CARRYB[28][48] , \CARRYB[28][47] , \CARRYB[28][46] ,
         \CARRYB[28][45] , \CARRYB[28][44] , \CARRYB[28][43] ,
         \CARRYB[28][42] , \CARRYB[28][41] , \CARRYB[28][40] ,
         \CARRYB[28][39] , \CARRYB[28][38] , \CARRYB[28][37] ,
         \CARRYB[28][36] , \CARRYB[28][35] , \CARRYB[28][34] ,
         \CARRYB[28][33] , \CARRYB[28][32] , \CARRYB[28][31] ,
         \CARRYB[28][30] , \CARRYB[28][29] , \CARRYB[28][28] ,
         \CARRYB[28][27] , \CARRYB[28][26] , \CARRYB[28][25] ,
         \CARRYB[28][24] , \CARRYB[28][23] , \CARRYB[28][22] ,
         \CARRYB[28][21] , \CARRYB[28][20] , \CARRYB[28][19] ,
         \CARRYB[28][18] , \CARRYB[28][17] , \CARRYB[28][16] ,
         \CARRYB[28][15] , \CARRYB[28][14] , \CARRYB[28][13] ,
         \CARRYB[28][12] , \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] ,
         \CARRYB[28][8] , \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] ,
         \CARRYB[28][4] , \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][94] , \CARRYB[27][93] , \CARRYB[27][92] ,
         \CARRYB[27][91] , \CARRYB[27][90] , \CARRYB[27][89] ,
         \CARRYB[27][88] , \CARRYB[27][87] , \CARRYB[27][86] ,
         \CARRYB[27][85] , \CARRYB[27][84] , \CARRYB[27][83] ,
         \CARRYB[27][82] , \CARRYB[27][81] , \CARRYB[27][80] ,
         \CARRYB[27][79] , \CARRYB[27][78] , \CARRYB[27][77] ,
         \CARRYB[27][76] , \CARRYB[27][75] , \CARRYB[27][74] ,
         \CARRYB[27][73] , \CARRYB[27][72] , \CARRYB[27][71] ,
         \CARRYB[27][70] , \CARRYB[27][69] , \CARRYB[27][68] ,
         \CARRYB[27][67] , \CARRYB[27][66] , \CARRYB[27][65] ,
         \CARRYB[27][64] , \CARRYB[27][63] , \CARRYB[27][62] ,
         \CARRYB[27][61] , \CARRYB[27][60] , \CARRYB[27][59] ,
         \CARRYB[27][58] , \CARRYB[27][57] , \CARRYB[27][56] ,
         \CARRYB[27][55] , \CARRYB[27][54] , \CARRYB[27][53] ,
         \CARRYB[27][52] , \CARRYB[27][51] , \CARRYB[27][50] ,
         \CARRYB[27][49] , \CARRYB[27][48] , \CARRYB[27][47] ,
         \CARRYB[27][46] , \CARRYB[27][45] , \CARRYB[27][44] ,
         \CARRYB[27][43] , \CARRYB[27][42] , \CARRYB[27][41] ,
         \CARRYB[27][40] , \CARRYB[27][39] , \CARRYB[27][38] ,
         \CARRYB[27][37] , \CARRYB[27][36] , \CARRYB[27][35] ,
         \CARRYB[27][34] , \CARRYB[27][33] , \CARRYB[27][32] ,
         \CARRYB[27][31] , \CARRYB[27][30] , \CARRYB[27][29] ,
         \CARRYB[27][28] , \CARRYB[27][27] , \CARRYB[27][26] ,
         \CARRYB[27][25] , \CARRYB[27][24] , \CARRYB[27][23] ,
         \CARRYB[27][22] , \CARRYB[27][21] , \CARRYB[27][20] ,
         \CARRYB[27][19] , \CARRYB[27][18] , \CARRYB[27][17] ,
         \CARRYB[27][16] , \CARRYB[27][15] , \CARRYB[27][14] ,
         \CARRYB[27][13] , \CARRYB[27][12] , \CARRYB[27][11] ,
         \CARRYB[27][10] , \CARRYB[27][9] , \CARRYB[27][8] , \CARRYB[27][7] ,
         \CARRYB[27][6] , \CARRYB[27][5] , \CARRYB[27][4] , \CARRYB[27][3] ,
         \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] , \CARRYB[26][94] ,
         \CARRYB[26][93] , \CARRYB[26][92] , \CARRYB[26][91] ,
         \CARRYB[26][90] , \CARRYB[26][89] , \CARRYB[26][88] ,
         \CARRYB[26][87] , \CARRYB[26][86] , \CARRYB[26][85] ,
         \CARRYB[26][84] , \CARRYB[26][83] , \CARRYB[26][82] ,
         \CARRYB[26][81] , \CARRYB[26][80] , \CARRYB[26][79] ,
         \CARRYB[26][78] , \CARRYB[26][77] , \CARRYB[26][76] ,
         \CARRYB[26][75] , \CARRYB[26][74] , \CARRYB[26][73] ,
         \CARRYB[26][72] , \CARRYB[26][71] , \CARRYB[26][70] ,
         \CARRYB[26][69] , \CARRYB[26][68] , \CARRYB[26][67] ,
         \CARRYB[26][66] , \CARRYB[26][65] , \CARRYB[26][64] ,
         \CARRYB[26][63] , \CARRYB[26][62] , \CARRYB[26][61] ,
         \CARRYB[26][60] , \CARRYB[26][59] , \CARRYB[26][58] ,
         \CARRYB[26][57] , \CARRYB[26][56] , \CARRYB[26][55] ,
         \CARRYB[26][54] , \CARRYB[26][53] , \CARRYB[26][52] ,
         \CARRYB[26][51] , \CARRYB[26][50] , \CARRYB[26][49] ,
         \CARRYB[26][48] , \CARRYB[26][47] , \CARRYB[26][46] ,
         \CARRYB[26][45] , \CARRYB[26][44] , \CARRYB[26][43] ,
         \CARRYB[26][42] , \CARRYB[26][41] , \CARRYB[26][40] ,
         \CARRYB[26][39] , \CARRYB[26][38] , \CARRYB[26][37] ,
         \CARRYB[26][36] , \CARRYB[26][35] , \CARRYB[26][34] ,
         \CARRYB[26][33] , \CARRYB[26][32] , \CARRYB[26][31] ,
         \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][94] , \CARRYB[25][93] , \CARRYB[25][92] ,
         \CARRYB[25][91] , \CARRYB[25][90] , \CARRYB[25][89] ,
         \CARRYB[25][88] , \CARRYB[25][87] , \CARRYB[25][86] ,
         \CARRYB[25][85] , \CARRYB[25][84] , \CARRYB[25][83] ,
         \CARRYB[25][82] , \CARRYB[25][81] , \CARRYB[25][80] ,
         \CARRYB[25][79] , \CARRYB[25][78] , \CARRYB[25][77] ,
         \CARRYB[25][76] , \CARRYB[25][75] , \CARRYB[25][74] ,
         \CARRYB[25][73] , \CARRYB[25][72] , \CARRYB[25][71] ,
         \CARRYB[25][70] , \CARRYB[25][69] , \CARRYB[25][68] ,
         \CARRYB[25][67] , \CARRYB[25][66] , \CARRYB[25][65] ,
         \CARRYB[25][64] , \CARRYB[25][63] , \CARRYB[25][62] ,
         \CARRYB[25][61] , \CARRYB[25][60] , \CARRYB[25][59] ,
         \CARRYB[25][58] , \CARRYB[25][57] , \CARRYB[25][56] ,
         \CARRYB[25][55] , \CARRYB[25][54] , \CARRYB[25][53] ,
         \CARRYB[25][52] , \CARRYB[25][51] , \CARRYB[25][50] ,
         \CARRYB[25][49] , \CARRYB[25][48] , \CARRYB[25][47] ,
         \CARRYB[25][46] , \CARRYB[25][45] , \CARRYB[25][44] ,
         \CARRYB[25][43] , \CARRYB[25][42] , \CARRYB[25][41] ,
         \CARRYB[25][40] , \CARRYB[25][39] , \CARRYB[25][38] ,
         \CARRYB[25][37] , \CARRYB[25][36] , \CARRYB[25][35] ,
         \CARRYB[25][34] , \CARRYB[25][33] , \CARRYB[25][32] ,
         \CARRYB[25][31] , \CARRYB[25][30] , \CARRYB[25][29] ,
         \CARRYB[25][28] , \CARRYB[25][27] , \CARRYB[25][26] ,
         \CARRYB[25][25] , \CARRYB[25][24] , \CARRYB[25][23] ,
         \CARRYB[25][22] , \CARRYB[25][21] , \CARRYB[25][20] ,
         \CARRYB[25][19] , \CARRYB[25][18] , \CARRYB[25][17] ,
         \CARRYB[25][16] , \CARRYB[25][15] , \CARRYB[25][14] ,
         \CARRYB[25][13] , \CARRYB[25][12] , \CARRYB[25][11] ,
         \CARRYB[25][10] , \CARRYB[25][9] , \CARRYB[25][8] , \CARRYB[25][7] ,
         \CARRYB[25][6] , \CARRYB[25][5] , \CARRYB[25][4] , \CARRYB[25][3] ,
         \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] , \CARRYB[24][94] ,
         \CARRYB[24][93] , \CARRYB[24][92] , \CARRYB[24][91] ,
         \CARRYB[24][90] , \CARRYB[24][89] , \CARRYB[24][88] ,
         \CARRYB[24][87] , \CARRYB[24][86] , \CARRYB[24][85] ,
         \CARRYB[24][84] , \CARRYB[24][83] , \CARRYB[24][82] ,
         \CARRYB[24][81] , \CARRYB[24][80] , \CARRYB[24][79] ,
         \CARRYB[24][78] , \CARRYB[24][77] , \CARRYB[24][76] ,
         \CARRYB[24][75] , \CARRYB[24][74] , \CARRYB[24][73] ,
         \CARRYB[24][72] , \CARRYB[24][71] , \CARRYB[24][70] ,
         \CARRYB[24][69] , \CARRYB[24][68] , \CARRYB[24][67] ,
         \CARRYB[24][66] , \CARRYB[24][65] , \CARRYB[24][64] , \SUMB[29][94] ,
         \SUMB[29][93] , \SUMB[29][92] , \SUMB[29][91] , \SUMB[29][90] ,
         \SUMB[29][89] , \SUMB[29][88] , \SUMB[29][87] , \SUMB[29][86] ,
         \SUMB[29][85] , \SUMB[29][84] , \SUMB[29][83] , \SUMB[29][82] ,
         \SUMB[29][81] , \SUMB[29][80] , \SUMB[29][79] , \SUMB[29][78] ,
         \SUMB[29][77] , \SUMB[29][76] , \SUMB[29][75] , \SUMB[29][74] ,
         \SUMB[29][73] , \SUMB[29][72] , \SUMB[29][71] , \SUMB[29][70] ,
         \SUMB[29][69] , \SUMB[29][68] , \SUMB[29][67] , \SUMB[29][66] ,
         \SUMB[29][65] , \SUMB[29][64] , \SUMB[29][63] , \SUMB[29][62] ,
         \SUMB[29][61] , \SUMB[29][60] , \SUMB[29][59] , \SUMB[29][58] ,
         \SUMB[29][57] , \SUMB[29][56] , \SUMB[29][55] , \SUMB[29][54] ,
         \SUMB[29][53] , \SUMB[29][52] , \SUMB[29][51] , \SUMB[29][50] ,
         \SUMB[29][49] , \SUMB[29][48] , \SUMB[29][47] , \SUMB[29][46] ,
         \SUMB[29][45] , \SUMB[29][44] , \SUMB[29][43] , \SUMB[29][42] ,
         \SUMB[29][41] , \SUMB[29][40] , \SUMB[29][39] , \SUMB[29][38] ,
         \SUMB[29][37] , \SUMB[29][36] , \SUMB[29][35] , \SUMB[29][34] ,
         \SUMB[29][33] , \SUMB[29][32] , \SUMB[29][31] , \SUMB[29][30] ,
         \SUMB[29][29] , \SUMB[29][28] , \SUMB[29][27] , \SUMB[29][26] ,
         \SUMB[29][25] , \SUMB[29][24] , \SUMB[29][23] , \SUMB[29][22] ,
         \SUMB[29][21] , \SUMB[29][20] , \SUMB[29][19] , \SUMB[29][18] ,
         \SUMB[29][17] , \SUMB[29][16] , \SUMB[29][15] , \SUMB[29][14] ,
         \SUMB[29][13] , \SUMB[29][12] , \SUMB[29][11] , \SUMB[29][10] ,
         \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] , \SUMB[29][6] ,
         \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] , \SUMB[29][2] ,
         \SUMB[29][1] , \SUMB[29][0] , \SUMB[28][94] , \SUMB[28][93] ,
         \SUMB[28][92] , \SUMB[28][91] , \SUMB[28][90] , \SUMB[28][89] ,
         \SUMB[28][88] , \SUMB[28][87] , \SUMB[28][86] , \SUMB[28][85] ,
         \SUMB[28][84] , \SUMB[28][83] , \SUMB[28][82] , \SUMB[28][81] ,
         \SUMB[28][80] , \SUMB[28][79] , \SUMB[28][78] , \SUMB[28][77] ,
         \SUMB[28][76] , \SUMB[28][75] , \SUMB[28][74] , \SUMB[28][73] ,
         \SUMB[28][72] , \SUMB[28][71] , \SUMB[28][70] , \SUMB[28][69] ,
         \SUMB[28][68] , \SUMB[28][67] , \SUMB[28][66] , \SUMB[28][65] ,
         \SUMB[28][64] , \SUMB[28][63] , \SUMB[28][62] , \SUMB[28][61] ,
         \SUMB[28][60] , \SUMB[28][59] , \SUMB[28][58] , \SUMB[28][57] ,
         \SUMB[28][56] , \SUMB[28][55] , \SUMB[28][54] , \SUMB[28][53] ,
         \SUMB[28][52] , \SUMB[28][51] , \SUMB[28][50] , \SUMB[28][49] ,
         \SUMB[28][48] , \SUMB[28][47] , \SUMB[28][46] , \SUMB[28][45] ,
         \SUMB[28][44] , \SUMB[28][43] , \SUMB[28][42] , \SUMB[28][41] ,
         \SUMB[28][40] , \SUMB[28][39] , \SUMB[28][38] , \SUMB[28][37] ,
         \SUMB[28][36] , \SUMB[28][35] , \SUMB[28][34] , \SUMB[28][33] ,
         \SUMB[28][32] , \SUMB[28][31] , \SUMB[28][30] , \SUMB[28][29] ,
         \SUMB[28][28] , \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] ,
         \SUMB[28][24] , \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] ,
         \SUMB[28][20] , \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] ,
         \SUMB[28][16] , \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] ,
         \SUMB[28][12] , \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] ,
         \SUMB[28][8] , \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] ,
         \SUMB[28][4] , \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] ,
         \SUMB[27][94] , \SUMB[27][93] , \SUMB[27][92] , \SUMB[27][91] ,
         \SUMB[27][90] , \SUMB[27][89] , \SUMB[27][88] , \SUMB[27][87] ,
         \SUMB[27][86] , \SUMB[27][85] , \SUMB[27][84] , \SUMB[27][83] ,
         \SUMB[27][82] , \SUMB[27][81] , \SUMB[27][80] , \SUMB[27][79] ,
         \SUMB[27][78] , \SUMB[27][77] , \SUMB[27][76] , \SUMB[27][75] ,
         \SUMB[27][74] , \SUMB[27][73] , \SUMB[27][72] , \SUMB[27][71] ,
         \SUMB[27][70] , \SUMB[27][69] , \SUMB[27][68] , \SUMB[27][67] ,
         \SUMB[27][66] , \SUMB[27][65] , \SUMB[27][64] , \SUMB[27][63] ,
         \SUMB[27][62] , \SUMB[27][61] , \SUMB[27][60] , \SUMB[27][59] ,
         \SUMB[27][58] , \SUMB[27][57] , \SUMB[27][56] , \SUMB[27][55] ,
         \SUMB[27][54] , \SUMB[27][53] , \SUMB[27][52] , \SUMB[27][51] ,
         \SUMB[27][50] , \SUMB[27][49] , \SUMB[27][48] , \SUMB[27][47] ,
         \SUMB[27][46] , \SUMB[27][45] , \SUMB[27][44] , \SUMB[27][43] ,
         \SUMB[27][42] , \SUMB[27][41] , \SUMB[27][40] , \SUMB[27][39] ,
         \SUMB[27][38] , \SUMB[27][37] , \SUMB[27][36] , \SUMB[27][35] ,
         \SUMB[27][34] , \SUMB[27][33] , \SUMB[27][32] , \SUMB[27][31] ,
         \SUMB[27][30] , \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] ,
         \SUMB[27][26] , \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] ,
         \SUMB[27][22] , \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] ,
         \SUMB[27][18] , \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] ,
         \SUMB[27][14] , \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] ,
         \SUMB[27][10] , \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] ,
         \SUMB[27][6] , \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][94] , \SUMB[26][93] ,
         \SUMB[26][92] , \SUMB[26][91] , \SUMB[26][90] , \SUMB[26][89] ,
         \SUMB[26][88] , \SUMB[26][87] , \SUMB[26][86] , \SUMB[26][85] ,
         \SUMB[26][84] , \SUMB[26][83] , \SUMB[26][82] , \SUMB[26][81] ,
         \SUMB[26][80] , \SUMB[26][79] , \SUMB[26][78] , \SUMB[26][77] ,
         \SUMB[26][76] , \SUMB[26][75] , \SUMB[26][74] , \SUMB[26][73] ,
         \SUMB[26][72] , \SUMB[26][71] , \SUMB[26][70] , \SUMB[26][69] ,
         \SUMB[26][68] , \SUMB[26][67] , \SUMB[26][66] , \SUMB[26][65] ,
         \SUMB[26][64] , \SUMB[26][63] , \SUMB[26][62] , \SUMB[26][61] ,
         \SUMB[26][60] , \SUMB[26][59] , \SUMB[26][58] , \SUMB[26][57] ,
         \SUMB[26][56] , \SUMB[26][55] , \SUMB[26][54] , \SUMB[26][53] ,
         \SUMB[26][52] , \SUMB[26][51] , \SUMB[26][50] , \SUMB[26][49] ,
         \SUMB[26][48] , \SUMB[26][47] , \SUMB[26][46] , \SUMB[26][45] ,
         \SUMB[26][44] , \SUMB[26][43] , \SUMB[26][42] , \SUMB[26][41] ,
         \SUMB[26][40] , \SUMB[26][39] , \SUMB[26][38] , \SUMB[26][37] ,
         \SUMB[26][36] , \SUMB[26][35] , \SUMB[26][34] , \SUMB[26][33] ,
         \SUMB[26][32] , \SUMB[26][31] , \SUMB[26][30] , \SUMB[26][29] ,
         \SUMB[26][28] , \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] ,
         \SUMB[26][24] , \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] ,
         \SUMB[26][20] , \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] ,
         \SUMB[26][16] , \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] ,
         \SUMB[26][12] , \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] ,
         \SUMB[26][8] , \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] ,
         \SUMB[26][4] , \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] ,
         \SUMB[25][94] , \SUMB[25][93] , \SUMB[25][92] , \SUMB[25][91] ,
         \SUMB[25][90] , \SUMB[25][89] , \SUMB[25][88] , \SUMB[25][87] ,
         \SUMB[25][86] , \SUMB[25][85] , \SUMB[25][84] , \SUMB[25][83] ,
         \SUMB[25][82] , \SUMB[25][81] , \SUMB[25][80] , \SUMB[25][79] ,
         \SUMB[25][78] , \SUMB[25][77] , \SUMB[25][76] , \SUMB[25][75] ,
         \SUMB[25][74] , \SUMB[25][73] , \SUMB[25][72] , \SUMB[25][71] ,
         \SUMB[25][70] , \SUMB[25][69] , \SUMB[25][68] , \SUMB[25][67] ,
         \SUMB[25][66] , \SUMB[25][65] , \SUMB[25][64] , \SUMB[25][63] ,
         \SUMB[25][62] , \SUMB[25][61] , \SUMB[25][60] , \SUMB[25][59] ,
         \SUMB[25][58] , \SUMB[25][57] , \SUMB[25][56] , \SUMB[25][55] ,
         \SUMB[25][54] , \SUMB[25][53] , \SUMB[25][52] , \SUMB[25][51] ,
         \SUMB[25][50] , \SUMB[25][49] , \SUMB[25][48] , \SUMB[25][47] ,
         \SUMB[25][46] , \SUMB[25][45] , \SUMB[25][44] , \SUMB[25][43] ,
         \SUMB[25][42] , \SUMB[25][41] , \SUMB[25][40] , \SUMB[25][39] ,
         \SUMB[25][38] , \SUMB[25][37] , \SUMB[25][36] , \SUMB[25][35] ,
         \SUMB[25][34] , \SUMB[25][33] , \SUMB[25][32] , \SUMB[25][31] ,
         \SUMB[25][30] , \SUMB[25][29] , \SUMB[25][28] , \SUMB[25][27] ,
         \SUMB[25][26] , \SUMB[25][25] , \SUMB[25][24] , \SUMB[25][23] ,
         \SUMB[25][22] , \SUMB[25][21] , \SUMB[25][20] , \SUMB[25][19] ,
         \SUMB[25][18] , \SUMB[25][17] , \SUMB[25][16] , \SUMB[25][15] ,
         \SUMB[25][14] , \SUMB[25][13] , \SUMB[25][12] , \SUMB[25][11] ,
         \SUMB[25][10] , \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] ,
         \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] ,
         \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][94] , \SUMB[24][93] ,
         \SUMB[24][92] , \SUMB[24][91] , \SUMB[24][90] , \SUMB[24][89] ,
         \SUMB[24][88] , \SUMB[24][87] , \SUMB[24][86] , \SUMB[24][85] ,
         \SUMB[24][84] , \SUMB[24][83] , \SUMB[24][82] , \SUMB[24][81] ,
         \SUMB[24][80] , \SUMB[24][79] , \SUMB[24][78] , \SUMB[24][77] ,
         \SUMB[24][76] , \SUMB[24][75] , \SUMB[24][74] , \SUMB[24][73] ,
         \SUMB[24][72] , \SUMB[24][71] , \SUMB[24][70] , \SUMB[24][69] ,
         \SUMB[24][68] , \SUMB[24][67] , \SUMB[24][66] , \SUMB[24][65] ,
         \SUMB[24][64] , \A1[122] , \A1[121] , \A1[120] , \A1[119] , \A1[118] ,
         \A1[117] , \A1[116] , \A1[115] , \A1[114] , \A1[113] , \A1[112] ,
         \A1[111] , \A1[110] , \A1[109] , \A1[108] , \A1[107] , \A1[106] ,
         \A1[105] , \A1[104] , \A1[103] , \A1[102] , \A1[101] , \A1[100] ,
         \A1[99] , \A1[98] , \A1[97] , \A1[96] , \A1[95] , \A1[94] , \A1[93] ,
         \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] ,
         \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] ,
         \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] ,
         \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] ,
         \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] ,
         \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] ,
         \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] ,
         \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] ,
         \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] ,
         \A1[29] , \A1[28] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[123] , \A2[122] , \A2[121] , \A2[120] , \A2[119] ,
         \A2[118] , \A2[117] , \A2[116] , \A2[115] , \A2[114] , \A2[113] ,
         \A2[112] , \A2[111] , \A2[110] , \A2[109] , \A2[108] , \A2[107] ,
         \A2[106] , \A2[105] , \A2[104] , \A2[103] , \A2[102] , \A2[101] ,
         \A2[100] , \A2[99] , \A2[98] , \A2[97] , \A2[96] , \A2[95] , \A2[94] ,
         \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] ,
         \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] ,
         \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] ,
         \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] ,
         \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] ,
         \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] ,
         \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         \A2[30] , \A2[29] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93;

  LOG_POLY_DW01_add_6 FS_1 ( .A({1'b0, \A1[122] , \A1[121] , \A1[120] , 
        \A1[119] , \A1[118] , \A1[117] , \A1[116] , \A1[115] , \A1[114] , 
        \A1[113] , \A1[112] , \A1[111] , \A1[110] , \A1[109] , \A1[108] , 
        \A1[107] , \A1[106] , \A1[105] , \A1[104] , \A1[103] , \A1[102] , 
        \A1[101] , \A1[100] , \A1[99] , \A1[98] , \A1[97] , \A1[96] , \A1[95] , 
        \A1[94] , \A1[93] , \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , 
        \A1[87] , \A1[86] , \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , 
        \A1[80] , \A1[79] , \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , 
        \A1[73] , \A1[72] , \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , 
        \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , 
        \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , 
        \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , 
        \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , 
        \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , 
        \A1[31] , \A1[30] , \A1[29] , \A1[28] , \SUMB[29][0] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , 
        \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , 
        \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[123] , 
        \A2[122] , \A2[121] , \A2[120] , \A2[119] , \A2[118] , \A2[117] , 
        \A2[116] , \A2[115] , \A2[114] , \A2[113] , \A2[112] , \A2[111] , 
        \A2[110] , \A2[109] , \A2[108] , \A2[107] , \A2[106] , \A2[105] , 
        \A2[104] , \A2[103] , \A2[102] , \A2[101] , \A2[100] , \A2[99] , 
        \A2[98] , \A2[97] , \A2[96] , \A2[95] , \A2[94] , \A2[93] , \A2[92] , 
        \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] , \A2[86] , \A2[85] , 
        \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] , \A2[79] , \A2[78] , 
        \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] , \A2[72] , \A2[71] , 
        \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] , \A2[65] , \A2[64] , 
        \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , \A2[57] , 
        \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , 
        \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] , \A2[44] , \A2[43] , 
        \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , 
        \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , \A2[29] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, PRODUCT[118:89], SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93}) );
  FA1A S2_14_57 ( .A(\ab[14][57] ), .B(\CARRYB[13][57] ), .CI(\SUMB[13][58] ), 
        .CO(\CARRYB[14][57] ), .S(\SUMB[14][57] ) );
  FA1A S2_13_57 ( .A(\ab[13][57] ), .B(\CARRYB[12][57] ), .CI(\SUMB[12][58] ), 
        .CO(\CARRYB[13][57] ), .S(\SUMB[13][57] ) );
  FA1A S2_12_57 ( .A(\ab[12][57] ), .B(\CARRYB[11][57] ), .CI(\SUMB[11][58] ), 
        .CO(\CARRYB[12][57] ), .S(\SUMB[12][57] ) );
  FA1A S2_11_57 ( .A(\ab[11][57] ), .B(\CARRYB[10][57] ), .CI(\SUMB[10][58] ), 
        .CO(\CARRYB[11][57] ), .S(\SUMB[11][57] ) );
  FA1A S2_10_57 ( .A(\ab[10][57] ), .B(\CARRYB[9][57] ), .CI(\SUMB[9][58] ), 
        .CO(\CARRYB[10][57] ), .S(\SUMB[10][57] ) );
  FA1A S2_9_57 ( .A(\ab[9][57] ), .B(\CARRYB[8][57] ), .CI(\SUMB[8][58] ), 
        .CO(\CARRYB[9][57] ), .S(\SUMB[9][57] ) );
  FA1A S2_8_57 ( .A(\ab[8][57] ), .B(\CARRYB[7][57] ), .CI(\SUMB[7][58] ), 
        .CO(\CARRYB[8][57] ), .S(\SUMB[8][57] ) );
  FA1A S2_7_57 ( .A(\ab[7][57] ), .B(\CARRYB[6][57] ), .CI(\SUMB[6][58] ), 
        .CO(\CARRYB[7][57] ), .S(\SUMB[7][57] ) );
  FA1A S2_6_57 ( .A(\ab[6][57] ), .B(\CARRYB[5][57] ), .CI(\SUMB[5][58] ), 
        .CO(\CARRYB[6][57] ), .S(\SUMB[6][57] ) );
  FA1A S2_5_57 ( .A(\ab[5][57] ), .B(\CARRYB[4][57] ), .CI(\SUMB[4][58] ), 
        .CO(\CARRYB[5][57] ), .S(\SUMB[5][57] ) );
  FA1A S2_4_57 ( .A(\ab[4][57] ), .B(\CARRYB[3][57] ), .CI(\SUMB[3][58] ), 
        .CO(\CARRYB[4][57] ), .S(\SUMB[4][57] ) );
  FA1A S2_3_57 ( .A(\ab[3][57] ), .B(\CARRYB[2][57] ), .CI(\SUMB[2][58] ), 
        .CO(\CARRYB[3][57] ), .S(\SUMB[3][57] ) );
  FA1A S2_2_57 ( .A(\ab[2][57] ), .B(\CARRYB[1][57] ), .CI(\SUMB[1][58] ), 
        .CO(\CARRYB[2][57] ), .S(\SUMB[2][57] ) );
  FA1A S2_14_56 ( .A(\ab[14][56] ), .B(\CARRYB[13][56] ), .CI(\SUMB[13][57] ), 
        .CO(\CARRYB[14][56] ), .S(\SUMB[14][56] ) );
  FA1A S2_14_54 ( .A(\ab[14][54] ), .B(\CARRYB[13][54] ), .CI(\SUMB[13][55] ), 
        .CO(\CARRYB[14][54] ), .S(\SUMB[14][54] ) );
  FA1A S2_14_53 ( .A(\ab[14][53] ), .B(\CARRYB[13][53] ), .CI(\SUMB[13][54] ), 
        .CO(\CARRYB[14][53] ), .S(\SUMB[14][53] ) );
  FA1A S2_14_59 ( .A(\ab[14][59] ), .B(\CARRYB[13][59] ), .CI(\SUMB[13][60] ), 
        .CO(\CARRYB[14][59] ), .S(\SUMB[14][59] ) );
  FA1A S2_14_58 ( .A(\ab[14][58] ), .B(\CARRYB[13][58] ), .CI(\SUMB[13][59] ), 
        .CO(\CARRYB[14][58] ), .S(\SUMB[14][58] ) );
  FA1A S2_13_58 ( .A(\ab[13][58] ), .B(\CARRYB[12][58] ), .CI(\SUMB[12][59] ), 
        .CO(\CARRYB[13][58] ), .S(\SUMB[13][58] ) );
  FA1A S2_13_56 ( .A(\ab[13][56] ), .B(\CARRYB[12][56] ), .CI(\SUMB[12][57] ), 
        .CO(\CARRYB[13][56] ), .S(\SUMB[13][56] ) );
  FA1A S2_13_54 ( .A(\ab[13][54] ), .B(\CARRYB[12][54] ), .CI(\SUMB[12][55] ), 
        .CO(\CARRYB[13][54] ), .S(\SUMB[13][54] ) );
  FA1A S2_13_53 ( .A(\ab[13][53] ), .B(\CARRYB[12][53] ), .CI(\SUMB[12][54] ), 
        .CO(\CARRYB[13][53] ), .S(\SUMB[13][53] ) );
  FA1A S2_13_59 ( .A(\ab[13][59] ), .B(\CARRYB[12][59] ), .CI(\SUMB[12][60] ), 
        .CO(\CARRYB[13][59] ), .S(\SUMB[13][59] ) );
  FA1A S2_12_59 ( .A(\ab[12][59] ), .B(\CARRYB[11][59] ), .CI(\SUMB[11][60] ), 
        .CO(\CARRYB[12][59] ), .S(\SUMB[12][59] ) );
  FA1A S2_12_58 ( .A(\ab[12][58] ), .B(\CARRYB[11][58] ), .CI(\SUMB[11][59] ), 
        .CO(\CARRYB[12][58] ), .S(\SUMB[12][58] ) );
  FA1A S2_12_56 ( .A(\ab[12][56] ), .B(\CARRYB[11][56] ), .CI(\SUMB[11][57] ), 
        .CO(\CARRYB[12][56] ), .S(\SUMB[12][56] ) );
  FA1A S2_12_54 ( .A(\ab[12][54] ), .B(\CARRYB[11][54] ), .CI(\SUMB[11][55] ), 
        .CO(\CARRYB[12][54] ), .S(\SUMB[12][54] ) );
  FA1A S2_12_53 ( .A(\ab[12][53] ), .B(\CARRYB[11][53] ), .CI(\SUMB[11][54] ), 
        .CO(\CARRYB[12][53] ), .S(\SUMB[12][53] ) );
  FA1A S2_11_59 ( .A(\ab[11][59] ), .B(\CARRYB[10][59] ), .CI(\SUMB[10][60] ), 
        .CO(\CARRYB[11][59] ), .S(\SUMB[11][59] ) );
  FA1A S2_11_58 ( .A(\ab[11][58] ), .B(\CARRYB[10][58] ), .CI(\SUMB[10][59] ), 
        .CO(\CARRYB[11][58] ), .S(\SUMB[11][58] ) );
  FA1A S2_11_56 ( .A(\ab[11][56] ), .B(\CARRYB[10][56] ), .CI(\SUMB[10][57] ), 
        .CO(\CARRYB[11][56] ), .S(\SUMB[11][56] ) );
  FA1A S2_11_54 ( .A(\ab[11][54] ), .B(\CARRYB[10][54] ), .CI(\SUMB[10][55] ), 
        .CO(\CARRYB[11][54] ), .S(\SUMB[11][54] ) );
  FA1A S2_11_53 ( .A(\ab[11][53] ), .B(\CARRYB[10][53] ), .CI(\SUMB[10][54] ), 
        .CO(\CARRYB[11][53] ), .S(\SUMB[11][53] ) );
  FA1A S2_10_59 ( .A(\ab[10][59] ), .B(\CARRYB[9][59] ), .CI(\SUMB[9][60] ), 
        .CO(\CARRYB[10][59] ), .S(\SUMB[10][59] ) );
  FA1A S2_10_58 ( .A(\ab[10][58] ), .B(\CARRYB[9][58] ), .CI(\SUMB[9][59] ), 
        .CO(\CARRYB[10][58] ), .S(\SUMB[10][58] ) );
  FA1A S2_10_56 ( .A(\ab[10][56] ), .B(\CARRYB[9][56] ), .CI(\SUMB[9][57] ), 
        .CO(\CARRYB[10][56] ), .S(\SUMB[10][56] ) );
  FA1A S2_10_54 ( .A(\ab[10][54] ), .B(\CARRYB[9][54] ), .CI(\SUMB[9][55] ), 
        .CO(\CARRYB[10][54] ), .S(\SUMB[10][54] ) );
  FA1A S2_10_53 ( .A(\ab[10][53] ), .B(\CARRYB[9][53] ), .CI(\SUMB[9][54] ), 
        .CO(\CARRYB[10][53] ), .S(\SUMB[10][53] ) );
  FA1A S2_9_59 ( .A(\ab[9][59] ), .B(\CARRYB[8][59] ), .CI(\SUMB[8][60] ), 
        .CO(\CARRYB[9][59] ), .S(\SUMB[9][59] ) );
  FA1A S2_9_58 ( .A(\ab[9][58] ), .B(\CARRYB[8][58] ), .CI(\SUMB[8][59] ), 
        .CO(\CARRYB[9][58] ), .S(\SUMB[9][58] ) );
  FA1A S2_9_56 ( .A(\ab[9][56] ), .B(\CARRYB[8][56] ), .CI(\SUMB[8][57] ), 
        .CO(\CARRYB[9][56] ), .S(\SUMB[9][56] ) );
  FA1A S2_9_54 ( .A(\ab[9][54] ), .B(\CARRYB[8][54] ), .CI(\SUMB[8][55] ), 
        .CO(\CARRYB[9][54] ), .S(\SUMB[9][54] ) );
  FA1A S2_9_53 ( .A(\ab[9][53] ), .B(\CARRYB[8][53] ), .CI(\SUMB[8][54] ), 
        .CO(\CARRYB[9][53] ), .S(\SUMB[9][53] ) );
  FA1A S2_8_59 ( .A(\ab[8][59] ), .B(\CARRYB[7][59] ), .CI(\SUMB[7][60] ), 
        .CO(\CARRYB[8][59] ), .S(\SUMB[8][59] ) );
  FA1A S2_8_58 ( .A(\ab[8][58] ), .B(\CARRYB[7][58] ), .CI(\SUMB[7][59] ), 
        .CO(\CARRYB[8][58] ), .S(\SUMB[8][58] ) );
  FA1A S2_8_56 ( .A(\ab[8][56] ), .B(\CARRYB[7][56] ), .CI(\SUMB[7][57] ), 
        .CO(\CARRYB[8][56] ), .S(\SUMB[8][56] ) );
  FA1A S2_8_54 ( .A(\ab[8][54] ), .B(\CARRYB[7][54] ), .CI(\SUMB[7][55] ), 
        .CO(\CARRYB[8][54] ), .S(\SUMB[8][54] ) );
  FA1A S2_8_53 ( .A(\ab[8][53] ), .B(\CARRYB[7][53] ), .CI(\SUMB[7][54] ), 
        .CO(\CARRYB[8][53] ), .S(\SUMB[8][53] ) );
  FA1A S2_7_59 ( .A(\ab[7][59] ), .B(\CARRYB[6][59] ), .CI(\SUMB[6][60] ), 
        .CO(\CARRYB[7][59] ), .S(\SUMB[7][59] ) );
  FA1A S2_7_58 ( .A(\ab[7][58] ), .B(\CARRYB[6][58] ), .CI(\SUMB[6][59] ), 
        .CO(\CARRYB[7][58] ), .S(\SUMB[7][58] ) );
  FA1A S2_7_56 ( .A(\ab[7][56] ), .B(\CARRYB[6][56] ), .CI(\SUMB[6][57] ), 
        .CO(\CARRYB[7][56] ), .S(\SUMB[7][56] ) );
  FA1A S2_7_54 ( .A(\ab[7][54] ), .B(\CARRYB[6][54] ), .CI(\SUMB[6][55] ), 
        .CO(\CARRYB[7][54] ), .S(\SUMB[7][54] ) );
  FA1A S2_7_53 ( .A(\ab[7][53] ), .B(\CARRYB[6][53] ), .CI(\SUMB[6][54] ), 
        .CO(\CARRYB[7][53] ), .S(\SUMB[7][53] ) );
  FA1A S2_6_59 ( .A(\ab[6][59] ), .B(\CARRYB[5][59] ), .CI(\SUMB[5][60] ), 
        .CO(\CARRYB[6][59] ), .S(\SUMB[6][59] ) );
  FA1A S2_6_58 ( .A(\ab[6][58] ), .B(\CARRYB[5][58] ), .CI(\SUMB[5][59] ), 
        .CO(\CARRYB[6][58] ), .S(\SUMB[6][58] ) );
  FA1A S2_6_56 ( .A(\ab[6][56] ), .B(\CARRYB[5][56] ), .CI(\SUMB[5][57] ), 
        .CO(\CARRYB[6][56] ), .S(\SUMB[6][56] ) );
  FA1A S2_6_54 ( .A(\ab[6][54] ), .B(\CARRYB[5][54] ), .CI(\SUMB[5][55] ), 
        .CO(\CARRYB[6][54] ), .S(\SUMB[6][54] ) );
  FA1A S2_6_53 ( .A(\ab[6][53] ), .B(\CARRYB[5][53] ), .CI(\SUMB[5][54] ), 
        .CO(\CARRYB[6][53] ), .S(\SUMB[6][53] ) );
  FA1A S2_5_59 ( .A(\ab[5][59] ), .B(\CARRYB[4][59] ), .CI(\SUMB[4][60] ), 
        .CO(\CARRYB[5][59] ), .S(\SUMB[5][59] ) );
  FA1A S2_5_58 ( .A(\ab[5][58] ), .B(\CARRYB[4][58] ), .CI(\SUMB[4][59] ), 
        .CO(\CARRYB[5][58] ), .S(\SUMB[5][58] ) );
  FA1A S2_5_56 ( .A(\ab[5][56] ), .B(\CARRYB[4][56] ), .CI(\SUMB[4][57] ), 
        .CO(\CARRYB[5][56] ), .S(\SUMB[5][56] ) );
  FA1A S2_5_54 ( .A(\ab[5][54] ), .B(\CARRYB[4][54] ), .CI(\SUMB[4][55] ), 
        .CO(\CARRYB[5][54] ), .S(\SUMB[5][54] ) );
  FA1A S2_5_53 ( .A(\ab[5][53] ), .B(\CARRYB[4][53] ), .CI(\SUMB[4][54] ), 
        .CO(\CARRYB[5][53] ), .S(\SUMB[5][53] ) );
  FA1A S2_4_59 ( .A(\ab[4][59] ), .B(\CARRYB[3][59] ), .CI(\SUMB[3][60] ), 
        .CO(\CARRYB[4][59] ), .S(\SUMB[4][59] ) );
  FA1A S2_4_58 ( .A(\ab[4][58] ), .B(\CARRYB[3][58] ), .CI(\SUMB[3][59] ), 
        .CO(\CARRYB[4][58] ), .S(\SUMB[4][58] ) );
  FA1A S2_4_56 ( .A(\ab[4][56] ), .B(\CARRYB[3][56] ), .CI(\SUMB[3][57] ), 
        .CO(\CARRYB[4][56] ), .S(\SUMB[4][56] ) );
  FA1A S2_4_54 ( .A(\ab[4][54] ), .B(\CARRYB[3][54] ), .CI(\SUMB[3][55] ), 
        .CO(\CARRYB[4][54] ), .S(\SUMB[4][54] ) );
  FA1A S2_4_53 ( .A(\ab[4][53] ), .B(\CARRYB[3][53] ), .CI(\SUMB[3][54] ), 
        .CO(\CARRYB[4][53] ), .S(\SUMB[4][53] ) );
  FA1A S2_3_59 ( .A(\ab[3][59] ), .B(\CARRYB[2][59] ), .CI(\SUMB[2][60] ), 
        .CO(\CARRYB[3][59] ), .S(\SUMB[3][59] ) );
  FA1A S2_3_58 ( .A(\ab[3][58] ), .B(\CARRYB[2][58] ), .CI(\SUMB[2][59] ), 
        .CO(\CARRYB[3][58] ), .S(\SUMB[3][58] ) );
  FA1A S2_3_56 ( .A(\ab[3][56] ), .B(\CARRYB[2][56] ), .CI(\SUMB[2][57] ), 
        .CO(\CARRYB[3][56] ), .S(\SUMB[3][56] ) );
  FA1A S2_3_54 ( .A(\ab[3][54] ), .B(\CARRYB[2][54] ), .CI(\SUMB[2][55] ), 
        .CO(\CARRYB[3][54] ), .S(\SUMB[3][54] ) );
  FA1A S2_3_53 ( .A(\ab[3][53] ), .B(\CARRYB[2][53] ), .CI(\SUMB[2][54] ), 
        .CO(\CARRYB[3][53] ), .S(\SUMB[3][53] ) );
  FA1A S2_2_59 ( .A(\ab[2][59] ), .B(\CARRYB[1][59] ), .CI(\SUMB[1][60] ), 
        .CO(\CARRYB[2][59] ), .S(\SUMB[2][59] ) );
  FA1A S2_2_58 ( .A(\ab[2][58] ), .B(\CARRYB[1][58] ), .CI(\SUMB[1][59] ), 
        .CO(\CARRYB[2][58] ), .S(\SUMB[2][58] ) );
  FA1A S2_2_56 ( .A(\ab[2][56] ), .B(\CARRYB[1][56] ), .CI(\SUMB[1][57] ), 
        .CO(\CARRYB[2][56] ), .S(\SUMB[2][56] ) );
  FA1A S2_2_54 ( .A(\ab[2][54] ), .B(\CARRYB[1][54] ), .CI(\SUMB[1][55] ), 
        .CO(\CARRYB[2][54] ), .S(\SUMB[2][54] ) );
  FA1A S2_2_53 ( .A(\ab[2][53] ), .B(\CARRYB[1][53] ), .CI(\SUMB[1][54] ), 
        .CO(\CARRYB[2][53] ), .S(\SUMB[2][53] ) );
  FA1A S2_14_52 ( .A(\ab[14][52] ), .B(\CARRYB[13][52] ), .CI(\SUMB[13][53] ), 
        .CO(\CARRYB[14][52] ), .S(\SUMB[14][52] ) );
  FA1A S2_14_44 ( .A(\ab[14][44] ), .B(\CARRYB[13][44] ), .CI(\SUMB[13][45] ), 
        .CO(\CARRYB[14][44] ), .S(\SUMB[14][44] ) );
  FA1A S2_14_43 ( .A(\ab[14][43] ), .B(\CARRYB[13][43] ), .CI(\SUMB[13][44] ), 
        .CO(\CARRYB[14][43] ), .S(\SUMB[14][43] ) );
  FA1A S2_14_42 ( .A(\ab[14][42] ), .B(\CARRYB[13][42] ), .CI(\SUMB[13][43] ), 
        .CO(\CARRYB[14][42] ), .S(\SUMB[14][42] ) );
  FA1A S2_14_41 ( .A(\ab[14][41] ), .B(\CARRYB[13][41] ), .CI(\SUMB[13][42] ), 
        .CO(\CARRYB[14][41] ), .S(\SUMB[14][41] ) );
  FA1A S2_13_52 ( .A(\ab[13][52] ), .B(\CARRYB[12][52] ), .CI(\SUMB[12][53] ), 
        .CO(\CARRYB[13][52] ), .S(\SUMB[13][52] ) );
  FA1A S2_13_44 ( .A(\ab[13][44] ), .B(\CARRYB[12][44] ), .CI(\SUMB[12][45] ), 
        .CO(\CARRYB[13][44] ), .S(\SUMB[13][44] ) );
  FA1A S2_13_43 ( .A(\ab[13][43] ), .B(\CARRYB[12][43] ), .CI(\SUMB[12][44] ), 
        .CO(\CARRYB[13][43] ), .S(\SUMB[13][43] ) );
  FA1A S2_13_42 ( .A(\ab[13][42] ), .B(\CARRYB[12][42] ), .CI(\SUMB[12][43] ), 
        .CO(\CARRYB[13][42] ), .S(\SUMB[13][42] ) );
  FA1A S2_14_39 ( .A(\ab[14][39] ), .B(\CARRYB[13][39] ), .CI(\SUMB[13][40] ), 
        .CO(\CARRYB[14][39] ), .S(\SUMB[14][39] ) );
  FA1A S2_14_40 ( .A(\ab[14][40] ), .B(\CARRYB[13][40] ), .CI(\SUMB[13][41] ), 
        .CO(\CARRYB[14][40] ), .S(\SUMB[14][40] ) );
  FA1A S2_12_52 ( .A(\ab[12][52] ), .B(\CARRYB[11][52] ), .CI(\SUMB[11][53] ), 
        .CO(\CARRYB[12][52] ), .S(\SUMB[12][52] ) );
  FA1A S2_12_44 ( .A(\ab[12][44] ), .B(\CARRYB[11][44] ), .CI(\SUMB[11][45] ), 
        .CO(\CARRYB[12][44] ), .S(\SUMB[12][44] ) );
  FA1A S2_12_43 ( .A(\ab[12][43] ), .B(\CARRYB[11][43] ), .CI(\SUMB[11][44] ), 
        .CO(\CARRYB[12][43] ), .S(\SUMB[12][43] ) );
  FA1A S2_13_40 ( .A(\ab[13][40] ), .B(\CARRYB[12][40] ), .CI(\SUMB[12][41] ), 
        .CO(\CARRYB[13][40] ), .S(\SUMB[13][40] ) );
  FA1A S2_13_41 ( .A(\ab[13][41] ), .B(\CARRYB[12][41] ), .CI(\SUMB[12][42] ), 
        .CO(\CARRYB[13][41] ), .S(\SUMB[13][41] ) );
  FA1A S2_11_52 ( .A(\ab[11][52] ), .B(\CARRYB[10][52] ), .CI(\SUMB[10][53] ), 
        .CO(\CARRYB[11][52] ), .S(\SUMB[11][52] ) );
  FA1A S2_11_44 ( .A(\ab[11][44] ), .B(\CARRYB[10][44] ), .CI(\SUMB[10][45] ), 
        .CO(\CARRYB[11][44] ), .S(\SUMB[11][44] ) );
  FA1A S2_12_41 ( .A(\ab[12][41] ), .B(\CARRYB[11][41] ), .CI(\SUMB[11][42] ), 
        .CO(\CARRYB[12][41] ), .S(\SUMB[12][41] ) );
  FA1A S2_12_42 ( .A(\ab[12][42] ), .B(\CARRYB[11][42] ), .CI(\SUMB[11][43] ), 
        .CO(\CARRYB[12][42] ), .S(\SUMB[12][42] ) );
  FA1A S2_13_39 ( .A(\ab[13][39] ), .B(\CARRYB[12][39] ), .CI(\SUMB[12][40] ), 
        .CO(\CARRYB[13][39] ), .S(\SUMB[13][39] ) );
  FA1A S2_10_52 ( .A(\ab[10][52] ), .B(\CARRYB[9][52] ), .CI(\SUMB[9][53] ), 
        .CO(\CARRYB[10][52] ), .S(\SUMB[10][52] ) );
  FA1A S2_11_42 ( .A(\ab[11][42] ), .B(\CARRYB[10][42] ), .CI(\SUMB[10][43] ), 
        .CO(\CARRYB[11][42] ), .S(\SUMB[11][42] ) );
  FA1A S2_11_43 ( .A(\ab[11][43] ), .B(\CARRYB[10][43] ), .CI(\SUMB[10][44] ), 
        .CO(\CARRYB[11][43] ), .S(\SUMB[11][43] ) );
  FA1A S2_12_40 ( .A(\ab[12][40] ), .B(\CARRYB[11][40] ), .CI(\SUMB[11][41] ), 
        .CO(\CARRYB[12][40] ), .S(\SUMB[12][40] ) );
  FA1A S2_12_39 ( .A(\ab[12][39] ), .B(\CARRYB[11][39] ), .CI(\SUMB[11][40] ), 
        .CO(\CARRYB[12][39] ), .S(\SUMB[12][39] ) );
  FA1A S2_9_52 ( .A(\ab[9][52] ), .B(\CARRYB[8][52] ), .CI(\SUMB[8][53] ), 
        .CO(\CARRYB[9][52] ), .S(\SUMB[9][52] ) );
  FA1A S2_10_43 ( .A(\ab[10][43] ), .B(\CARRYB[9][43] ), .CI(\SUMB[9][44] ), 
        .CO(\CARRYB[10][43] ), .S(\SUMB[10][43] ) );
  FA1A S2_10_44 ( .A(\ab[10][44] ), .B(\CARRYB[9][44] ), .CI(\SUMB[9][45] ), 
        .CO(\CARRYB[10][44] ), .S(\SUMB[10][44] ) );
  FA1A S2_11_41 ( .A(\ab[11][41] ), .B(\CARRYB[10][41] ), .CI(\SUMB[10][42] ), 
        .CO(\CARRYB[11][41] ), .S(\SUMB[11][41] ) );
  FA1A S2_11_40 ( .A(\ab[11][40] ), .B(\CARRYB[10][40] ), .CI(\SUMB[10][41] ), 
        .CO(\CARRYB[11][40] ), .S(\SUMB[11][40] ) );
  FA1A S2_11_39 ( .A(\ab[11][39] ), .B(\CARRYB[10][39] ), .CI(\SUMB[10][40] ), 
        .CO(\CARRYB[11][39] ), .S(\SUMB[11][39] ) );
  FA1A S2_8_52 ( .A(\ab[8][52] ), .B(\CARRYB[7][52] ), .CI(\SUMB[7][53] ), 
        .CO(\CARRYB[8][52] ), .S(\SUMB[8][52] ) );
  FA1A S2_9_44 ( .A(\ab[9][44] ), .B(\CARRYB[8][44] ), .CI(\SUMB[8][45] ), 
        .CO(\CARRYB[9][44] ), .S(\SUMB[9][44] ) );
  FA1A S2_10_42 ( .A(\ab[10][42] ), .B(\CARRYB[9][42] ), .CI(\SUMB[9][43] ), 
        .CO(\CARRYB[10][42] ), .S(\SUMB[10][42] ) );
  FA1A S2_10_41 ( .A(\ab[10][41] ), .B(\CARRYB[9][41] ), .CI(\SUMB[9][42] ), 
        .CO(\CARRYB[10][41] ), .S(\SUMB[10][41] ) );
  FA1A S2_10_40 ( .A(\ab[10][40] ), .B(\CARRYB[9][40] ), .CI(\SUMB[9][41] ), 
        .CO(\CARRYB[10][40] ), .S(\SUMB[10][40] ) );
  FA1A S2_10_39 ( .A(\ab[10][39] ), .B(\CARRYB[9][39] ), .CI(\SUMB[9][40] ), 
        .CO(\CARRYB[10][39] ), .S(\SUMB[10][39] ) );
  FA1A S2_7_52 ( .A(\ab[7][52] ), .B(\CARRYB[6][52] ), .CI(\SUMB[6][53] ), 
        .CO(\CARRYB[7][52] ), .S(\SUMB[7][52] ) );
  FA1A S2_9_43 ( .A(\ab[9][43] ), .B(\CARRYB[8][43] ), .CI(\SUMB[8][44] ), 
        .CO(\CARRYB[9][43] ), .S(\SUMB[9][43] ) );
  FA1A S2_9_42 ( .A(\ab[9][42] ), .B(\CARRYB[8][42] ), .CI(\SUMB[8][43] ), 
        .CO(\CARRYB[9][42] ), .S(\SUMB[9][42] ) );
  FA1A S2_9_41 ( .A(\ab[9][41] ), .B(\CARRYB[8][41] ), .CI(\SUMB[8][42] ), 
        .CO(\CARRYB[9][41] ), .S(\SUMB[9][41] ) );
  FA1A S2_9_40 ( .A(\ab[9][40] ), .B(\CARRYB[8][40] ), .CI(\SUMB[8][41] ), 
        .CO(\CARRYB[9][40] ), .S(\SUMB[9][40] ) );
  FA1A S2_9_39 ( .A(\ab[9][39] ), .B(\CARRYB[8][39] ), .CI(\SUMB[8][40] ), 
        .CO(\CARRYB[9][39] ), .S(\SUMB[9][39] ) );
  FA1A S2_6_52 ( .A(\ab[6][52] ), .B(\CARRYB[5][52] ), .CI(\SUMB[5][53] ), 
        .CO(\CARRYB[6][52] ), .S(\SUMB[6][52] ) );
  FA1A S2_8_44 ( .A(\ab[8][44] ), .B(\CARRYB[7][44] ), .CI(\SUMB[7][45] ), 
        .CO(\CARRYB[8][44] ), .S(\SUMB[8][44] ) );
  FA1A S2_8_43 ( .A(\ab[8][43] ), .B(\CARRYB[7][43] ), .CI(\SUMB[7][44] ), 
        .CO(\CARRYB[8][43] ), .S(\SUMB[8][43] ) );
  FA1A S2_8_42 ( .A(\ab[8][42] ), .B(\CARRYB[7][42] ), .CI(\SUMB[7][43] ), 
        .CO(\CARRYB[8][42] ), .S(\SUMB[8][42] ) );
  FA1A S2_8_41 ( .A(\ab[8][41] ), .B(\CARRYB[7][41] ), .CI(\SUMB[7][42] ), 
        .CO(\CARRYB[8][41] ), .S(\SUMB[8][41] ) );
  FA1A S2_8_40 ( .A(\ab[8][40] ), .B(\CARRYB[7][40] ), .CI(\SUMB[7][41] ), 
        .CO(\CARRYB[8][40] ), .S(\SUMB[8][40] ) );
  FA1A S2_8_39 ( .A(\ab[8][39] ), .B(\CARRYB[7][39] ), .CI(\SUMB[7][40] ), 
        .CO(\CARRYB[8][39] ), .S(\SUMB[8][39] ) );
  FA1A S2_5_52 ( .A(\ab[5][52] ), .B(\CARRYB[4][52] ), .CI(\SUMB[4][53] ), 
        .CO(\CARRYB[5][52] ), .S(\SUMB[5][52] ) );
  FA1A S2_7_44 ( .A(\ab[7][44] ), .B(\CARRYB[6][44] ), .CI(\SUMB[6][45] ), 
        .CO(\CARRYB[7][44] ), .S(\SUMB[7][44] ) );
  FA1A S2_7_43 ( .A(\ab[7][43] ), .B(\CARRYB[6][43] ), .CI(\SUMB[6][44] ), 
        .CO(\CARRYB[7][43] ), .S(\SUMB[7][43] ) );
  FA1A S2_7_42 ( .A(\ab[7][42] ), .B(\CARRYB[6][42] ), .CI(\SUMB[6][43] ), 
        .CO(\CARRYB[7][42] ), .S(\SUMB[7][42] ) );
  FA1A S2_7_41 ( .A(\ab[7][41] ), .B(\CARRYB[6][41] ), .CI(\SUMB[6][42] ), 
        .CO(\CARRYB[7][41] ), .S(\SUMB[7][41] ) );
  FA1A S2_7_40 ( .A(\ab[7][40] ), .B(\CARRYB[6][40] ), .CI(\SUMB[6][41] ), 
        .CO(\CARRYB[7][40] ), .S(\SUMB[7][40] ) );
  FA1A S2_7_39 ( .A(\ab[7][39] ), .B(\CARRYB[6][39] ), .CI(\SUMB[6][40] ), 
        .CO(\CARRYB[7][39] ), .S(\SUMB[7][39] ) );
  FA1A S2_4_52 ( .A(\ab[4][52] ), .B(\CARRYB[3][52] ), .CI(\SUMB[3][53] ), 
        .CO(\CARRYB[4][52] ), .S(\SUMB[4][52] ) );
  FA1A S2_6_44 ( .A(\ab[6][44] ), .B(\CARRYB[5][44] ), .CI(\SUMB[5][45] ), 
        .CO(\CARRYB[6][44] ), .S(\SUMB[6][44] ) );
  FA1A S2_6_43 ( .A(\ab[6][43] ), .B(\CARRYB[5][43] ), .CI(\SUMB[5][44] ), 
        .CO(\CARRYB[6][43] ), .S(\SUMB[6][43] ) );
  FA1A S2_6_42 ( .A(\ab[6][42] ), .B(\CARRYB[5][42] ), .CI(\SUMB[5][43] ), 
        .CO(\CARRYB[6][42] ), .S(\SUMB[6][42] ) );
  FA1A S2_6_41 ( .A(\ab[6][41] ), .B(\CARRYB[5][41] ), .CI(\SUMB[5][42] ), 
        .CO(\CARRYB[6][41] ), .S(\SUMB[6][41] ) );
  FA1A S2_6_40 ( .A(\ab[6][40] ), .B(\CARRYB[5][40] ), .CI(\SUMB[5][41] ), 
        .CO(\CARRYB[6][40] ), .S(\SUMB[6][40] ) );
  FA1A S2_6_39 ( .A(\ab[6][39] ), .B(\CARRYB[5][39] ), .CI(\SUMB[5][40] ), 
        .CO(\CARRYB[6][39] ), .S(\SUMB[6][39] ) );
  FA1A S2_3_52 ( .A(\ab[3][52] ), .B(\CARRYB[2][52] ), .CI(\SUMB[2][53] ), 
        .CO(\CARRYB[3][52] ), .S(\SUMB[3][52] ) );
  FA1A S2_5_44 ( .A(\ab[5][44] ), .B(\CARRYB[4][44] ), .CI(\SUMB[4][45] ), 
        .CO(\CARRYB[5][44] ), .S(\SUMB[5][44] ) );
  FA1A S2_5_43 ( .A(\ab[5][43] ), .B(\CARRYB[4][43] ), .CI(\SUMB[4][44] ), 
        .CO(\CARRYB[5][43] ), .S(\SUMB[5][43] ) );
  FA1A S2_5_42 ( .A(\ab[5][42] ), .B(\CARRYB[4][42] ), .CI(\SUMB[4][43] ), 
        .CO(\CARRYB[5][42] ), .S(\SUMB[5][42] ) );
  FA1A S2_5_41 ( .A(\ab[5][41] ), .B(\CARRYB[4][41] ), .CI(\SUMB[4][42] ), 
        .CO(\CARRYB[5][41] ), .S(\SUMB[5][41] ) );
  FA1A S2_5_40 ( .A(\ab[5][40] ), .B(\CARRYB[4][40] ), .CI(\SUMB[4][41] ), 
        .CO(\CARRYB[5][40] ), .S(\SUMB[5][40] ) );
  FA1A S2_5_39 ( .A(\ab[5][39] ), .B(\CARRYB[4][39] ), .CI(\SUMB[4][40] ), 
        .CO(\CARRYB[5][39] ), .S(\SUMB[5][39] ) );
  FA1A S2_4_44 ( .A(\ab[4][44] ), .B(\CARRYB[3][44] ), .CI(\SUMB[3][45] ), 
        .CO(\CARRYB[4][44] ), .S(\SUMB[4][44] ) );
  FA1A S2_4_43 ( .A(\ab[4][43] ), .B(\CARRYB[3][43] ), .CI(\SUMB[3][44] ), 
        .CO(\CARRYB[4][43] ), .S(\SUMB[4][43] ) );
  FA1A S2_4_42 ( .A(\ab[4][42] ), .B(\CARRYB[3][42] ), .CI(\SUMB[3][43] ), 
        .CO(\CARRYB[4][42] ), .S(\SUMB[4][42] ) );
  FA1A S2_4_41 ( .A(\ab[4][41] ), .B(\CARRYB[3][41] ), .CI(\SUMB[3][42] ), 
        .CO(\CARRYB[4][41] ), .S(\SUMB[4][41] ) );
  FA1A S2_4_40 ( .A(\ab[4][40] ), .B(\CARRYB[3][40] ), .CI(\SUMB[3][41] ), 
        .CO(\CARRYB[4][40] ), .S(\SUMB[4][40] ) );
  FA1A S2_4_39 ( .A(\ab[4][39] ), .B(\CARRYB[3][39] ), .CI(\SUMB[3][40] ), 
        .CO(\CARRYB[4][39] ), .S(\SUMB[4][39] ) );
  FA1A S2_2_52 ( .A(\ab[2][52] ), .B(\CARRYB[1][52] ), .CI(\SUMB[1][53] ), 
        .CO(\CARRYB[2][52] ), .S(\SUMB[2][52] ) );
  FA1A S2_3_44 ( .A(\ab[3][44] ), .B(\CARRYB[2][44] ), .CI(\SUMB[2][45] ), 
        .CO(\CARRYB[3][44] ), .S(\SUMB[3][44] ) );
  FA1A S2_3_43 ( .A(\ab[3][43] ), .B(\CARRYB[2][43] ), .CI(\SUMB[2][44] ), 
        .CO(\CARRYB[3][43] ), .S(\SUMB[3][43] ) );
  FA1A S2_3_42 ( .A(\ab[3][42] ), .B(\CARRYB[2][42] ), .CI(\SUMB[2][43] ), 
        .CO(\CARRYB[3][42] ), .S(\SUMB[3][42] ) );
  FA1A S2_3_41 ( .A(\ab[3][41] ), .B(\CARRYB[2][41] ), .CI(\SUMB[2][42] ), 
        .CO(\CARRYB[3][41] ), .S(\SUMB[3][41] ) );
  FA1A S2_3_40 ( .A(\ab[3][40] ), .B(\CARRYB[2][40] ), .CI(\SUMB[2][41] ), 
        .CO(\CARRYB[3][40] ), .S(\SUMB[3][40] ) );
  FA1A S2_3_39 ( .A(\ab[3][39] ), .B(\CARRYB[2][39] ), .CI(\SUMB[2][40] ), 
        .CO(\CARRYB[3][39] ), .S(\SUMB[3][39] ) );
  FA1A S2_2_44 ( .A(\ab[2][44] ), .B(\CARRYB[1][44] ), .CI(\SUMB[1][45] ), 
        .CO(\CARRYB[2][44] ), .S(\SUMB[2][44] ) );
  FA1A S2_2_43 ( .A(\ab[2][43] ), .B(\CARRYB[1][43] ), .CI(\SUMB[1][44] ), 
        .CO(\CARRYB[2][43] ), .S(\SUMB[2][43] ) );
  FA1A S2_2_42 ( .A(\ab[2][42] ), .B(\CARRYB[1][42] ), .CI(\SUMB[1][43] ), 
        .CO(\CARRYB[2][42] ), .S(\SUMB[2][42] ) );
  FA1A S2_2_41 ( .A(\ab[2][41] ), .B(\CARRYB[1][41] ), .CI(\SUMB[1][42] ), 
        .CO(\CARRYB[2][41] ), .S(\SUMB[2][41] ) );
  FA1A S2_2_40 ( .A(\ab[2][40] ), .B(\CARRYB[1][40] ), .CI(\SUMB[1][41] ), 
        .CO(\CARRYB[2][40] ), .S(\SUMB[2][40] ) );
  FA1A S2_2_39 ( .A(\ab[2][39] ), .B(\CARRYB[1][39] ), .CI(\SUMB[1][40] ), 
        .CO(\CARRYB[2][39] ), .S(\SUMB[2][39] ) );
  FA1A S2_14_51 ( .A(\ab[14][51] ), .B(\CARRYB[13][51] ), .CI(\SUMB[13][52] ), 
        .CO(\CARRYB[14][51] ), .S(\SUMB[14][51] ) );
  FA1A S2_14_50 ( .A(\ab[14][50] ), .B(\CARRYB[13][50] ), .CI(\SUMB[13][51] ), 
        .CO(\CARRYB[14][50] ), .S(\SUMB[14][50] ) );
  FA1A S2_14_49 ( .A(\ab[14][49] ), .B(\CARRYB[13][49] ), .CI(\SUMB[13][50] ), 
        .CO(\CARRYB[14][49] ), .S(\SUMB[14][49] ) );
  FA1A S2_14_48 ( .A(\ab[14][48] ), .B(\CARRYB[13][48] ), .CI(\SUMB[13][49] ), 
        .CO(\CARRYB[14][48] ), .S(\SUMB[14][48] ) );
  FA1A S2_14_47 ( .A(\ab[14][47] ), .B(\CARRYB[13][47] ), .CI(\SUMB[13][48] ), 
        .CO(\CARRYB[14][47] ), .S(\SUMB[14][47] ) );
  FA1A S2_14_46 ( .A(\ab[14][46] ), .B(\CARRYB[13][46] ), .CI(\SUMB[13][47] ), 
        .CO(\CARRYB[14][46] ), .S(\SUMB[14][46] ) );
  FA1A S2_14_45 ( .A(\ab[14][45] ), .B(\CARRYB[13][45] ), .CI(\SUMB[13][46] ), 
        .CO(\CARRYB[14][45] ), .S(\SUMB[14][45] ) );
  FA1A S2_13_51 ( .A(\ab[13][51] ), .B(\CARRYB[12][51] ), .CI(\SUMB[12][52] ), 
        .CO(\CARRYB[13][51] ), .S(\SUMB[13][51] ) );
  FA1A S2_13_50 ( .A(\ab[13][50] ), .B(\CARRYB[12][50] ), .CI(\SUMB[12][51] ), 
        .CO(\CARRYB[13][50] ), .S(\SUMB[13][50] ) );
  FA1A S2_13_49 ( .A(\ab[13][49] ), .B(\CARRYB[12][49] ), .CI(\SUMB[12][50] ), 
        .CO(\CARRYB[13][49] ), .S(\SUMB[13][49] ) );
  FA1A S2_13_48 ( .A(\ab[13][48] ), .B(\CARRYB[12][48] ), .CI(\SUMB[12][49] ), 
        .CO(\CARRYB[13][48] ), .S(\SUMB[13][48] ) );
  FA1A S2_13_47 ( .A(\ab[13][47] ), .B(\CARRYB[12][47] ), .CI(\SUMB[12][48] ), 
        .CO(\CARRYB[13][47] ), .S(\SUMB[13][47] ) );
  FA1A S2_13_46 ( .A(\ab[13][46] ), .B(\CARRYB[12][46] ), .CI(\SUMB[12][47] ), 
        .CO(\CARRYB[13][46] ), .S(\SUMB[13][46] ) );
  FA1A S2_13_45 ( .A(\ab[13][45] ), .B(\CARRYB[12][45] ), .CI(\SUMB[12][46] ), 
        .CO(\CARRYB[13][45] ), .S(\SUMB[13][45] ) );
  FA1A S2_12_51 ( .A(\ab[12][51] ), .B(\CARRYB[11][51] ), .CI(\SUMB[11][52] ), 
        .CO(\CARRYB[12][51] ), .S(\SUMB[12][51] ) );
  FA1A S2_12_50 ( .A(\ab[12][50] ), .B(\CARRYB[11][50] ), .CI(\SUMB[11][51] ), 
        .CO(\CARRYB[12][50] ), .S(\SUMB[12][50] ) );
  FA1A S2_12_49 ( .A(\ab[12][49] ), .B(\CARRYB[11][49] ), .CI(\SUMB[11][50] ), 
        .CO(\CARRYB[12][49] ), .S(\SUMB[12][49] ) );
  FA1A S2_12_48 ( .A(\ab[12][48] ), .B(\CARRYB[11][48] ), .CI(\SUMB[11][49] ), 
        .CO(\CARRYB[12][48] ), .S(\SUMB[12][48] ) );
  FA1A S2_12_47 ( .A(\ab[12][47] ), .B(\CARRYB[11][47] ), .CI(\SUMB[11][48] ), 
        .CO(\CARRYB[12][47] ), .S(\SUMB[12][47] ) );
  FA1A S2_12_46 ( .A(\ab[12][46] ), .B(\CARRYB[11][46] ), .CI(\SUMB[11][47] ), 
        .CO(\CARRYB[12][46] ), .S(\SUMB[12][46] ) );
  FA1A S2_12_45 ( .A(\ab[12][45] ), .B(\CARRYB[11][45] ), .CI(\SUMB[11][46] ), 
        .CO(\CARRYB[12][45] ), .S(\SUMB[12][45] ) );
  FA1A S2_11_51 ( .A(\ab[11][51] ), .B(\CARRYB[10][51] ), .CI(\SUMB[10][52] ), 
        .CO(\CARRYB[11][51] ), .S(\SUMB[11][51] ) );
  FA1A S2_11_50 ( .A(\ab[11][50] ), .B(\CARRYB[10][50] ), .CI(\SUMB[10][51] ), 
        .CO(\CARRYB[11][50] ), .S(\SUMB[11][50] ) );
  FA1A S2_11_49 ( .A(\ab[11][49] ), .B(\CARRYB[10][49] ), .CI(\SUMB[10][50] ), 
        .CO(\CARRYB[11][49] ), .S(\SUMB[11][49] ) );
  FA1A S2_11_48 ( .A(\ab[11][48] ), .B(\CARRYB[10][48] ), .CI(\SUMB[10][49] ), 
        .CO(\CARRYB[11][48] ), .S(\SUMB[11][48] ) );
  FA1A S2_11_47 ( .A(\ab[11][47] ), .B(\CARRYB[10][47] ), .CI(\SUMB[10][48] ), 
        .CO(\CARRYB[11][47] ), .S(\SUMB[11][47] ) );
  FA1A S2_11_46 ( .A(\ab[11][46] ), .B(\CARRYB[10][46] ), .CI(\SUMB[10][47] ), 
        .CO(\CARRYB[11][46] ), .S(\SUMB[11][46] ) );
  FA1A S2_11_45 ( .A(\ab[11][45] ), .B(\CARRYB[10][45] ), .CI(\SUMB[10][46] ), 
        .CO(\CARRYB[11][45] ), .S(\SUMB[11][45] ) );
  FA1A S2_10_51 ( .A(\ab[10][51] ), .B(\CARRYB[9][51] ), .CI(\SUMB[9][52] ), 
        .CO(\CARRYB[10][51] ), .S(\SUMB[10][51] ) );
  FA1A S2_10_50 ( .A(\ab[10][50] ), .B(\CARRYB[9][50] ), .CI(\SUMB[9][51] ), 
        .CO(\CARRYB[10][50] ), .S(\SUMB[10][50] ) );
  FA1A S2_10_49 ( .A(\ab[10][49] ), .B(\CARRYB[9][49] ), .CI(\SUMB[9][50] ), 
        .CO(\CARRYB[10][49] ), .S(\SUMB[10][49] ) );
  FA1A S2_10_48 ( .A(\ab[10][48] ), .B(\CARRYB[9][48] ), .CI(\SUMB[9][49] ), 
        .CO(\CARRYB[10][48] ), .S(\SUMB[10][48] ) );
  FA1A S2_10_47 ( .A(\ab[10][47] ), .B(\CARRYB[9][47] ), .CI(\SUMB[9][48] ), 
        .CO(\CARRYB[10][47] ), .S(\SUMB[10][47] ) );
  FA1A S2_10_46 ( .A(\ab[10][46] ), .B(\CARRYB[9][46] ), .CI(\SUMB[9][47] ), 
        .CO(\CARRYB[10][46] ), .S(\SUMB[10][46] ) );
  FA1A S2_10_45 ( .A(\ab[10][45] ), .B(\CARRYB[9][45] ), .CI(\SUMB[9][46] ), 
        .CO(\CARRYB[10][45] ), .S(\SUMB[10][45] ) );
  FA1A S2_9_51 ( .A(\ab[9][51] ), .B(\CARRYB[8][51] ), .CI(\SUMB[8][52] ), 
        .CO(\CARRYB[9][51] ), .S(\SUMB[9][51] ) );
  FA1A S2_9_50 ( .A(\ab[9][50] ), .B(\CARRYB[8][50] ), .CI(\SUMB[8][51] ), 
        .CO(\CARRYB[9][50] ), .S(\SUMB[9][50] ) );
  FA1A S2_9_49 ( .A(\ab[9][49] ), .B(\CARRYB[8][49] ), .CI(\SUMB[8][50] ), 
        .CO(\CARRYB[9][49] ), .S(\SUMB[9][49] ) );
  FA1A S2_9_48 ( .A(\ab[9][48] ), .B(\CARRYB[8][48] ), .CI(\SUMB[8][49] ), 
        .CO(\CARRYB[9][48] ), .S(\SUMB[9][48] ) );
  FA1A S2_9_47 ( .A(\ab[9][47] ), .B(\CARRYB[8][47] ), .CI(\SUMB[8][48] ), 
        .CO(\CARRYB[9][47] ), .S(\SUMB[9][47] ) );
  FA1A S2_9_46 ( .A(\ab[9][46] ), .B(\CARRYB[8][46] ), .CI(\SUMB[8][47] ), 
        .CO(\CARRYB[9][46] ), .S(\SUMB[9][46] ) );
  FA1A S2_8_51 ( .A(\ab[8][51] ), .B(\CARRYB[7][51] ), .CI(\SUMB[7][52] ), 
        .CO(\CARRYB[8][51] ), .S(\SUMB[8][51] ) );
  FA1A S2_8_50 ( .A(\ab[8][50] ), .B(\CARRYB[7][50] ), .CI(\SUMB[7][51] ), 
        .CO(\CARRYB[8][50] ), .S(\SUMB[8][50] ) );
  FA1A S2_8_49 ( .A(\ab[8][49] ), .B(\CARRYB[7][49] ), .CI(\SUMB[7][50] ), 
        .CO(\CARRYB[8][49] ), .S(\SUMB[8][49] ) );
  FA1A S2_8_48 ( .A(\ab[8][48] ), .B(\CARRYB[7][48] ), .CI(\SUMB[7][49] ), 
        .CO(\CARRYB[8][48] ), .S(\SUMB[8][48] ) );
  FA1A S2_8_47 ( .A(\ab[8][47] ), .B(\CARRYB[7][47] ), .CI(\SUMB[7][48] ), 
        .CO(\CARRYB[8][47] ), .S(\SUMB[8][47] ) );
  FA1A S2_9_45 ( .A(\ab[9][45] ), .B(\CARRYB[8][45] ), .CI(\SUMB[8][46] ), 
        .CO(\CARRYB[9][45] ), .S(\SUMB[9][45] ) );
  FA1A S2_7_51 ( .A(\ab[7][51] ), .B(\CARRYB[6][51] ), .CI(\SUMB[6][52] ), 
        .CO(\CARRYB[7][51] ), .S(\SUMB[7][51] ) );
  FA1A S2_7_50 ( .A(\ab[7][50] ), .B(\CARRYB[6][50] ), .CI(\SUMB[6][51] ), 
        .CO(\CARRYB[7][50] ), .S(\SUMB[7][50] ) );
  FA1A S2_7_49 ( .A(\ab[7][49] ), .B(\CARRYB[6][49] ), .CI(\SUMB[6][50] ), 
        .CO(\CARRYB[7][49] ), .S(\SUMB[7][49] ) );
  FA1A S2_7_48 ( .A(\ab[7][48] ), .B(\CARRYB[6][48] ), .CI(\SUMB[6][49] ), 
        .CO(\CARRYB[7][48] ), .S(\SUMB[7][48] ) );
  FA1A S2_8_45 ( .A(\ab[8][45] ), .B(\CARRYB[7][45] ), .CI(\SUMB[7][46] ), 
        .CO(\CARRYB[8][45] ), .S(\SUMB[8][45] ) );
  FA1A S2_8_46 ( .A(\ab[8][46] ), .B(\CARRYB[7][46] ), .CI(\SUMB[7][47] ), 
        .CO(\CARRYB[8][46] ), .S(\SUMB[8][46] ) );
  FA1A S2_6_51 ( .A(\ab[6][51] ), .B(\CARRYB[5][51] ), .CI(\SUMB[5][52] ), 
        .CO(\CARRYB[6][51] ), .S(\SUMB[6][51] ) );
  FA1A S2_6_50 ( .A(\ab[6][50] ), .B(\CARRYB[5][50] ), .CI(\SUMB[5][51] ), 
        .CO(\CARRYB[6][50] ), .S(\SUMB[6][50] ) );
  FA1A S2_6_49 ( .A(\ab[6][49] ), .B(\CARRYB[5][49] ), .CI(\SUMB[5][50] ), 
        .CO(\CARRYB[6][49] ), .S(\SUMB[6][49] ) );
  FA1A S2_7_46 ( .A(\ab[7][46] ), .B(\CARRYB[6][46] ), .CI(\SUMB[6][47] ), 
        .CO(\CARRYB[7][46] ), .S(\SUMB[7][46] ) );
  FA1A S2_7_47 ( .A(\ab[7][47] ), .B(\CARRYB[6][47] ), .CI(\SUMB[6][48] ), 
        .CO(\CARRYB[7][47] ), .S(\SUMB[7][47] ) );
  FA1A S2_5_51 ( .A(\ab[5][51] ), .B(\CARRYB[4][51] ), .CI(\SUMB[4][52] ), 
        .CO(\CARRYB[5][51] ), .S(\SUMB[5][51] ) );
  FA1A S2_5_50 ( .A(\ab[5][50] ), .B(\CARRYB[4][50] ), .CI(\SUMB[4][51] ), 
        .CO(\CARRYB[5][50] ), .S(\SUMB[5][50] ) );
  FA1A S2_6_47 ( .A(\ab[6][47] ), .B(\CARRYB[5][47] ), .CI(\SUMB[5][48] ), 
        .CO(\CARRYB[6][47] ), .S(\SUMB[6][47] ) );
  FA1A S2_6_48 ( .A(\ab[6][48] ), .B(\CARRYB[5][48] ), .CI(\SUMB[5][49] ), 
        .CO(\CARRYB[6][48] ), .S(\SUMB[6][48] ) );
  FA1A S2_7_45 ( .A(\ab[7][45] ), .B(\CARRYB[6][45] ), .CI(\SUMB[6][46] ), 
        .CO(\CARRYB[7][45] ), .S(\SUMB[7][45] ) );
  FA1A S2_4_51 ( .A(\ab[4][51] ), .B(\CARRYB[3][51] ), .CI(\SUMB[3][52] ), 
        .CO(\CARRYB[4][51] ), .S(\SUMB[4][51] ) );
  FA1A S2_5_48 ( .A(\ab[5][48] ), .B(\CARRYB[4][48] ), .CI(\SUMB[4][49] ), 
        .CO(\CARRYB[5][48] ), .S(\SUMB[5][48] ) );
  FA1A S2_5_49 ( .A(\ab[5][49] ), .B(\CARRYB[4][49] ), .CI(\SUMB[4][50] ), 
        .CO(\CARRYB[5][49] ), .S(\SUMB[5][49] ) );
  FA1A S2_6_46 ( .A(\ab[6][46] ), .B(\CARRYB[5][46] ), .CI(\SUMB[5][47] ), 
        .CO(\CARRYB[6][46] ), .S(\SUMB[6][46] ) );
  FA1A S2_6_45 ( .A(\ab[6][45] ), .B(\CARRYB[5][45] ), .CI(\SUMB[5][46] ), 
        .CO(\CARRYB[6][45] ), .S(\SUMB[6][45] ) );
  FA1A S2_4_49 ( .A(\ab[4][49] ), .B(\CARRYB[3][49] ), .CI(\SUMB[3][50] ), 
        .CO(\CARRYB[4][49] ), .S(\SUMB[4][49] ) );
  FA1A S2_4_50 ( .A(\ab[4][50] ), .B(\CARRYB[3][50] ), .CI(\SUMB[3][51] ), 
        .CO(\CARRYB[4][50] ), .S(\SUMB[4][50] ) );
  FA1A S2_5_47 ( .A(\ab[5][47] ), .B(\CARRYB[4][47] ), .CI(\SUMB[4][48] ), 
        .CO(\CARRYB[5][47] ), .S(\SUMB[5][47] ) );
  FA1A S2_5_46 ( .A(\ab[5][46] ), .B(\CARRYB[4][46] ), .CI(\SUMB[4][47] ), 
        .CO(\CARRYB[5][46] ), .S(\SUMB[5][46] ) );
  FA1A S2_5_45 ( .A(\ab[5][45] ), .B(\CARRYB[4][45] ), .CI(\SUMB[4][46] ), 
        .CO(\CARRYB[5][45] ), .S(\SUMB[5][45] ) );
  FA1A S2_3_50 ( .A(\ab[3][50] ), .B(\CARRYB[2][50] ), .CI(\SUMB[2][51] ), 
        .CO(\CARRYB[3][50] ), .S(\SUMB[3][50] ) );
  FA1A S2_3_51 ( .A(\ab[3][51] ), .B(\CARRYB[2][51] ), .CI(\SUMB[2][52] ), 
        .CO(\CARRYB[3][51] ), .S(\SUMB[3][51] ) );
  FA1A S2_4_48 ( .A(\ab[4][48] ), .B(\CARRYB[3][48] ), .CI(\SUMB[3][49] ), 
        .CO(\CARRYB[4][48] ), .S(\SUMB[4][48] ) );
  FA1A S2_4_47 ( .A(\ab[4][47] ), .B(\CARRYB[3][47] ), .CI(\SUMB[3][48] ), 
        .CO(\CARRYB[4][47] ), .S(\SUMB[4][47] ) );
  FA1A S2_4_46 ( .A(\ab[4][46] ), .B(\CARRYB[3][46] ), .CI(\SUMB[3][47] ), 
        .CO(\CARRYB[4][46] ), .S(\SUMB[4][46] ) );
  FA1A S2_4_45 ( .A(\ab[4][45] ), .B(\CARRYB[3][45] ), .CI(\SUMB[3][46] ), 
        .CO(\CARRYB[4][45] ), .S(\SUMB[4][45] ) );
  FA1A S2_2_51 ( .A(\ab[2][51] ), .B(\CARRYB[1][51] ), .CI(\SUMB[1][52] ), 
        .CO(\CARRYB[2][51] ), .S(\SUMB[2][51] ) );
  FA1A S2_3_49 ( .A(\ab[3][49] ), .B(\CARRYB[2][49] ), .CI(\SUMB[2][50] ), 
        .CO(\CARRYB[3][49] ), .S(\SUMB[3][49] ) );
  FA1A S2_3_48 ( .A(\ab[3][48] ), .B(\CARRYB[2][48] ), .CI(\SUMB[2][49] ), 
        .CO(\CARRYB[3][48] ), .S(\SUMB[3][48] ) );
  FA1A S2_3_47 ( .A(\ab[3][47] ), .B(\CARRYB[2][47] ), .CI(\SUMB[2][48] ), 
        .CO(\CARRYB[3][47] ), .S(\SUMB[3][47] ) );
  FA1A S2_3_46 ( .A(\ab[3][46] ), .B(\CARRYB[2][46] ), .CI(\SUMB[2][47] ), 
        .CO(\CARRYB[3][46] ), .S(\SUMB[3][46] ) );
  FA1A S2_3_45 ( .A(\ab[3][45] ), .B(\CARRYB[2][45] ), .CI(\SUMB[2][46] ), 
        .CO(\CARRYB[3][45] ), .S(\SUMB[3][45] ) );
  FA1A S2_2_50 ( .A(\ab[2][50] ), .B(\CARRYB[1][50] ), .CI(\SUMB[1][51] ), 
        .CO(\CARRYB[2][50] ), .S(\SUMB[2][50] ) );
  FA1A S2_2_49 ( .A(\ab[2][49] ), .B(\CARRYB[1][49] ), .CI(\SUMB[1][50] ), 
        .CO(\CARRYB[2][49] ), .S(\SUMB[2][49] ) );
  FA1A S2_2_48 ( .A(\ab[2][48] ), .B(\CARRYB[1][48] ), .CI(\SUMB[1][49] ), 
        .CO(\CARRYB[2][48] ), .S(\SUMB[2][48] ) );
  FA1A S2_2_47 ( .A(\ab[2][47] ), .B(\CARRYB[1][47] ), .CI(\SUMB[1][48] ), 
        .CO(\CARRYB[2][47] ), .S(\SUMB[2][47] ) );
  FA1A S2_2_46 ( .A(\ab[2][46] ), .B(\CARRYB[1][46] ), .CI(\SUMB[1][47] ), 
        .CO(\CARRYB[2][46] ), .S(\SUMB[2][46] ) );
  FA1A S2_2_45 ( .A(\ab[2][45] ), .B(\CARRYB[1][45] ), .CI(\SUMB[1][46] ), 
        .CO(\CARRYB[2][45] ), .S(\SUMB[2][45] ) );
  FA1A S5_94 ( .A(\ab[29][94] ), .B(\CARRYB[28][94] ), .CI(\ab[28][95] ), .CO(
        \CARRYB[29][94] ), .S(\SUMB[29][94] ) );
  FA1A S4_93 ( .A(\ab[29][93] ), .B(\CARRYB[28][93] ), .CI(\SUMB[28][94] ), 
        .CO(\CARRYB[29][93] ), .S(\SUMB[29][93] ) );
  FA1A S4_92 ( .A(\ab[29][92] ), .B(\CARRYB[28][92] ), .CI(\SUMB[28][93] ), 
        .CO(\CARRYB[29][92] ), .S(\SUMB[29][92] ) );
  FA1A S4_91 ( .A(\ab[29][91] ), .B(\CARRYB[28][91] ), .CI(\SUMB[28][92] ), 
        .CO(\CARRYB[29][91] ), .S(\SUMB[29][91] ) );
  FA1A S4_90 ( .A(\ab[29][90] ), .B(\CARRYB[28][90] ), .CI(\SUMB[28][91] ), 
        .CO(\CARRYB[29][90] ), .S(\SUMB[29][90] ) );
  FA1A S3_28_94 ( .A(\ab[28][94] ), .B(\CARRYB[27][94] ), .CI(\ab[27][95] ), 
        .CO(\CARRYB[28][94] ), .S(\SUMB[28][94] ) );
  FA1A S2_28_93 ( .A(\ab[28][93] ), .B(\CARRYB[27][93] ), .CI(\SUMB[27][94] ), 
        .CO(\CARRYB[28][93] ), .S(\SUMB[28][93] ) );
  FA1A S2_28_92 ( .A(\ab[28][92] ), .B(\CARRYB[27][92] ), .CI(\SUMB[27][93] ), 
        .CO(\CARRYB[28][92] ), .S(\SUMB[28][92] ) );
  FA1A S2_28_91 ( .A(\ab[28][91] ), .B(\CARRYB[27][91] ), .CI(\SUMB[27][92] ), 
        .CO(\CARRYB[28][91] ), .S(\SUMB[28][91] ) );
  FA1A S3_27_94 ( .A(\ab[27][94] ), .B(\CARRYB[26][94] ), .CI(\ab[26][95] ), 
        .CO(\CARRYB[27][94] ), .S(\SUMB[27][94] ) );
  FA1A S2_27_93 ( .A(\ab[27][93] ), .B(\CARRYB[26][93] ), .CI(\SUMB[26][94] ), 
        .CO(\CARRYB[27][93] ), .S(\SUMB[27][93] ) );
  FA1A S2_27_92 ( .A(\ab[27][92] ), .B(\CARRYB[26][92] ), .CI(\SUMB[26][93] ), 
        .CO(\CARRYB[27][92] ), .S(\SUMB[27][92] ) );
  FA1A S3_26_94 ( .A(\ab[26][94] ), .B(\CARRYB[25][94] ), .CI(\ab[25][95] ), 
        .CO(\CARRYB[26][94] ), .S(\SUMB[26][94] ) );
  FA1A S2_26_93 ( .A(\ab[26][93] ), .B(\CARRYB[25][93] ), .CI(\SUMB[25][94] ), 
        .CO(\CARRYB[26][93] ), .S(\SUMB[26][93] ) );
  FA1A S3_25_94 ( .A(\ab[25][94] ), .B(\CARRYB[24][94] ), .CI(\ab[24][95] ), 
        .CO(\CARRYB[25][94] ), .S(\SUMB[25][94] ) );
  FA1A S3_24_94 ( .A(\ab[24][94] ), .B(\CARRYB[23][94] ), .CI(\ab[23][95] ), 
        .CO(\CARRYB[24][94] ), .S(\SUMB[24][94] ) );
  FA1A S3_23_94 ( .A(\ab[23][94] ), .B(\CARRYB[22][94] ), .CI(\ab[22][95] ), 
        .CO(\CARRYB[23][94] ), .S(\SUMB[23][94] ) );
  FA1A S3_22_94 ( .A(\ab[22][94] ), .B(\CARRYB[21][94] ), .CI(\ab[21][95] ), 
        .CO(\CARRYB[22][94] ), .S(\SUMB[22][94] ) );
  FA1A S3_21_94 ( .A(\ab[21][94] ), .B(\CARRYB[20][94] ), .CI(\ab[20][95] ), 
        .CO(\CARRYB[21][94] ), .S(\SUMB[21][94] ) );
  FA1A S3_20_94 ( .A(\ab[20][94] ), .B(\CARRYB[19][94] ), .CI(\ab[19][95] ), 
        .CO(\CARRYB[20][94] ), .S(\SUMB[20][94] ) );
  FA1A S2_25_93 ( .A(\ab[25][93] ), .B(\CARRYB[24][93] ), .CI(\SUMB[24][94] ), 
        .CO(\CARRYB[25][93] ), .S(\SUMB[25][93] ) );
  FA1A S2_24_93 ( .A(\ab[24][93] ), .B(\CARRYB[23][93] ), .CI(\SUMB[23][94] ), 
        .CO(\CARRYB[24][93] ), .S(\SUMB[24][93] ) );
  FA1A S2_23_93 ( .A(\ab[23][93] ), .B(\CARRYB[22][93] ), .CI(\SUMB[22][94] ), 
        .CO(\CARRYB[23][93] ), .S(\SUMB[23][93] ) );
  FA1A S2_22_93 ( .A(\ab[22][93] ), .B(\CARRYB[21][93] ), .CI(\SUMB[21][94] ), 
        .CO(\CARRYB[22][93] ), .S(\SUMB[22][93] ) );
  FA1A S2_21_93 ( .A(\ab[21][93] ), .B(\CARRYB[20][93] ), .CI(\SUMB[20][94] ), 
        .CO(\CARRYB[21][93] ), .S(\SUMB[21][93] ) );
  FA1A S3_19_94 ( .A(\ab[19][94] ), .B(\CARRYB[18][94] ), .CI(\ab[18][95] ), 
        .CO(\CARRYB[19][94] ), .S(\SUMB[19][94] ) );
  FA1A S3_18_94 ( .A(\ab[18][94] ), .B(\CARRYB[17][94] ), .CI(\ab[17][95] ), 
        .CO(\CARRYB[18][94] ), .S(\SUMB[18][94] ) );
  FA1A S3_17_94 ( .A(\ab[17][94] ), .B(\CARRYB[16][94] ), .CI(\ab[16][95] ), 
        .CO(\CARRYB[17][94] ), .S(\SUMB[17][94] ) );
  FA1A S3_16_94 ( .A(\ab[16][94] ), .B(\CARRYB[15][94] ), .CI(\ab[15][95] ), 
        .CO(\CARRYB[16][94] ), .S(\SUMB[16][94] ) );
  FA1A S3_15_94 ( .A(\ab[15][94] ), .B(\CARRYB[14][94] ), .CI(\ab[14][95] ), 
        .CO(\CARRYB[15][94] ), .S(\SUMB[15][94] ) );
  FA1A S2_20_93 ( .A(\ab[20][93] ), .B(\CARRYB[19][93] ), .CI(\SUMB[19][94] ), 
        .CO(\CARRYB[20][93] ), .S(\SUMB[20][93] ) );
  FA1A S2_19_93 ( .A(\ab[19][93] ), .B(\CARRYB[18][93] ), .CI(\SUMB[18][94] ), 
        .CO(\CARRYB[19][93] ), .S(\SUMB[19][93] ) );
  FA1A S2_18_93 ( .A(\ab[18][93] ), .B(\CARRYB[17][93] ), .CI(\SUMB[17][94] ), 
        .CO(\CARRYB[18][93] ), .S(\SUMB[18][93] ) );
  FA1A S2_17_93 ( .A(\ab[17][93] ), .B(\CARRYB[16][93] ), .CI(\SUMB[16][94] ), 
        .CO(\CARRYB[17][93] ), .S(\SUMB[17][93] ) );
  FA1A S2_16_93 ( .A(\ab[16][93] ), .B(\CARRYB[15][93] ), .CI(\SUMB[15][94] ), 
        .CO(\CARRYB[16][93] ), .S(\SUMB[16][93] ) );
  FA1A S2_15_93 ( .A(\ab[15][93] ), .B(\CARRYB[14][93] ), .CI(\SUMB[14][94] ), 
        .CO(\CARRYB[15][93] ), .S(\SUMB[15][93] ) );
  FA1A S2_26_92 ( .A(\ab[26][92] ), .B(\CARRYB[25][92] ), .CI(\SUMB[25][93] ), 
        .CO(\CARRYB[26][92] ), .S(\SUMB[26][92] ) );
  FA1A S2_25_92 ( .A(\ab[25][92] ), .B(\CARRYB[24][92] ), .CI(\SUMB[24][93] ), 
        .CO(\CARRYB[25][92] ), .S(\SUMB[25][92] ) );
  FA1A S2_24_92 ( .A(\ab[24][92] ), .B(\CARRYB[23][92] ), .CI(\SUMB[23][93] ), 
        .CO(\CARRYB[24][92] ), .S(\SUMB[24][92] ) );
  FA1A S2_23_92 ( .A(\ab[23][92] ), .B(\CARRYB[22][92] ), .CI(\SUMB[22][93] ), 
        .CO(\CARRYB[23][92] ), .S(\SUMB[23][92] ) );
  FA1A S2_22_92 ( .A(\ab[22][92] ), .B(\CARRYB[21][92] ), .CI(\SUMB[21][93] ), 
        .CO(\CARRYB[22][92] ), .S(\SUMB[22][92] ) );
  FA1A S2_27_91 ( .A(\ab[27][91] ), .B(\CARRYB[26][91] ), .CI(\SUMB[26][92] ), 
        .CO(\CARRYB[27][91] ), .S(\SUMB[27][91] ) );
  FA1A S2_26_91 ( .A(\ab[26][91] ), .B(\CARRYB[25][91] ), .CI(\SUMB[25][92] ), 
        .CO(\CARRYB[26][91] ), .S(\SUMB[26][91] ) );
  FA1A S2_25_91 ( .A(\ab[25][91] ), .B(\CARRYB[24][91] ), .CI(\SUMB[24][92] ), 
        .CO(\CARRYB[25][91] ), .S(\SUMB[25][91] ) );
  FA1A S2_24_91 ( .A(\ab[24][91] ), .B(\CARRYB[23][91] ), .CI(\SUMB[23][92] ), 
        .CO(\CARRYB[24][91] ), .S(\SUMB[24][91] ) );
  FA1A S2_23_91 ( .A(\ab[23][91] ), .B(\CARRYB[22][91] ), .CI(\SUMB[22][92] ), 
        .CO(\CARRYB[23][91] ), .S(\SUMB[23][91] ) );
  FA1A S2_21_92 ( .A(\ab[21][92] ), .B(\CARRYB[20][92] ), .CI(\SUMB[20][93] ), 
        .CO(\CARRYB[21][92] ), .S(\SUMB[21][92] ) );
  FA1A S2_20_92 ( .A(\ab[20][92] ), .B(\CARRYB[19][92] ), .CI(\SUMB[19][93] ), 
        .CO(\CARRYB[20][92] ), .S(\SUMB[20][92] ) );
  FA1A S2_19_92 ( .A(\ab[19][92] ), .B(\CARRYB[18][92] ), .CI(\SUMB[18][93] ), 
        .CO(\CARRYB[19][92] ), .S(\SUMB[19][92] ) );
  FA1A S2_18_92 ( .A(\ab[18][92] ), .B(\CARRYB[17][92] ), .CI(\SUMB[17][93] ), 
        .CO(\CARRYB[18][92] ), .S(\SUMB[18][92] ) );
  FA1A S2_17_92 ( .A(\ab[17][92] ), .B(\CARRYB[16][92] ), .CI(\SUMB[16][93] ), 
        .CO(\CARRYB[17][92] ), .S(\SUMB[17][92] ) );
  FA1A S2_16_92 ( .A(\ab[16][92] ), .B(\CARRYB[15][92] ), .CI(\SUMB[15][93] ), 
        .CO(\CARRYB[16][92] ), .S(\SUMB[16][92] ) );
  FA1A S2_15_92 ( .A(\ab[15][92] ), .B(\CARRYB[14][92] ), .CI(\SUMB[14][93] ), 
        .CO(\CARRYB[15][92] ), .S(\SUMB[15][92] ) );
  FA1A S2_28_90 ( .A(\ab[28][90] ), .B(\CARRYB[27][90] ), .CI(\SUMB[27][91] ), 
        .CO(\CARRYB[28][90] ), .S(\SUMB[28][90] ) );
  FA1A S2_27_90 ( .A(\ab[27][90] ), .B(\CARRYB[26][90] ), .CI(\SUMB[26][91] ), 
        .CO(\CARRYB[27][90] ), .S(\SUMB[27][90] ) );
  FA1A S2_26_90 ( .A(\ab[26][90] ), .B(\CARRYB[25][90] ), .CI(\SUMB[25][91] ), 
        .CO(\CARRYB[26][90] ), .S(\SUMB[26][90] ) );
  FA1A S2_25_90 ( .A(\ab[25][90] ), .B(\CARRYB[24][90] ), .CI(\SUMB[24][91] ), 
        .CO(\CARRYB[25][90] ), .S(\SUMB[25][90] ) );
  FA1A S2_24_90 ( .A(\ab[24][90] ), .B(\CARRYB[23][90] ), .CI(\SUMB[23][91] ), 
        .CO(\CARRYB[24][90] ), .S(\SUMB[24][90] ) );
  FA1A S2_22_91 ( .A(\ab[22][91] ), .B(\CARRYB[21][91] ), .CI(\SUMB[21][92] ), 
        .CO(\CARRYB[22][91] ), .S(\SUMB[22][91] ) );
  FA1A S2_21_91 ( .A(\ab[21][91] ), .B(\CARRYB[20][91] ), .CI(\SUMB[20][92] ), 
        .CO(\CARRYB[21][91] ), .S(\SUMB[21][91] ) );
  FA1A S2_20_91 ( .A(\ab[20][91] ), .B(\CARRYB[19][91] ), .CI(\SUMB[19][92] ), 
        .CO(\CARRYB[20][91] ), .S(\SUMB[20][91] ) );
  FA1A S2_19_91 ( .A(\ab[19][91] ), .B(\CARRYB[18][91] ), .CI(\SUMB[18][92] ), 
        .CO(\CARRYB[19][91] ), .S(\SUMB[19][91] ) );
  FA1A S2_18_91 ( .A(\ab[18][91] ), .B(\CARRYB[17][91] ), .CI(\SUMB[17][92] ), 
        .CO(\CARRYB[18][91] ), .S(\SUMB[18][91] ) );
  FA1A S2_17_91 ( .A(\ab[17][91] ), .B(\CARRYB[16][91] ), .CI(\SUMB[16][92] ), 
        .CO(\CARRYB[17][91] ), .S(\SUMB[17][91] ) );
  FA1A S2_16_91 ( .A(\ab[16][91] ), .B(\CARRYB[15][91] ), .CI(\SUMB[15][92] ), 
        .CO(\CARRYB[16][91] ), .S(\SUMB[16][91] ) );
  FA1A S2_15_91 ( .A(\ab[15][91] ), .B(\CARRYB[14][91] ), .CI(\SUMB[14][92] ), 
        .CO(\CARRYB[15][91] ), .S(\SUMB[15][91] ) );
  FA1A S2_28_89 ( .A(\ab[28][89] ), .B(\CARRYB[27][89] ), .CI(\SUMB[27][90] ), 
        .CO(\CARRYB[28][89] ), .S(\SUMB[28][89] ) );
  FA1A S2_27_89 ( .A(\ab[27][89] ), .B(\CARRYB[26][89] ), .CI(\SUMB[26][90] ), 
        .CO(\CARRYB[27][89] ), .S(\SUMB[27][89] ) );
  FA1A S2_26_89 ( .A(\ab[26][89] ), .B(\CARRYB[25][89] ), .CI(\SUMB[25][90] ), 
        .CO(\CARRYB[26][89] ), .S(\SUMB[26][89] ) );
  FA1A S2_25_89 ( .A(\ab[25][89] ), .B(\CARRYB[24][89] ), .CI(\SUMB[24][90] ), 
        .CO(\CARRYB[25][89] ), .S(\SUMB[25][89] ) );
  FA1A S2_23_90 ( .A(\ab[23][90] ), .B(\CARRYB[22][90] ), .CI(\SUMB[22][91] ), 
        .CO(\CARRYB[23][90] ), .S(\SUMB[23][90] ) );
  FA1A S2_22_90 ( .A(\ab[22][90] ), .B(\CARRYB[21][90] ), .CI(\SUMB[21][91] ), 
        .CO(\CARRYB[22][90] ), .S(\SUMB[22][90] ) );
  FA1A S2_21_90 ( .A(\ab[21][90] ), .B(\CARRYB[20][90] ), .CI(\SUMB[20][91] ), 
        .CO(\CARRYB[21][90] ), .S(\SUMB[21][90] ) );
  FA1A S2_20_90 ( .A(\ab[20][90] ), .B(\CARRYB[19][90] ), .CI(\SUMB[19][91] ), 
        .CO(\CARRYB[20][90] ), .S(\SUMB[20][90] ) );
  FA1A S2_19_90 ( .A(\ab[19][90] ), .B(\CARRYB[18][90] ), .CI(\SUMB[18][91] ), 
        .CO(\CARRYB[19][90] ), .S(\SUMB[19][90] ) );
  FA1A S2_18_90 ( .A(\ab[18][90] ), .B(\CARRYB[17][90] ), .CI(\SUMB[17][91] ), 
        .CO(\CARRYB[18][90] ), .S(\SUMB[18][90] ) );
  FA1A S2_17_90 ( .A(\ab[17][90] ), .B(\CARRYB[16][90] ), .CI(\SUMB[16][91] ), 
        .CO(\CARRYB[17][90] ), .S(\SUMB[17][90] ) );
  FA1A S2_16_90 ( .A(\ab[16][90] ), .B(\CARRYB[15][90] ), .CI(\SUMB[15][91] ), 
        .CO(\CARRYB[16][90] ), .S(\SUMB[16][90] ) );
  FA1A S2_15_90 ( .A(\ab[15][90] ), .B(\CARRYB[14][90] ), .CI(\SUMB[14][91] ), 
        .CO(\CARRYB[15][90] ), .S(\SUMB[15][90] ) );
  FA1A S4_89 ( .A(\ab[29][89] ), .B(\CARRYB[28][89] ), .CI(\SUMB[28][90] ), 
        .CO(\CARRYB[29][89] ), .S(\SUMB[29][89] ) );
  FA1A S2_28_88 ( .A(\ab[28][88] ), .B(\CARRYB[27][88] ), .CI(\SUMB[27][89] ), 
        .CO(\CARRYB[28][88] ), .S(\SUMB[28][88] ) );
  FA1A S2_27_88 ( .A(\ab[27][88] ), .B(\CARRYB[26][88] ), .CI(\SUMB[26][89] ), 
        .CO(\CARRYB[27][88] ), .S(\SUMB[27][88] ) );
  FA1A S2_26_88 ( .A(\ab[26][88] ), .B(\CARRYB[25][88] ), .CI(\SUMB[25][89] ), 
        .CO(\CARRYB[26][88] ), .S(\SUMB[26][88] ) );
  FA1A S2_24_89 ( .A(\ab[24][89] ), .B(\CARRYB[23][89] ), .CI(\SUMB[23][90] ), 
        .CO(\CARRYB[24][89] ), .S(\SUMB[24][89] ) );
  FA1A S2_23_89 ( .A(\ab[23][89] ), .B(\CARRYB[22][89] ), .CI(\SUMB[22][90] ), 
        .CO(\CARRYB[23][89] ), .S(\SUMB[23][89] ) );
  FA1A S2_22_89 ( .A(\ab[22][89] ), .B(\CARRYB[21][89] ), .CI(\SUMB[21][90] ), 
        .CO(\CARRYB[22][89] ), .S(\SUMB[22][89] ) );
  FA1A S2_21_89 ( .A(\ab[21][89] ), .B(\CARRYB[20][89] ), .CI(\SUMB[20][90] ), 
        .CO(\CARRYB[21][89] ), .S(\SUMB[21][89] ) );
  FA1A S2_20_89 ( .A(\ab[20][89] ), .B(\CARRYB[19][89] ), .CI(\SUMB[19][90] ), 
        .CO(\CARRYB[20][89] ), .S(\SUMB[20][89] ) );
  FA1A S2_19_89 ( .A(\ab[19][89] ), .B(\CARRYB[18][89] ), .CI(\SUMB[18][90] ), 
        .CO(\CARRYB[19][89] ), .S(\SUMB[19][89] ) );
  FA1A S2_18_89 ( .A(\ab[18][89] ), .B(\CARRYB[17][89] ), .CI(\SUMB[17][90] ), 
        .CO(\CARRYB[18][89] ), .S(\SUMB[18][89] ) );
  FA1A S2_17_89 ( .A(\ab[17][89] ), .B(\CARRYB[16][89] ), .CI(\SUMB[16][90] ), 
        .CO(\CARRYB[17][89] ), .S(\SUMB[17][89] ) );
  FA1A S2_16_89 ( .A(\ab[16][89] ), .B(\CARRYB[15][89] ), .CI(\SUMB[15][90] ), 
        .CO(\CARRYB[16][89] ), .S(\SUMB[16][89] ) );
  FA1A S2_15_89 ( .A(\ab[15][89] ), .B(\CARRYB[14][89] ), .CI(\SUMB[14][90] ), 
        .CO(\CARRYB[15][89] ), .S(\SUMB[15][89] ) );
  FA1A S4_88 ( .A(\ab[29][88] ), .B(\CARRYB[28][88] ), .CI(\SUMB[28][89] ), 
        .CO(\CARRYB[29][88] ), .S(\SUMB[29][88] ) );
  FA1A S2_28_87 ( .A(\ab[28][87] ), .B(\CARRYB[27][87] ), .CI(\SUMB[27][88] ), 
        .CO(\CARRYB[28][87] ), .S(\SUMB[28][87] ) );
  FA1A S2_27_87 ( .A(\ab[27][87] ), .B(\CARRYB[26][87] ), .CI(\SUMB[26][88] ), 
        .CO(\CARRYB[27][87] ), .S(\SUMB[27][87] ) );
  FA1A S4_87 ( .A(\ab[29][87] ), .B(\CARRYB[28][87] ), .CI(\SUMB[28][88] ), 
        .CO(\CARRYB[29][87] ), .S(\SUMB[29][87] ) );
  FA1A S2_28_86 ( .A(\ab[28][86] ), .B(\CARRYB[27][86] ), .CI(\SUMB[27][87] ), 
        .CO(\CARRYB[28][86] ), .S(\SUMB[28][86] ) );
  FA1A S2_25_88 ( .A(\ab[25][88] ), .B(\CARRYB[24][88] ), .CI(\SUMB[24][89] ), 
        .CO(\CARRYB[25][88] ), .S(\SUMB[25][88] ) );
  FA1A S2_24_88 ( .A(\ab[24][88] ), .B(\CARRYB[23][88] ), .CI(\SUMB[23][89] ), 
        .CO(\CARRYB[24][88] ), .S(\SUMB[24][88] ) );
  FA1A S2_23_88 ( .A(\ab[23][88] ), .B(\CARRYB[22][88] ), .CI(\SUMB[22][89] ), 
        .CO(\CARRYB[23][88] ), .S(\SUMB[23][88] ) );
  FA1A S2_22_88 ( .A(\ab[22][88] ), .B(\CARRYB[21][88] ), .CI(\SUMB[21][89] ), 
        .CO(\CARRYB[22][88] ), .S(\SUMB[22][88] ) );
  FA1A S2_21_88 ( .A(\ab[21][88] ), .B(\CARRYB[20][88] ), .CI(\SUMB[20][89] ), 
        .CO(\CARRYB[21][88] ), .S(\SUMB[21][88] ) );
  FA1A S2_20_88 ( .A(\ab[20][88] ), .B(\CARRYB[19][88] ), .CI(\SUMB[19][89] ), 
        .CO(\CARRYB[20][88] ), .S(\SUMB[20][88] ) );
  FA1A S2_19_88 ( .A(\ab[19][88] ), .B(\CARRYB[18][88] ), .CI(\SUMB[18][89] ), 
        .CO(\CARRYB[19][88] ), .S(\SUMB[19][88] ) );
  FA1A S2_18_88 ( .A(\ab[18][88] ), .B(\CARRYB[17][88] ), .CI(\SUMB[17][89] ), 
        .CO(\CARRYB[18][88] ), .S(\SUMB[18][88] ) );
  FA1A S2_17_88 ( .A(\ab[17][88] ), .B(\CARRYB[16][88] ), .CI(\SUMB[16][89] ), 
        .CO(\CARRYB[17][88] ), .S(\SUMB[17][88] ) );
  FA1A S2_16_88 ( .A(\ab[16][88] ), .B(\CARRYB[15][88] ), .CI(\SUMB[15][89] ), 
        .CO(\CARRYB[16][88] ), .S(\SUMB[16][88] ) );
  FA1A S2_15_88 ( .A(\ab[15][88] ), .B(\CARRYB[14][88] ), .CI(\SUMB[14][89] ), 
        .CO(\CARRYB[15][88] ), .S(\SUMB[15][88] ) );
  FA1A S4_86 ( .A(\ab[29][86] ), .B(\CARRYB[28][86] ), .CI(\SUMB[28][87] ), 
        .CO(\CARRYB[29][86] ), .S(\SUMB[29][86] ) );
  FA1A S2_26_87 ( .A(\ab[26][87] ), .B(\CARRYB[25][87] ), .CI(\SUMB[25][88] ), 
        .CO(\CARRYB[26][87] ), .S(\SUMB[26][87] ) );
  FA1A S2_25_87 ( .A(\ab[25][87] ), .B(\CARRYB[24][87] ), .CI(\SUMB[24][88] ), 
        .CO(\CARRYB[25][87] ), .S(\SUMB[25][87] ) );
  FA1A S2_24_87 ( .A(\ab[24][87] ), .B(\CARRYB[23][87] ), .CI(\SUMB[23][88] ), 
        .CO(\CARRYB[24][87] ), .S(\SUMB[24][87] ) );
  FA1A S2_23_87 ( .A(\ab[23][87] ), .B(\CARRYB[22][87] ), .CI(\SUMB[22][88] ), 
        .CO(\CARRYB[23][87] ), .S(\SUMB[23][87] ) );
  FA1A S2_22_87 ( .A(\ab[22][87] ), .B(\CARRYB[21][87] ), .CI(\SUMB[21][88] ), 
        .CO(\CARRYB[22][87] ), .S(\SUMB[22][87] ) );
  FA1A S2_21_87 ( .A(\ab[21][87] ), .B(\CARRYB[20][87] ), .CI(\SUMB[20][88] ), 
        .CO(\CARRYB[21][87] ), .S(\SUMB[21][87] ) );
  FA1A S2_20_87 ( .A(\ab[20][87] ), .B(\CARRYB[19][87] ), .CI(\SUMB[19][88] ), 
        .CO(\CARRYB[20][87] ), .S(\SUMB[20][87] ) );
  FA1A S2_19_87 ( .A(\ab[19][87] ), .B(\CARRYB[18][87] ), .CI(\SUMB[18][88] ), 
        .CO(\CARRYB[19][87] ), .S(\SUMB[19][87] ) );
  FA1A S2_18_87 ( .A(\ab[18][87] ), .B(\CARRYB[17][87] ), .CI(\SUMB[17][88] ), 
        .CO(\CARRYB[18][87] ), .S(\SUMB[18][87] ) );
  FA1A S2_17_87 ( .A(\ab[17][87] ), .B(\CARRYB[16][87] ), .CI(\SUMB[16][88] ), 
        .CO(\CARRYB[17][87] ), .S(\SUMB[17][87] ) );
  FA1A S2_16_87 ( .A(\ab[16][87] ), .B(\CARRYB[15][87] ), .CI(\SUMB[15][88] ), 
        .CO(\CARRYB[16][87] ), .S(\SUMB[16][87] ) );
  FA1A S2_15_87 ( .A(\ab[15][87] ), .B(\CARRYB[14][87] ), .CI(\SUMB[14][88] ), 
        .CO(\CARRYB[15][87] ), .S(\SUMB[15][87] ) );
  FA1A S4_85 ( .A(\ab[29][85] ), .B(\CARRYB[28][85] ), .CI(\SUMB[28][86] ), 
        .CO(\CARRYB[29][85] ), .S(\SUMB[29][85] ) );
  FA1A S2_27_86 ( .A(\ab[27][86] ), .B(\CARRYB[26][86] ), .CI(\SUMB[26][87] ), 
        .CO(\CARRYB[27][86] ), .S(\SUMB[27][86] ) );
  FA1A S2_26_86 ( .A(\ab[26][86] ), .B(\CARRYB[25][86] ), .CI(\SUMB[25][87] ), 
        .CO(\CARRYB[26][86] ), .S(\SUMB[26][86] ) );
  FA1A S2_25_86 ( .A(\ab[25][86] ), .B(\CARRYB[24][86] ), .CI(\SUMB[24][87] ), 
        .CO(\CARRYB[25][86] ), .S(\SUMB[25][86] ) );
  FA1A S2_24_86 ( .A(\ab[24][86] ), .B(\CARRYB[23][86] ), .CI(\SUMB[23][87] ), 
        .CO(\CARRYB[24][86] ), .S(\SUMB[24][86] ) );
  FA1A S2_23_86 ( .A(\ab[23][86] ), .B(\CARRYB[22][86] ), .CI(\SUMB[22][87] ), 
        .CO(\CARRYB[23][86] ), .S(\SUMB[23][86] ) );
  FA1A S2_22_86 ( .A(\ab[22][86] ), .B(\CARRYB[21][86] ), .CI(\SUMB[21][87] ), 
        .CO(\CARRYB[22][86] ), .S(\SUMB[22][86] ) );
  FA1A S2_21_86 ( .A(\ab[21][86] ), .B(\CARRYB[20][86] ), .CI(\SUMB[20][87] ), 
        .CO(\CARRYB[21][86] ), .S(\SUMB[21][86] ) );
  FA1A S2_20_86 ( .A(\ab[20][86] ), .B(\CARRYB[19][86] ), .CI(\SUMB[19][87] ), 
        .CO(\CARRYB[20][86] ), .S(\SUMB[20][86] ) );
  FA1A S2_19_86 ( .A(\ab[19][86] ), .B(\CARRYB[18][86] ), .CI(\SUMB[18][87] ), 
        .CO(\CARRYB[19][86] ), .S(\SUMB[19][86] ) );
  FA1A S2_18_86 ( .A(\ab[18][86] ), .B(\CARRYB[17][86] ), .CI(\SUMB[17][87] ), 
        .CO(\CARRYB[18][86] ), .S(\SUMB[18][86] ) );
  FA1A S2_17_86 ( .A(\ab[17][86] ), .B(\CARRYB[16][86] ), .CI(\SUMB[16][87] ), 
        .CO(\CARRYB[17][86] ), .S(\SUMB[17][86] ) );
  FA1A S2_16_86 ( .A(\ab[16][86] ), .B(\CARRYB[15][86] ), .CI(\SUMB[15][87] ), 
        .CO(\CARRYB[16][86] ), .S(\SUMB[16][86] ) );
  FA1A S2_15_86 ( .A(\ab[15][86] ), .B(\CARRYB[14][86] ), .CI(\SUMB[14][87] ), 
        .CO(\CARRYB[15][86] ), .S(\SUMB[15][86] ) );
  FA1A S2_28_85 ( .A(\ab[28][85] ), .B(\CARRYB[27][85] ), .CI(\SUMB[27][86] ), 
        .CO(\CARRYB[28][85] ), .S(\SUMB[28][85] ) );
  FA1A S2_27_85 ( .A(\ab[27][85] ), .B(\CARRYB[26][85] ), .CI(\SUMB[26][86] ), 
        .CO(\CARRYB[27][85] ), .S(\SUMB[27][85] ) );
  FA1A S2_26_85 ( .A(\ab[26][85] ), .B(\CARRYB[25][85] ), .CI(\SUMB[25][86] ), 
        .CO(\CARRYB[26][85] ), .S(\SUMB[26][85] ) );
  FA1A S2_25_85 ( .A(\ab[25][85] ), .B(\CARRYB[24][85] ), .CI(\SUMB[24][86] ), 
        .CO(\CARRYB[25][85] ), .S(\SUMB[25][85] ) );
  FA1A S2_24_85 ( .A(\ab[24][85] ), .B(\CARRYB[23][85] ), .CI(\SUMB[23][86] ), 
        .CO(\CARRYB[24][85] ), .S(\SUMB[24][85] ) );
  FA1A S2_23_85 ( .A(\ab[23][85] ), .B(\CARRYB[22][85] ), .CI(\SUMB[22][86] ), 
        .CO(\CARRYB[23][85] ), .S(\SUMB[23][85] ) );
  FA1A S2_22_85 ( .A(\ab[22][85] ), .B(\CARRYB[21][85] ), .CI(\SUMB[21][86] ), 
        .CO(\CARRYB[22][85] ), .S(\SUMB[22][85] ) );
  FA1A S2_21_85 ( .A(\ab[21][85] ), .B(\CARRYB[20][85] ), .CI(\SUMB[20][86] ), 
        .CO(\CARRYB[21][85] ), .S(\SUMB[21][85] ) );
  FA1A S2_20_85 ( .A(\ab[20][85] ), .B(\CARRYB[19][85] ), .CI(\SUMB[19][86] ), 
        .CO(\CARRYB[20][85] ), .S(\SUMB[20][85] ) );
  FA1A S2_19_85 ( .A(\ab[19][85] ), .B(\CARRYB[18][85] ), .CI(\SUMB[18][86] ), 
        .CO(\CARRYB[19][85] ), .S(\SUMB[19][85] ) );
  FA1A S2_18_85 ( .A(\ab[18][85] ), .B(\CARRYB[17][85] ), .CI(\SUMB[17][86] ), 
        .CO(\CARRYB[18][85] ), .S(\SUMB[18][85] ) );
  FA1A S2_17_85 ( .A(\ab[17][85] ), .B(\CARRYB[16][85] ), .CI(\SUMB[16][86] ), 
        .CO(\CARRYB[17][85] ), .S(\SUMB[17][85] ) );
  FA1A S2_16_85 ( .A(\ab[16][85] ), .B(\CARRYB[15][85] ), .CI(\SUMB[15][86] ), 
        .CO(\CARRYB[16][85] ), .S(\SUMB[16][85] ) );
  FA1A S2_15_85 ( .A(\ab[15][85] ), .B(\CARRYB[14][85] ), .CI(\SUMB[14][86] ), 
        .CO(\CARRYB[15][85] ), .S(\SUMB[15][85] ) );
  FA1A S4_80 ( .A(\ab[29][80] ), .B(\CARRYB[28][80] ), .CI(\SUMB[28][81] ), 
        .CO(\CARRYB[29][80] ), .S(\SUMB[29][80] ) );
  FA1A S4_81 ( .A(\ab[29][81] ), .B(\CARRYB[28][81] ), .CI(\SUMB[28][82] ), 
        .CO(\CARRYB[29][81] ), .S(\SUMB[29][81] ) );
  FA1A S2_28_81 ( .A(\ab[28][81] ), .B(\CARRYB[27][81] ), .CI(\SUMB[27][82] ), 
        .CO(\CARRYB[28][81] ), .S(\SUMB[28][81] ) );
  FA1A S2_27_81 ( .A(\ab[27][81] ), .B(\CARRYB[26][81] ), .CI(\SUMB[26][82] ), 
        .CO(\CARRYB[27][81] ), .S(\SUMB[27][81] ) );
  FA1A S2_26_81 ( .A(\ab[26][81] ), .B(\CARRYB[25][81] ), .CI(\SUMB[25][82] ), 
        .CO(\CARRYB[26][81] ), .S(\SUMB[26][81] ) );
  FA1A S2_25_81 ( .A(\ab[25][81] ), .B(\CARRYB[24][81] ), .CI(\SUMB[24][82] ), 
        .CO(\CARRYB[25][81] ), .S(\SUMB[25][81] ) );
  FA1A S2_24_81 ( .A(\ab[24][81] ), .B(\CARRYB[23][81] ), .CI(\SUMB[23][82] ), 
        .CO(\CARRYB[24][81] ), .S(\SUMB[24][81] ) );
  FA1A S2_23_81 ( .A(\ab[23][81] ), .B(\CARRYB[22][81] ), .CI(\SUMB[22][82] ), 
        .CO(\CARRYB[23][81] ), .S(\SUMB[23][81] ) );
  FA1A S2_22_81 ( .A(\ab[22][81] ), .B(\CARRYB[21][81] ), .CI(\SUMB[21][82] ), 
        .CO(\CARRYB[22][81] ), .S(\SUMB[22][81] ) );
  FA1A S2_21_81 ( .A(\ab[21][81] ), .B(\CARRYB[20][81] ), .CI(\SUMB[20][82] ), 
        .CO(\CARRYB[21][81] ), .S(\SUMB[21][81] ) );
  FA1A S2_20_81 ( .A(\ab[20][81] ), .B(\CARRYB[19][81] ), .CI(\SUMB[19][82] ), 
        .CO(\CARRYB[20][81] ), .S(\SUMB[20][81] ) );
  FA1A S2_19_81 ( .A(\ab[19][81] ), .B(\CARRYB[18][81] ), .CI(\SUMB[18][82] ), 
        .CO(\CARRYB[19][81] ), .S(\SUMB[19][81] ) );
  FA1A S2_18_81 ( .A(\ab[18][81] ), .B(\CARRYB[17][81] ), .CI(\SUMB[17][82] ), 
        .CO(\CARRYB[18][81] ), .S(\SUMB[18][81] ) );
  FA1A S2_17_81 ( .A(\ab[17][81] ), .B(\CARRYB[16][81] ), .CI(\SUMB[16][82] ), 
        .CO(\CARRYB[17][81] ), .S(\SUMB[17][81] ) );
  FA1A S2_16_81 ( .A(\ab[16][81] ), .B(\CARRYB[15][81] ), .CI(\SUMB[15][82] ), 
        .CO(\CARRYB[16][81] ), .S(\SUMB[16][81] ) );
  FA1A S2_15_81 ( .A(\ab[15][81] ), .B(\CARRYB[14][81] ), .CI(\SUMB[14][82] ), 
        .CO(\CARRYB[15][81] ), .S(\SUMB[15][81] ) );
  FA1A S2_28_80 ( .A(\ab[28][80] ), .B(\CARRYB[27][80] ), .CI(\SUMB[27][81] ), 
        .CO(\CARRYB[28][80] ), .S(\SUMB[28][80] ) );
  FA1A S4_82 ( .A(\ab[29][82] ), .B(\CARRYB[28][82] ), .CI(\SUMB[28][83] ), 
        .CO(\CARRYB[29][82] ), .S(\SUMB[29][82] ) );
  FA1A S2_27_80 ( .A(\ab[27][80] ), .B(\CARRYB[26][80] ), .CI(\SUMB[26][81] ), 
        .CO(\CARRYB[27][80] ), .S(\SUMB[27][80] ) );
  FA1A S2_28_82 ( .A(\ab[28][82] ), .B(\CARRYB[27][82] ), .CI(\SUMB[27][83] ), 
        .CO(\CARRYB[28][82] ), .S(\SUMB[28][82] ) );
  FA1A S4_83 ( .A(\ab[29][83] ), .B(\CARRYB[28][83] ), .CI(\SUMB[28][84] ), 
        .CO(\CARRYB[29][83] ), .S(\SUMB[29][83] ) );
  FA1A S2_26_80 ( .A(\ab[26][80] ), .B(\CARRYB[25][80] ), .CI(\SUMB[25][81] ), 
        .CO(\CARRYB[26][80] ), .S(\SUMB[26][80] ) );
  FA1A S2_27_82 ( .A(\ab[27][82] ), .B(\CARRYB[26][82] ), .CI(\SUMB[26][83] ), 
        .CO(\CARRYB[27][82] ), .S(\SUMB[27][82] ) );
  FA1A S2_28_84 ( .A(\ab[28][84] ), .B(\CARRYB[27][84] ), .CI(\SUMB[27][85] ), 
        .CO(\CARRYB[28][84] ), .S(\SUMB[28][84] ) );
  FA1A S2_28_83 ( .A(\ab[28][83] ), .B(\CARRYB[27][83] ), .CI(\SUMB[27][84] ), 
        .CO(\CARRYB[28][83] ), .S(\SUMB[28][83] ) );
  FA1A S2_25_80 ( .A(\ab[25][80] ), .B(\CARRYB[24][80] ), .CI(\SUMB[24][81] ), 
        .CO(\CARRYB[25][80] ), .S(\SUMB[25][80] ) );
  FA1A S2_26_82 ( .A(\ab[26][82] ), .B(\CARRYB[25][82] ), .CI(\SUMB[25][83] ), 
        .CO(\CARRYB[26][82] ), .S(\SUMB[26][82] ) );
  FA1A S2_27_84 ( .A(\ab[27][84] ), .B(\CARRYB[26][84] ), .CI(\SUMB[26][85] ), 
        .CO(\CARRYB[27][84] ), .S(\SUMB[27][84] ) );
  FA1A S2_27_83 ( .A(\ab[27][83] ), .B(\CARRYB[26][83] ), .CI(\SUMB[26][84] ), 
        .CO(\CARRYB[27][83] ), .S(\SUMB[27][83] ) );
  FA1A S2_25_82 ( .A(\ab[25][82] ), .B(\CARRYB[24][82] ), .CI(\SUMB[24][83] ), 
        .CO(\CARRYB[25][82] ), .S(\SUMB[25][82] ) );
  FA1A S2_26_84 ( .A(\ab[26][84] ), .B(\CARRYB[25][84] ), .CI(\SUMB[25][85] ), 
        .CO(\CARRYB[26][84] ), .S(\SUMB[26][84] ) );
  FA1A S2_26_83 ( .A(\ab[26][83] ), .B(\CARRYB[25][83] ), .CI(\SUMB[25][84] ), 
        .CO(\CARRYB[26][83] ), .S(\SUMB[26][83] ) );
  FA1A S2_24_80 ( .A(\ab[24][80] ), .B(\CARRYB[23][80] ), .CI(\SUMB[23][81] ), 
        .CO(\CARRYB[24][80] ), .S(\SUMB[24][80] ) );
  FA1A S2_24_82 ( .A(\ab[24][82] ), .B(\CARRYB[23][82] ), .CI(\SUMB[23][83] ), 
        .CO(\CARRYB[24][82] ), .S(\SUMB[24][82] ) );
  FA1A S2_25_84 ( .A(\ab[25][84] ), .B(\CARRYB[24][84] ), .CI(\SUMB[24][85] ), 
        .CO(\CARRYB[25][84] ), .S(\SUMB[25][84] ) );
  FA1A S2_25_83 ( .A(\ab[25][83] ), .B(\CARRYB[24][83] ), .CI(\SUMB[24][84] ), 
        .CO(\CARRYB[25][83] ), .S(\SUMB[25][83] ) );
  FA1A S2_23_80 ( .A(\ab[23][80] ), .B(\CARRYB[22][80] ), .CI(\SUMB[22][81] ), 
        .CO(\CARRYB[23][80] ), .S(\SUMB[23][80] ) );
  FA1A S2_23_82 ( .A(\ab[23][82] ), .B(\CARRYB[22][82] ), .CI(\SUMB[22][83] ), 
        .CO(\CARRYB[23][82] ), .S(\SUMB[23][82] ) );
  FA1A S2_24_84 ( .A(\ab[24][84] ), .B(\CARRYB[23][84] ), .CI(\SUMB[23][85] ), 
        .CO(\CARRYB[24][84] ), .S(\SUMB[24][84] ) );
  FA1A S2_24_83 ( .A(\ab[24][83] ), .B(\CARRYB[23][83] ), .CI(\SUMB[23][84] ), 
        .CO(\CARRYB[24][83] ), .S(\SUMB[24][83] ) );
  FA1A S2_22_82 ( .A(\ab[22][82] ), .B(\CARRYB[21][82] ), .CI(\SUMB[21][83] ), 
        .CO(\CARRYB[22][82] ), .S(\SUMB[22][82] ) );
  FA1A S2_22_80 ( .A(\ab[22][80] ), .B(\CARRYB[21][80] ), .CI(\SUMB[21][81] ), 
        .CO(\CARRYB[22][80] ), .S(\SUMB[22][80] ) );
  FA1A S2_23_84 ( .A(\ab[23][84] ), .B(\CARRYB[22][84] ), .CI(\SUMB[22][85] ), 
        .CO(\CARRYB[23][84] ), .S(\SUMB[23][84] ) );
  FA1A S2_23_83 ( .A(\ab[23][83] ), .B(\CARRYB[22][83] ), .CI(\SUMB[22][84] ), 
        .CO(\CARRYB[23][83] ), .S(\SUMB[23][83] ) );
  FA1A S2_21_82 ( .A(\ab[21][82] ), .B(\CARRYB[20][82] ), .CI(\SUMB[20][83] ), 
        .CO(\CARRYB[21][82] ), .S(\SUMB[21][82] ) );
  FA1A S2_21_80 ( .A(\ab[21][80] ), .B(\CARRYB[20][80] ), .CI(\SUMB[20][81] ), 
        .CO(\CARRYB[21][80] ), .S(\SUMB[21][80] ) );
  FA1A S2_22_84 ( .A(\ab[22][84] ), .B(\CARRYB[21][84] ), .CI(\SUMB[21][85] ), 
        .CO(\CARRYB[22][84] ), .S(\SUMB[22][84] ) );
  FA1A S2_22_83 ( .A(\ab[22][83] ), .B(\CARRYB[21][83] ), .CI(\SUMB[21][84] ), 
        .CO(\CARRYB[22][83] ), .S(\SUMB[22][83] ) );
  FA1A S2_20_82 ( .A(\ab[20][82] ), .B(\CARRYB[19][82] ), .CI(\SUMB[19][83] ), 
        .CO(\CARRYB[20][82] ), .S(\SUMB[20][82] ) );
  FA1A S2_20_80 ( .A(\ab[20][80] ), .B(\CARRYB[19][80] ), .CI(\SUMB[19][81] ), 
        .CO(\CARRYB[20][80] ), .S(\SUMB[20][80] ) );
  FA1A S2_21_84 ( .A(\ab[21][84] ), .B(\CARRYB[20][84] ), .CI(\SUMB[20][85] ), 
        .CO(\CARRYB[21][84] ), .S(\SUMB[21][84] ) );
  FA1A S2_21_83 ( .A(\ab[21][83] ), .B(\CARRYB[20][83] ), .CI(\SUMB[20][84] ), 
        .CO(\CARRYB[21][83] ), .S(\SUMB[21][83] ) );
  FA1A S2_19_82 ( .A(\ab[19][82] ), .B(\CARRYB[18][82] ), .CI(\SUMB[18][83] ), 
        .CO(\CARRYB[19][82] ), .S(\SUMB[19][82] ) );
  FA1A S2_20_84 ( .A(\ab[20][84] ), .B(\CARRYB[19][84] ), .CI(\SUMB[19][85] ), 
        .CO(\CARRYB[20][84] ), .S(\SUMB[20][84] ) );
  FA1A S2_20_83 ( .A(\ab[20][83] ), .B(\CARRYB[19][83] ), .CI(\SUMB[19][84] ), 
        .CO(\CARRYB[20][83] ), .S(\SUMB[20][83] ) );
  FA1A S2_18_82 ( .A(\ab[18][82] ), .B(\CARRYB[17][82] ), .CI(\SUMB[17][83] ), 
        .CO(\CARRYB[18][82] ), .S(\SUMB[18][82] ) );
  FA1A S2_19_84 ( .A(\ab[19][84] ), .B(\CARRYB[18][84] ), .CI(\SUMB[18][85] ), 
        .CO(\CARRYB[19][84] ), .S(\SUMB[19][84] ) );
  FA1A S2_19_83 ( .A(\ab[19][83] ), .B(\CARRYB[18][83] ), .CI(\SUMB[18][84] ), 
        .CO(\CARRYB[19][83] ), .S(\SUMB[19][83] ) );
  FA1A S2_18_84 ( .A(\ab[18][84] ), .B(\CARRYB[17][84] ), .CI(\SUMB[17][85] ), 
        .CO(\CARRYB[18][84] ), .S(\SUMB[18][84] ) );
  FA1A S2_18_83 ( .A(\ab[18][83] ), .B(\CARRYB[17][83] ), .CI(\SUMB[17][84] ), 
        .CO(\CARRYB[18][83] ), .S(\SUMB[18][83] ) );
  FA1A S2_17_84 ( .A(\ab[17][84] ), .B(\CARRYB[16][84] ), .CI(\SUMB[16][85] ), 
        .CO(\CARRYB[17][84] ), .S(\SUMB[17][84] ) );
  FA1A S2_17_83 ( .A(\ab[17][83] ), .B(\CARRYB[16][83] ), .CI(\SUMB[16][84] ), 
        .CO(\CARRYB[17][83] ), .S(\SUMB[17][83] ) );
  FA1A S2_16_84 ( .A(\ab[16][84] ), .B(\CARRYB[15][84] ), .CI(\SUMB[15][85] ), 
        .CO(\CARRYB[16][84] ), .S(\SUMB[16][84] ) );
  FA1A S2_19_80 ( .A(\ab[19][80] ), .B(\CARRYB[18][80] ), .CI(\SUMB[18][81] ), 
        .CO(\CARRYB[19][80] ), .S(\SUMB[19][80] ) );
  FA1A S2_18_80 ( .A(\ab[18][80] ), .B(\CARRYB[17][80] ), .CI(\SUMB[17][81] ), 
        .CO(\CARRYB[18][80] ), .S(\SUMB[18][80] ) );
  FA1A S2_17_82 ( .A(\ab[17][82] ), .B(\CARRYB[16][82] ), .CI(\SUMB[16][83] ), 
        .CO(\CARRYB[17][82] ), .S(\SUMB[17][82] ) );
  FA1A S2_17_80 ( .A(\ab[17][80] ), .B(\CARRYB[16][80] ), .CI(\SUMB[16][81] ), 
        .CO(\CARRYB[17][80] ), .S(\SUMB[17][80] ) );
  FA1A S2_16_83 ( .A(\ab[16][83] ), .B(\CARRYB[15][83] ), .CI(\SUMB[15][84] ), 
        .CO(\CARRYB[16][83] ), .S(\SUMB[16][83] ) );
  FA1A S2_16_82 ( .A(\ab[16][82] ), .B(\CARRYB[15][82] ), .CI(\SUMB[15][83] ), 
        .CO(\CARRYB[16][82] ), .S(\SUMB[16][82] ) );
  FA1A S2_15_84 ( .A(\ab[15][84] ), .B(\CARRYB[14][84] ), .CI(\SUMB[14][85] ), 
        .CO(\CARRYB[15][84] ), .S(\SUMB[15][84] ) );
  FA1A S2_15_83 ( .A(\ab[15][83] ), .B(\CARRYB[14][83] ), .CI(\SUMB[14][84] ), 
        .CO(\CARRYB[15][83] ), .S(\SUMB[15][83] ) );
  FA1A S2_15_82 ( .A(\ab[15][82] ), .B(\CARRYB[14][82] ), .CI(\SUMB[14][83] ), 
        .CO(\CARRYB[15][82] ), .S(\SUMB[15][82] ) );
  FA1A S2_16_80 ( .A(\ab[16][80] ), .B(\CARRYB[15][80] ), .CI(\SUMB[15][81] ), 
        .CO(\CARRYB[16][80] ), .S(\SUMB[16][80] ) );
  FA1A S2_15_80 ( .A(\ab[15][80] ), .B(\CARRYB[14][80] ), .CI(\SUMB[14][81] ), 
        .CO(\CARRYB[15][80] ), .S(\SUMB[15][80] ) );
  FA1A S4_84 ( .A(\ab[29][84] ), .B(\CARRYB[28][84] ), .CI(\SUMB[28][85] ), 
        .CO(\CARRYB[29][84] ), .S(\SUMB[29][84] ) );
  FA1A S4_73 ( .A(\ab[29][73] ), .B(\CARRYB[28][73] ), .CI(\SUMB[28][74] ), 
        .CO(\CARRYB[29][73] ), .S(\SUMB[29][73] ) );
  FA1A S4_78 ( .A(\ab[29][78] ), .B(\CARRYB[28][78] ), .CI(\SUMB[28][79] ), 
        .CO(\CARRYB[29][78] ), .S(\SUMB[29][78] ) );
  FA1A S4_77 ( .A(\ab[29][77] ), .B(\CARRYB[28][77] ), .CI(\SUMB[28][78] ), 
        .CO(\CARRYB[29][77] ), .S(\SUMB[29][77] ) );
  FA1A S2_28_73 ( .A(\ab[28][73] ), .B(\CARRYB[27][73] ), .CI(\SUMB[27][74] ), 
        .CO(\CARRYB[28][73] ), .S(\SUMB[28][73] ) );
  FA1A S2_28_79 ( .A(\ab[28][79] ), .B(\CARRYB[27][79] ), .CI(\SUMB[27][80] ), 
        .CO(\CARRYB[28][79] ), .S(\SUMB[28][79] ) );
  FA1A S2_28_78 ( .A(\ab[28][78] ), .B(\CARRYB[27][78] ), .CI(\SUMB[27][79] ), 
        .CO(\CARRYB[28][78] ), .S(\SUMB[28][78] ) );
  FA1A S2_28_77 ( .A(\ab[28][77] ), .B(\CARRYB[27][77] ), .CI(\SUMB[27][78] ), 
        .CO(\CARRYB[28][77] ), .S(\SUMB[28][77] ) );
  FA1A S4_75 ( .A(\ab[29][75] ), .B(\CARRYB[28][75] ), .CI(\SUMB[28][76] ), 
        .CO(\CARRYB[29][75] ), .S(\SUMB[29][75] ) );
  FA1A S4_71 ( .A(\ab[29][71] ), .B(\CARRYB[28][71] ), .CI(\SUMB[28][72] ), 
        .CO(\CARRYB[29][71] ), .S(\SUMB[29][71] ) );
  FA1A S2_27_79 ( .A(\ab[27][79] ), .B(\CARRYB[26][79] ), .CI(\SUMB[26][80] ), 
        .CO(\CARRYB[27][79] ), .S(\SUMB[27][79] ) );
  FA1A S2_27_78 ( .A(\ab[27][78] ), .B(\CARRYB[26][78] ), .CI(\SUMB[26][79] ), 
        .CO(\CARRYB[27][78] ), .S(\SUMB[27][78] ) );
  FA1A S2_28_76 ( .A(\ab[28][76] ), .B(\CARRYB[27][76] ), .CI(\SUMB[27][77] ), 
        .CO(\CARRYB[28][76] ), .S(\SUMB[28][76] ) );
  FA1A S2_28_75 ( .A(\ab[28][75] ), .B(\CARRYB[27][75] ), .CI(\SUMB[27][76] ), 
        .CO(\CARRYB[28][75] ), .S(\SUMB[28][75] ) );
  FA1A S2_28_74 ( .A(\ab[28][74] ), .B(\CARRYB[27][74] ), .CI(\SUMB[27][75] ), 
        .CO(\CARRYB[28][74] ), .S(\SUMB[28][74] ) );
  FA1A S2_28_72 ( .A(\ab[28][72] ), .B(\CARRYB[27][72] ), .CI(\SUMB[27][73] ), 
        .CO(\CARRYB[28][72] ), .S(\SUMB[28][72] ) );
  FA1A S4_69 ( .A(\ab[29][69] ), .B(\CARRYB[28][69] ), .CI(\SUMB[28][70] ), 
        .CO(\CARRYB[29][69] ), .S(\SUMB[29][69] ) );
  FA1A S2_26_79 ( .A(\ab[26][79] ), .B(\CARRYB[25][79] ), .CI(\SUMB[25][80] ), 
        .CO(\CARRYB[26][79] ), .S(\SUMB[26][79] ) );
  FA1A S2_27_77 ( .A(\ab[27][77] ), .B(\CARRYB[26][77] ), .CI(\SUMB[26][78] ), 
        .CO(\CARRYB[27][77] ), .S(\SUMB[27][77] ) );
  FA1A S2_27_76 ( .A(\ab[27][76] ), .B(\CARRYB[26][76] ), .CI(\SUMB[26][77] ), 
        .CO(\CARRYB[27][76] ), .S(\SUMB[27][76] ) );
  FA1A S2_27_75 ( .A(\ab[27][75] ), .B(\CARRYB[26][75] ), .CI(\SUMB[26][76] ), 
        .CO(\CARRYB[27][75] ), .S(\SUMB[27][75] ) );
  FA1A S2_27_74 ( .A(\ab[27][74] ), .B(\CARRYB[26][74] ), .CI(\SUMB[26][75] ), 
        .CO(\CARRYB[27][74] ), .S(\SUMB[27][74] ) );
  FA1A S2_27_73 ( .A(\ab[27][73] ), .B(\CARRYB[26][73] ), .CI(\SUMB[26][74] ), 
        .CO(\CARRYB[27][73] ), .S(\SUMB[27][73] ) );
  FA1A S2_28_69 ( .A(\ab[28][69] ), .B(\CARRYB[27][69] ), .CI(\SUMB[27][70] ), 
        .CO(\CARRYB[28][69] ), .S(\SUMB[28][69] ) );
  FA1A S2_26_78 ( .A(\ab[26][78] ), .B(\CARRYB[25][78] ), .CI(\SUMB[25][79] ), 
        .CO(\CARRYB[26][78] ), .S(\SUMB[26][78] ) );
  FA1A S2_26_77 ( .A(\ab[26][77] ), .B(\CARRYB[25][77] ), .CI(\SUMB[25][78] ), 
        .CO(\CARRYB[26][77] ), .S(\SUMB[26][77] ) );
  FA1A S2_26_76 ( .A(\ab[26][76] ), .B(\CARRYB[25][76] ), .CI(\SUMB[25][77] ), 
        .CO(\CARRYB[26][76] ), .S(\SUMB[26][76] ) );
  FA1A S2_26_75 ( .A(\ab[26][75] ), .B(\CARRYB[25][75] ), .CI(\SUMB[25][76] ), 
        .CO(\CARRYB[26][75] ), .S(\SUMB[26][75] ) );
  FA1A S2_26_74 ( .A(\ab[26][74] ), .B(\CARRYB[25][74] ), .CI(\SUMB[25][75] ), 
        .CO(\CARRYB[26][74] ), .S(\SUMB[26][74] ) );
  FA1A S2_25_79 ( .A(\ab[25][79] ), .B(\CARRYB[24][79] ), .CI(\SUMB[24][80] ), 
        .CO(\CARRYB[25][79] ), .S(\SUMB[25][79] ) );
  FA1A S2_25_78 ( .A(\ab[25][78] ), .B(\CARRYB[24][78] ), .CI(\SUMB[24][79] ), 
        .CO(\CARRYB[25][78] ), .S(\SUMB[25][78] ) );
  FA1A S2_25_77 ( .A(\ab[25][77] ), .B(\CARRYB[24][77] ), .CI(\SUMB[24][78] ), 
        .CO(\CARRYB[25][77] ), .S(\SUMB[25][77] ) );
  FA1A S2_25_76 ( .A(\ab[25][76] ), .B(\CARRYB[24][76] ), .CI(\SUMB[24][77] ), 
        .CO(\CARRYB[25][76] ), .S(\SUMB[25][76] ) );
  FA1A S2_25_75 ( .A(\ab[25][75] ), .B(\CARRYB[24][75] ), .CI(\SUMB[24][76] ), 
        .CO(\CARRYB[25][75] ), .S(\SUMB[25][75] ) );
  FA1A S2_24_79 ( .A(\ab[24][79] ), .B(\CARRYB[23][79] ), .CI(\SUMB[23][80] ), 
        .CO(\CARRYB[24][79] ), .S(\SUMB[24][79] ) );
  FA1A S2_24_78 ( .A(\ab[24][78] ), .B(\CARRYB[23][78] ), .CI(\SUMB[23][79] ), 
        .CO(\CARRYB[24][78] ), .S(\SUMB[24][78] ) );
  FA1A S2_24_77 ( .A(\ab[24][77] ), .B(\CARRYB[23][77] ), .CI(\SUMB[23][78] ), 
        .CO(\CARRYB[24][77] ), .S(\SUMB[24][77] ) );
  FA1A S2_24_76 ( .A(\ab[24][76] ), .B(\CARRYB[23][76] ), .CI(\SUMB[23][77] ), 
        .CO(\CARRYB[24][76] ), .S(\SUMB[24][76] ) );
  FA1A S4_57 ( .A(\ab[29][57] ), .B(\CARRYB[28][57] ), .CI(\SUMB[28][58] ), 
        .CO(\CARRYB[29][57] ), .S(\SUMB[29][57] ) );
  FA1A S2_23_79 ( .A(\ab[23][79] ), .B(\CARRYB[22][79] ), .CI(\SUMB[22][80] ), 
        .CO(\CARRYB[23][79] ), .S(\SUMB[23][79] ) );
  FA1A S2_23_78 ( .A(\ab[23][78] ), .B(\CARRYB[22][78] ), .CI(\SUMB[22][79] ), 
        .CO(\CARRYB[23][78] ), .S(\SUMB[23][78] ) );
  FA1A S2_23_77 ( .A(\ab[23][77] ), .B(\CARRYB[22][77] ), .CI(\SUMB[22][78] ), 
        .CO(\CARRYB[23][77] ), .S(\SUMB[23][77] ) );
  FA1A S2_28_57 ( .A(\ab[28][57] ), .B(\CARRYB[27][57] ), .CI(\SUMB[27][58] ), 
        .CO(\CARRYB[28][57] ), .S(\SUMB[28][57] ) );
  FA1A S2_22_79 ( .A(\ab[22][79] ), .B(\CARRYB[21][79] ), .CI(\SUMB[21][80] ), 
        .CO(\CARRYB[22][79] ), .S(\SUMB[22][79] ) );
  FA1A S2_22_78 ( .A(\ab[22][78] ), .B(\CARRYB[21][78] ), .CI(\SUMB[21][79] ), 
        .CO(\CARRYB[22][78] ), .S(\SUMB[22][78] ) );
  FA1A S2_28_71 ( .A(\ab[28][71] ), .B(\CARRYB[27][71] ), .CI(\SUMB[27][72] ), 
        .CO(\CARRYB[28][71] ), .S(\SUMB[28][71] ) );
  FA1A S2_28_70 ( .A(\ab[28][70] ), .B(\CARRYB[27][70] ), .CI(\SUMB[27][71] ), 
        .CO(\CARRYB[28][70] ), .S(\SUMB[28][70] ) );
  FA1A S2_21_79 ( .A(\ab[21][79] ), .B(\CARRYB[20][79] ), .CI(\SUMB[20][80] ), 
        .CO(\CARRYB[21][79] ), .S(\SUMB[21][79] ) );
  FA1A S2_27_72 ( .A(\ab[27][72] ), .B(\CARRYB[26][72] ), .CI(\SUMB[26][73] ), 
        .CO(\CARRYB[27][72] ), .S(\SUMB[27][72] ) );
  FA1A S2_27_71 ( .A(\ab[27][71] ), .B(\CARRYB[26][71] ), .CI(\SUMB[26][72] ), 
        .CO(\CARRYB[27][71] ), .S(\SUMB[27][71] ) );
  FA1A S2_27_70 ( .A(\ab[27][70] ), .B(\CARRYB[26][70] ), .CI(\SUMB[26][71] ), 
        .CO(\CARRYB[27][70] ), .S(\SUMB[27][70] ) );
  FA1A S2_27_57 ( .A(\ab[27][57] ), .B(\CARRYB[26][57] ), .CI(\SUMB[26][58] ), 
        .CO(\CARRYB[27][57] ), .S(\SUMB[27][57] ) );
  FA1A S2_26_73 ( .A(\ab[26][73] ), .B(\CARRYB[25][73] ), .CI(\SUMB[25][74] ), 
        .CO(\CARRYB[26][73] ), .S(\SUMB[26][73] ) );
  FA1A S2_26_72 ( .A(\ab[26][72] ), .B(\CARRYB[25][72] ), .CI(\SUMB[25][73] ), 
        .CO(\CARRYB[26][72] ), .S(\SUMB[26][72] ) );
  FA1A S2_26_71 ( .A(\ab[26][71] ), .B(\CARRYB[25][71] ), .CI(\SUMB[25][72] ), 
        .CO(\CARRYB[26][71] ), .S(\SUMB[26][71] ) );
  FA1A S2_25_74 ( .A(\ab[25][74] ), .B(\CARRYB[24][74] ), .CI(\SUMB[24][75] ), 
        .CO(\CARRYB[25][74] ), .S(\SUMB[25][74] ) );
  FA1A S2_25_73 ( .A(\ab[25][73] ), .B(\CARRYB[24][73] ), .CI(\SUMB[24][74] ), 
        .CO(\CARRYB[25][73] ), .S(\SUMB[25][73] ) );
  FA1A S2_25_72 ( .A(\ab[25][72] ), .B(\CARRYB[24][72] ), .CI(\SUMB[24][73] ), 
        .CO(\CARRYB[25][72] ), .S(\SUMB[25][72] ) );
  FA1A S2_27_69 ( .A(\ab[27][69] ), .B(\CARRYB[26][69] ), .CI(\SUMB[26][70] ), 
        .CO(\CARRYB[27][69] ), .S(\SUMB[27][69] ) );
  FA1A S2_26_57 ( .A(\ab[26][57] ), .B(\CARRYB[25][57] ), .CI(\SUMB[25][58] ), 
        .CO(\CARRYB[26][57] ), .S(\SUMB[26][57] ) );
  FA1A S2_24_75 ( .A(\ab[24][75] ), .B(\CARRYB[23][75] ), .CI(\SUMB[23][76] ), 
        .CO(\CARRYB[24][75] ), .S(\SUMB[24][75] ) );
  FA1A S2_24_74 ( .A(\ab[24][74] ), .B(\CARRYB[23][74] ), .CI(\SUMB[23][75] ), 
        .CO(\CARRYB[24][74] ), .S(\SUMB[24][74] ) );
  FA1A S2_24_73 ( .A(\ab[24][73] ), .B(\CARRYB[23][73] ), .CI(\SUMB[23][74] ), 
        .CO(\CARRYB[24][73] ), .S(\SUMB[24][73] ) );
  FA1A S2_26_69 ( .A(\ab[26][69] ), .B(\CARRYB[25][69] ), .CI(\SUMB[25][70] ), 
        .CO(\CARRYB[26][69] ), .S(\SUMB[26][69] ) );
  FA1A S2_26_70 ( .A(\ab[26][70] ), .B(\CARRYB[25][70] ), .CI(\SUMB[25][71] ), 
        .CO(\CARRYB[26][70] ), .S(\SUMB[26][70] ) );
  FA1A S2_25_57 ( .A(\ab[25][57] ), .B(\CARRYB[24][57] ), .CI(\SUMB[24][58] ), 
        .CO(\CARRYB[25][57] ), .S(\SUMB[25][57] ) );
  FA1A S2_23_76 ( .A(\ab[23][76] ), .B(\CARRYB[22][76] ), .CI(\SUMB[22][77] ), 
        .CO(\CARRYB[23][76] ), .S(\SUMB[23][76] ) );
  FA1A S2_23_75 ( .A(\ab[23][75] ), .B(\CARRYB[22][75] ), .CI(\SUMB[22][76] ), 
        .CO(\CARRYB[23][75] ), .S(\SUMB[23][75] ) );
  FA1A S2_23_74 ( .A(\ab[23][74] ), .B(\CARRYB[22][74] ), .CI(\SUMB[22][75] ), 
        .CO(\CARRYB[23][74] ), .S(\SUMB[23][74] ) );
  FA1A S2_25_69 ( .A(\ab[25][69] ), .B(\CARRYB[24][69] ), .CI(\SUMB[24][70] ), 
        .CO(\CARRYB[25][69] ), .S(\SUMB[25][69] ) );
  FA1A S2_25_70 ( .A(\ab[25][70] ), .B(\CARRYB[24][70] ), .CI(\SUMB[24][71] ), 
        .CO(\CARRYB[25][70] ), .S(\SUMB[25][70] ) );
  FA1A S2_25_71 ( .A(\ab[25][71] ), .B(\CARRYB[24][71] ), .CI(\SUMB[24][72] ), 
        .CO(\CARRYB[25][71] ), .S(\SUMB[25][71] ) );
  FA1A S2_24_57 ( .A(\ab[24][57] ), .B(\CARRYB[23][57] ), .CI(\SUMB[23][58] ), 
        .CO(\CARRYB[24][57] ), .S(\SUMB[24][57] ) );
  FA1A S2_22_77 ( .A(\ab[22][77] ), .B(\CARRYB[21][77] ), .CI(\SUMB[21][78] ), 
        .CO(\CARRYB[22][77] ), .S(\SUMB[22][77] ) );
  FA1A S2_22_76 ( .A(\ab[22][76] ), .B(\CARRYB[21][76] ), .CI(\SUMB[21][77] ), 
        .CO(\CARRYB[22][76] ), .S(\SUMB[22][76] ) );
  FA1A S2_22_75 ( .A(\ab[22][75] ), .B(\CARRYB[21][75] ), .CI(\SUMB[21][76] ), 
        .CO(\CARRYB[22][75] ), .S(\SUMB[22][75] ) );
  FA1A S2_24_69 ( .A(\ab[24][69] ), .B(\CARRYB[23][69] ), .CI(\SUMB[23][70] ), 
        .CO(\CARRYB[24][69] ), .S(\SUMB[24][69] ) );
  FA1A S2_24_70 ( .A(\ab[24][70] ), .B(\CARRYB[23][70] ), .CI(\SUMB[23][71] ), 
        .CO(\CARRYB[24][70] ), .S(\SUMB[24][70] ) );
  FA1A S2_24_71 ( .A(\ab[24][71] ), .B(\CARRYB[23][71] ), .CI(\SUMB[23][72] ), 
        .CO(\CARRYB[24][71] ), .S(\SUMB[24][71] ) );
  FA1A S2_24_72 ( .A(\ab[24][72] ), .B(\CARRYB[23][72] ), .CI(\SUMB[23][73] ), 
        .CO(\CARRYB[24][72] ), .S(\SUMB[24][72] ) );
  FA1A S2_21_78 ( .A(\ab[21][78] ), .B(\CARRYB[20][78] ), .CI(\SUMB[20][79] ), 
        .CO(\CARRYB[21][78] ), .S(\SUMB[21][78] ) );
  FA1A S2_21_77 ( .A(\ab[21][77] ), .B(\CARRYB[20][77] ), .CI(\SUMB[20][78] ), 
        .CO(\CARRYB[21][77] ), .S(\SUMB[21][77] ) );
  FA1A S2_21_76 ( .A(\ab[21][76] ), .B(\CARRYB[20][76] ), .CI(\SUMB[20][77] ), 
        .CO(\CARRYB[21][76] ), .S(\SUMB[21][76] ) );
  FA1A S2_23_69 ( .A(\ab[23][69] ), .B(\CARRYB[22][69] ), .CI(\SUMB[22][70] ), 
        .CO(\CARRYB[23][69] ), .S(\SUMB[23][69] ) );
  FA1A S2_23_70 ( .A(\ab[23][70] ), .B(\CARRYB[22][70] ), .CI(\SUMB[22][71] ), 
        .CO(\CARRYB[23][70] ), .S(\SUMB[23][70] ) );
  FA1A S2_23_71 ( .A(\ab[23][71] ), .B(\CARRYB[22][71] ), .CI(\SUMB[22][72] ), 
        .CO(\CARRYB[23][71] ), .S(\SUMB[23][71] ) );
  FA1A S2_23_72 ( .A(\ab[23][72] ), .B(\CARRYB[22][72] ), .CI(\SUMB[22][73] ), 
        .CO(\CARRYB[23][72] ), .S(\SUMB[23][72] ) );
  FA1A S2_23_73 ( .A(\ab[23][73] ), .B(\CARRYB[22][73] ), .CI(\SUMB[22][74] ), 
        .CO(\CARRYB[23][73] ), .S(\SUMB[23][73] ) );
  FA1A S2_23_57 ( .A(\ab[23][57] ), .B(\CARRYB[22][57] ), .CI(\SUMB[22][58] ), 
        .CO(\CARRYB[23][57] ), .S(\SUMB[23][57] ) );
  FA1A S2_20_79 ( .A(\ab[20][79] ), .B(\CARRYB[19][79] ), .CI(\SUMB[19][80] ), 
        .CO(\CARRYB[20][79] ), .S(\SUMB[20][79] ) );
  FA1A S2_20_78 ( .A(\ab[20][78] ), .B(\CARRYB[19][78] ), .CI(\SUMB[19][79] ), 
        .CO(\CARRYB[20][78] ), .S(\SUMB[20][78] ) );
  FA1A S2_20_77 ( .A(\ab[20][77] ), .B(\CARRYB[19][77] ), .CI(\SUMB[19][78] ), 
        .CO(\CARRYB[20][77] ), .S(\SUMB[20][77] ) );
  FA1A S2_22_70 ( .A(\ab[22][70] ), .B(\CARRYB[21][70] ), .CI(\SUMB[21][71] ), 
        .CO(\CARRYB[22][70] ), .S(\SUMB[22][70] ) );
  FA1A S2_22_71 ( .A(\ab[22][71] ), .B(\CARRYB[21][71] ), .CI(\SUMB[21][72] ), 
        .CO(\CARRYB[22][71] ), .S(\SUMB[22][71] ) );
  FA1A S2_22_72 ( .A(\ab[22][72] ), .B(\CARRYB[21][72] ), .CI(\SUMB[21][73] ), 
        .CO(\CARRYB[22][72] ), .S(\SUMB[22][72] ) );
  FA1A S2_22_73 ( .A(\ab[22][73] ), .B(\CARRYB[21][73] ), .CI(\SUMB[21][74] ), 
        .CO(\CARRYB[22][73] ), .S(\SUMB[22][73] ) );
  FA1A S2_22_74 ( .A(\ab[22][74] ), .B(\CARRYB[21][74] ), .CI(\SUMB[21][75] ), 
        .CO(\CARRYB[22][74] ), .S(\SUMB[22][74] ) );
  FA1A S2_19_79 ( .A(\ab[19][79] ), .B(\CARRYB[18][79] ), .CI(\SUMB[18][80] ), 
        .CO(\CARRYB[19][79] ), .S(\SUMB[19][79] ) );
  FA1A S2_19_78 ( .A(\ab[19][78] ), .B(\CARRYB[18][78] ), .CI(\SUMB[18][79] ), 
        .CO(\CARRYB[19][78] ), .S(\SUMB[19][78] ) );
  FA1A S2_21_71 ( .A(\ab[21][71] ), .B(\CARRYB[20][71] ), .CI(\SUMB[20][72] ), 
        .CO(\CARRYB[21][71] ), .S(\SUMB[21][71] ) );
  FA1A S2_21_72 ( .A(\ab[21][72] ), .B(\CARRYB[20][72] ), .CI(\SUMB[20][73] ), 
        .CO(\CARRYB[21][72] ), .S(\SUMB[21][72] ) );
  FA1A S2_21_73 ( .A(\ab[21][73] ), .B(\CARRYB[20][73] ), .CI(\SUMB[20][74] ), 
        .CO(\CARRYB[21][73] ), .S(\SUMB[21][73] ) );
  FA1A S2_21_74 ( .A(\ab[21][74] ), .B(\CARRYB[20][74] ), .CI(\SUMB[20][75] ), 
        .CO(\CARRYB[21][74] ), .S(\SUMB[21][74] ) );
  FA1A S2_21_75 ( .A(\ab[21][75] ), .B(\CARRYB[20][75] ), .CI(\SUMB[20][76] ), 
        .CO(\CARRYB[21][75] ), .S(\SUMB[21][75] ) );
  FA1A S2_18_79 ( .A(\ab[18][79] ), .B(\CARRYB[17][79] ), .CI(\SUMB[17][80] ), 
        .CO(\CARRYB[18][79] ), .S(\SUMB[18][79] ) );
  FA1A S2_20_72 ( .A(\ab[20][72] ), .B(\CARRYB[19][72] ), .CI(\SUMB[19][73] ), 
        .CO(\CARRYB[20][72] ), .S(\SUMB[20][72] ) );
  FA1A S2_20_73 ( .A(\ab[20][73] ), .B(\CARRYB[19][73] ), .CI(\SUMB[19][74] ), 
        .CO(\CARRYB[20][73] ), .S(\SUMB[20][73] ) );
  FA1A S2_20_74 ( .A(\ab[20][74] ), .B(\CARRYB[19][74] ), .CI(\SUMB[19][75] ), 
        .CO(\CARRYB[20][74] ), .S(\SUMB[20][74] ) );
  FA1A S2_20_75 ( .A(\ab[20][75] ), .B(\CARRYB[19][75] ), .CI(\SUMB[19][76] ), 
        .CO(\CARRYB[20][75] ), .S(\SUMB[20][75] ) );
  FA1A S2_20_76 ( .A(\ab[20][76] ), .B(\CARRYB[19][76] ), .CI(\SUMB[19][77] ), 
        .CO(\CARRYB[20][76] ), .S(\SUMB[20][76] ) );
  FA1A S2_22_69 ( .A(\ab[22][69] ), .B(\CARRYB[21][69] ), .CI(\SUMB[21][70] ), 
        .CO(\CARRYB[22][69] ), .S(\SUMB[22][69] ) );
  FA1A S2_22_57 ( .A(\ab[22][57] ), .B(\CARRYB[21][57] ), .CI(\SUMB[21][58] ), 
        .CO(\CARRYB[22][57] ), .S(\SUMB[22][57] ) );
  FA1A S2_19_73 ( .A(\ab[19][73] ), .B(\CARRYB[18][73] ), .CI(\SUMB[18][74] ), 
        .CO(\CARRYB[19][73] ), .S(\SUMB[19][73] ) );
  FA1A S2_19_74 ( .A(\ab[19][74] ), .B(\CARRYB[18][74] ), .CI(\SUMB[18][75] ), 
        .CO(\CARRYB[19][74] ), .S(\SUMB[19][74] ) );
  FA1A S2_19_75 ( .A(\ab[19][75] ), .B(\CARRYB[18][75] ), .CI(\SUMB[18][76] ), 
        .CO(\CARRYB[19][75] ), .S(\SUMB[19][75] ) );
  FA1A S2_19_76 ( .A(\ab[19][76] ), .B(\CARRYB[18][76] ), .CI(\SUMB[18][77] ), 
        .CO(\CARRYB[19][76] ), .S(\SUMB[19][76] ) );
  FA1A S2_19_77 ( .A(\ab[19][77] ), .B(\CARRYB[18][77] ), .CI(\SUMB[18][78] ), 
        .CO(\CARRYB[19][77] ), .S(\SUMB[19][77] ) );
  FA1A S2_21_69 ( .A(\ab[21][69] ), .B(\CARRYB[20][69] ), .CI(\SUMB[20][70] ), 
        .CO(\CARRYB[21][69] ), .S(\SUMB[21][69] ) );
  FA1A S2_21_70 ( .A(\ab[21][70] ), .B(\CARRYB[20][70] ), .CI(\SUMB[20][71] ), 
        .CO(\CARRYB[21][70] ), .S(\SUMB[21][70] ) );
  FA1A S2_21_57 ( .A(\ab[21][57] ), .B(\CARRYB[20][57] ), .CI(\SUMB[20][58] ), 
        .CO(\CARRYB[21][57] ), .S(\SUMB[21][57] ) );
  FA1A S2_18_74 ( .A(\ab[18][74] ), .B(\CARRYB[17][74] ), .CI(\SUMB[17][75] ), 
        .CO(\CARRYB[18][74] ), .S(\SUMB[18][74] ) );
  FA1A S2_18_75 ( .A(\ab[18][75] ), .B(\CARRYB[17][75] ), .CI(\SUMB[17][76] ), 
        .CO(\CARRYB[18][75] ), .S(\SUMB[18][75] ) );
  FA1A S2_18_76 ( .A(\ab[18][76] ), .B(\CARRYB[17][76] ), .CI(\SUMB[17][77] ), 
        .CO(\CARRYB[18][76] ), .S(\SUMB[18][76] ) );
  FA1A S2_18_77 ( .A(\ab[18][77] ), .B(\CARRYB[17][77] ), .CI(\SUMB[17][78] ), 
        .CO(\CARRYB[18][77] ), .S(\SUMB[18][77] ) );
  FA1A S2_18_78 ( .A(\ab[18][78] ), .B(\CARRYB[17][78] ), .CI(\SUMB[17][79] ), 
        .CO(\CARRYB[18][78] ), .S(\SUMB[18][78] ) );
  FA1A S2_20_69 ( .A(\ab[20][69] ), .B(\CARRYB[19][69] ), .CI(\SUMB[19][70] ), 
        .CO(\CARRYB[20][69] ), .S(\SUMB[20][69] ) );
  FA1A S2_20_70 ( .A(\ab[20][70] ), .B(\CARRYB[19][70] ), .CI(\SUMB[19][71] ), 
        .CO(\CARRYB[20][70] ), .S(\SUMB[20][70] ) );
  FA1A S2_20_71 ( .A(\ab[20][71] ), .B(\CARRYB[19][71] ), .CI(\SUMB[19][72] ), 
        .CO(\CARRYB[20][71] ), .S(\SUMB[20][71] ) );
  FA1A S2_20_57 ( .A(\ab[20][57] ), .B(\CARRYB[19][57] ), .CI(\SUMB[19][58] ), 
        .CO(\CARRYB[20][57] ), .S(\SUMB[20][57] ) );
  FA1A S2_17_75 ( .A(\ab[17][75] ), .B(\CARRYB[16][75] ), .CI(\SUMB[16][76] ), 
        .CO(\CARRYB[17][75] ), .S(\SUMB[17][75] ) );
  FA1A S2_17_76 ( .A(\ab[17][76] ), .B(\CARRYB[16][76] ), .CI(\SUMB[16][77] ), 
        .CO(\CARRYB[17][76] ), .S(\SUMB[17][76] ) );
  FA1A S2_17_77 ( .A(\ab[17][77] ), .B(\CARRYB[16][77] ), .CI(\SUMB[16][78] ), 
        .CO(\CARRYB[17][77] ), .S(\SUMB[17][77] ) );
  FA1A S2_17_78 ( .A(\ab[17][78] ), .B(\CARRYB[16][78] ), .CI(\SUMB[16][79] ), 
        .CO(\CARRYB[17][78] ), .S(\SUMB[17][78] ) );
  FA1A S2_17_79 ( .A(\ab[17][79] ), .B(\CARRYB[16][79] ), .CI(\SUMB[16][80] ), 
        .CO(\CARRYB[17][79] ), .S(\SUMB[17][79] ) );
  FA1A S2_19_70 ( .A(\ab[19][70] ), .B(\CARRYB[18][70] ), .CI(\SUMB[18][71] ), 
        .CO(\CARRYB[19][70] ), .S(\SUMB[19][70] ) );
  FA1A S2_19_69 ( .A(\ab[19][69] ), .B(\CARRYB[18][69] ), .CI(\SUMB[18][70] ), 
        .CO(\CARRYB[19][69] ), .S(\SUMB[19][69] ) );
  FA1A S2_19_71 ( .A(\ab[19][71] ), .B(\CARRYB[18][71] ), .CI(\SUMB[18][72] ), 
        .CO(\CARRYB[19][71] ), .S(\SUMB[19][71] ) );
  FA1A S2_19_72 ( .A(\ab[19][72] ), .B(\CARRYB[18][72] ), .CI(\SUMB[18][73] ), 
        .CO(\CARRYB[19][72] ), .S(\SUMB[19][72] ) );
  FA1A S2_19_57 ( .A(\ab[19][57] ), .B(\CARRYB[18][57] ), .CI(\SUMB[18][58] ), 
        .CO(\CARRYB[19][57] ), .S(\SUMB[19][57] ) );
  FA1A S2_16_76 ( .A(\ab[16][76] ), .B(\CARRYB[15][76] ), .CI(\SUMB[15][77] ), 
        .CO(\CARRYB[16][76] ), .S(\SUMB[16][76] ) );
  FA1A S2_16_77 ( .A(\ab[16][77] ), .B(\CARRYB[15][77] ), .CI(\SUMB[15][78] ), 
        .CO(\CARRYB[16][77] ), .S(\SUMB[16][77] ) );
  FA1A S2_16_78 ( .A(\ab[16][78] ), .B(\CARRYB[15][78] ), .CI(\SUMB[15][79] ), 
        .CO(\CARRYB[16][78] ), .S(\SUMB[16][78] ) );
  FA1A S2_16_79 ( .A(\ab[16][79] ), .B(\CARRYB[15][79] ), .CI(\SUMB[15][80] ), 
        .CO(\CARRYB[16][79] ), .S(\SUMB[16][79] ) );
  FA1A S2_18_71 ( .A(\ab[18][71] ), .B(\CARRYB[17][71] ), .CI(\SUMB[17][72] ), 
        .CO(\CARRYB[18][71] ), .S(\SUMB[18][71] ) );
  FA1A S2_18_70 ( .A(\ab[18][70] ), .B(\CARRYB[17][70] ), .CI(\SUMB[17][71] ), 
        .CO(\CARRYB[18][70] ), .S(\SUMB[18][70] ) );
  FA1A S2_18_69 ( .A(\ab[18][69] ), .B(\CARRYB[17][69] ), .CI(\SUMB[17][70] ), 
        .CO(\CARRYB[18][69] ), .S(\SUMB[18][69] ) );
  FA1A S2_18_72 ( .A(\ab[18][72] ), .B(\CARRYB[17][72] ), .CI(\SUMB[17][73] ), 
        .CO(\CARRYB[18][72] ), .S(\SUMB[18][72] ) );
  FA1A S2_18_73 ( .A(\ab[18][73] ), .B(\CARRYB[17][73] ), .CI(\SUMB[17][74] ), 
        .CO(\CARRYB[18][73] ), .S(\SUMB[18][73] ) );
  FA1A S2_18_57 ( .A(\ab[18][57] ), .B(\CARRYB[17][57] ), .CI(\SUMB[17][58] ), 
        .CO(\CARRYB[18][57] ), .S(\SUMB[18][57] ) );
  FA1A S2_15_77 ( .A(\ab[15][77] ), .B(\CARRYB[14][77] ), .CI(\SUMB[14][78] ), 
        .CO(\CARRYB[15][77] ), .S(\SUMB[15][77] ) );
  FA1A S2_15_78 ( .A(\ab[15][78] ), .B(\CARRYB[14][78] ), .CI(\SUMB[14][79] ), 
        .CO(\CARRYB[15][78] ), .S(\SUMB[15][78] ) );
  FA1A S2_15_79 ( .A(\ab[15][79] ), .B(\CARRYB[14][79] ), .CI(\SUMB[14][80] ), 
        .CO(\CARRYB[15][79] ), .S(\SUMB[15][79] ) );
  FA1A S2_17_72 ( .A(\ab[17][72] ), .B(\CARRYB[16][72] ), .CI(\SUMB[16][73] ), 
        .CO(\CARRYB[17][72] ), .S(\SUMB[17][72] ) );
  FA1A S2_17_71 ( .A(\ab[17][71] ), .B(\CARRYB[16][71] ), .CI(\SUMB[16][72] ), 
        .CO(\CARRYB[17][71] ), .S(\SUMB[17][71] ) );
  FA1A S2_17_70 ( .A(\ab[17][70] ), .B(\CARRYB[16][70] ), .CI(\SUMB[16][71] ), 
        .CO(\CARRYB[17][70] ), .S(\SUMB[17][70] ) );
  FA1A S2_17_69 ( .A(\ab[17][69] ), .B(\CARRYB[16][69] ), .CI(\SUMB[16][70] ), 
        .CO(\CARRYB[17][69] ), .S(\SUMB[17][69] ) );
  FA1A S2_17_73 ( .A(\ab[17][73] ), .B(\CARRYB[16][73] ), .CI(\SUMB[16][74] ), 
        .CO(\CARRYB[17][73] ), .S(\SUMB[17][73] ) );
  FA1A S2_17_74 ( .A(\ab[17][74] ), .B(\CARRYB[16][74] ), .CI(\SUMB[16][75] ), 
        .CO(\CARRYB[17][74] ), .S(\SUMB[17][74] ) );
  FA1A S2_17_57 ( .A(\ab[17][57] ), .B(\CARRYB[16][57] ), .CI(\SUMB[16][58] ), 
        .CO(\CARRYB[17][57] ), .S(\SUMB[17][57] ) );
  FA1A S2_16_73 ( .A(\ab[16][73] ), .B(\CARRYB[15][73] ), .CI(\SUMB[15][74] ), 
        .CO(\CARRYB[16][73] ), .S(\SUMB[16][73] ) );
  FA1A S2_16_72 ( .A(\ab[16][72] ), .B(\CARRYB[15][72] ), .CI(\SUMB[15][73] ), 
        .CO(\CARRYB[16][72] ), .S(\SUMB[16][72] ) );
  FA1A S2_16_71 ( .A(\ab[16][71] ), .B(\CARRYB[15][71] ), .CI(\SUMB[15][72] ), 
        .CO(\CARRYB[16][71] ), .S(\SUMB[16][71] ) );
  FA1A S2_16_70 ( .A(\ab[16][70] ), .B(\CARRYB[15][70] ), .CI(\SUMB[15][71] ), 
        .CO(\CARRYB[16][70] ), .S(\SUMB[16][70] ) );
  FA1A S2_16_69 ( .A(\ab[16][69] ), .B(\CARRYB[15][69] ), .CI(\SUMB[15][70] ), 
        .CO(\CARRYB[16][69] ), .S(\SUMB[16][69] ) );
  FA1A S2_16_74 ( .A(\ab[16][74] ), .B(\CARRYB[15][74] ), .CI(\SUMB[15][75] ), 
        .CO(\CARRYB[16][74] ), .S(\SUMB[16][74] ) );
  FA1A S2_16_75 ( .A(\ab[16][75] ), .B(\CARRYB[15][75] ), .CI(\SUMB[15][76] ), 
        .CO(\CARRYB[16][75] ), .S(\SUMB[16][75] ) );
  FA1A S2_16_57 ( .A(\ab[16][57] ), .B(\CARRYB[15][57] ), .CI(\SUMB[15][58] ), 
        .CO(\CARRYB[16][57] ), .S(\SUMB[16][57] ) );
  FA1A S2_15_74 ( .A(\ab[15][74] ), .B(\CARRYB[14][74] ), .CI(\SUMB[14][75] ), 
        .CO(\CARRYB[15][74] ), .S(\SUMB[15][74] ) );
  FA1A S2_15_73 ( .A(\ab[15][73] ), .B(\CARRYB[14][73] ), .CI(\SUMB[14][74] ), 
        .CO(\CARRYB[15][73] ), .S(\SUMB[15][73] ) );
  FA1A S2_15_72 ( .A(\ab[15][72] ), .B(\CARRYB[14][72] ), .CI(\SUMB[14][73] ), 
        .CO(\CARRYB[15][72] ), .S(\SUMB[15][72] ) );
  FA1A S2_15_71 ( .A(\ab[15][71] ), .B(\CARRYB[14][71] ), .CI(\SUMB[14][72] ), 
        .CO(\CARRYB[15][71] ), .S(\SUMB[15][71] ) );
  FA1A S2_15_70 ( .A(\ab[15][70] ), .B(\CARRYB[14][70] ), .CI(\SUMB[14][71] ), 
        .CO(\CARRYB[15][70] ), .S(\SUMB[15][70] ) );
  FA1A S2_15_69 ( .A(\ab[15][69] ), .B(\CARRYB[14][69] ), .CI(\SUMB[14][70] ), 
        .CO(\CARRYB[15][69] ), .S(\SUMB[15][69] ) );
  FA1A S2_15_75 ( .A(\ab[15][75] ), .B(\CARRYB[14][75] ), .CI(\SUMB[14][76] ), 
        .CO(\CARRYB[15][75] ), .S(\SUMB[15][75] ) );
  FA1A S2_15_76 ( .A(\ab[15][76] ), .B(\CARRYB[14][76] ), .CI(\SUMB[14][77] ), 
        .CO(\CARRYB[15][76] ), .S(\SUMB[15][76] ) );
  FA1A S2_15_57 ( .A(\ab[15][57] ), .B(\CARRYB[14][57] ), .CI(\SUMB[14][58] ), 
        .CO(\CARRYB[15][57] ), .S(\SUMB[15][57] ) );
  FA1A S4_79 ( .A(\ab[29][79] ), .B(\CARRYB[28][79] ), .CI(\SUMB[28][80] ), 
        .CO(\CARRYB[29][79] ), .S(\SUMB[29][79] ) );
  FA1A S4_72 ( .A(\ab[29][72] ), .B(\CARRYB[28][72] ), .CI(\SUMB[28][73] ), 
        .CO(\CARRYB[29][72] ), .S(\SUMB[29][72] ) );
  FA1A S4_76 ( .A(\ab[29][76] ), .B(\CARRYB[28][76] ), .CI(\SUMB[28][77] ), 
        .CO(\CARRYB[29][76] ), .S(\SUMB[29][76] ) );
  FA1A S4_74 ( .A(\ab[29][74] ), .B(\CARRYB[28][74] ), .CI(\SUMB[28][75] ), 
        .CO(\CARRYB[29][74] ), .S(\SUMB[29][74] ) );
  FA1A S4_70 ( .A(\ab[29][70] ), .B(\CARRYB[28][70] ), .CI(\SUMB[28][71] ), 
        .CO(\CARRYB[29][70] ), .S(\SUMB[29][70] ) );
  FA1A S2_28_56 ( .A(\ab[28][56] ), .B(\CARRYB[27][56] ), .CI(\SUMB[27][57] ), 
        .CO(\CARRYB[28][56] ), .S(\SUMB[28][56] ) );
  FA1A S4_54 ( .A(\ab[29][54] ), .B(\CARRYB[28][54] ), .CI(\SUMB[28][55] ), 
        .CO(\CARRYB[29][54] ), .S(\SUMB[29][54] ) );
  FA1A S4_53 ( .A(\ab[29][53] ), .B(\CARRYB[28][53] ), .CI(\SUMB[28][54] ), 
        .CO(\CARRYB[29][53] ), .S(\SUMB[29][53] ) );
  FA1A S4_64 ( .A(\ab[29][64] ), .B(\CARRYB[28][64] ), .CI(\SUMB[28][65] ), 
        .CO(\CARRYB[29][64] ), .S(\SUMB[29][64] ) );
  FA1A S4_65 ( .A(\ab[29][65] ), .B(\CARRYB[28][65] ), .CI(\SUMB[28][66] ), 
        .CO(\CARRYB[29][65] ), .S(\SUMB[29][65] ) );
  FA1A S4_66 ( .A(\ab[29][66] ), .B(\CARRYB[28][66] ), .CI(\SUMB[28][67] ), 
        .CO(\CARRYB[29][66] ), .S(\SUMB[29][66] ) );
  FA1A S4_67 ( .A(\ab[29][67] ), .B(\CARRYB[28][67] ), .CI(\SUMB[28][68] ), 
        .CO(\CARRYB[29][67] ), .S(\SUMB[29][67] ) );
  FA1A S4_58 ( .A(\ab[29][58] ), .B(\CARRYB[28][58] ), .CI(\SUMB[28][59] ), 
        .CO(\CARRYB[29][58] ), .S(\SUMB[29][58] ) );
  FA1A S2_28_55 ( .A(\ab[28][55] ), .B(\CARRYB[27][55] ), .CI(\SUMB[27][56] ), 
        .CO(\CARRYB[28][55] ), .S(\SUMB[28][55] ) );
  FA1A S2_28_54 ( .A(\ab[28][54] ), .B(\CARRYB[27][54] ), .CI(\SUMB[27][55] ), 
        .CO(\CARRYB[28][54] ), .S(\SUMB[28][54] ) );
  FA1A S2_28_53 ( .A(\ab[28][53] ), .B(\CARRYB[27][53] ), .CI(\SUMB[27][54] ), 
        .CO(\CARRYB[28][53] ), .S(\SUMB[28][53] ) );
  FA1A S2_28_59 ( .A(\ab[28][59] ), .B(\CARRYB[27][59] ), .CI(\SUMB[27][60] ), 
        .CO(\CARRYB[28][59] ), .S(\SUMB[28][59] ) );
  FA1A S2_28_64 ( .A(\ab[28][64] ), .B(\CARRYB[27][64] ), .CI(\SUMB[27][65] ), 
        .CO(\CARRYB[28][64] ), .S(\SUMB[28][64] ) );
  FA1A S2_28_65 ( .A(\ab[28][65] ), .B(\CARRYB[27][65] ), .CI(\SUMB[27][66] ), 
        .CO(\CARRYB[28][65] ), .S(\SUMB[28][65] ) );
  FA1A S2_28_66 ( .A(\ab[28][66] ), .B(\CARRYB[27][66] ), .CI(\SUMB[27][67] ), 
        .CO(\CARRYB[28][66] ), .S(\SUMB[28][66] ) );
  FA1A S2_28_67 ( .A(\ab[28][67] ), .B(\CARRYB[27][67] ), .CI(\SUMB[27][68] ), 
        .CO(\CARRYB[28][67] ), .S(\SUMB[28][67] ) );
  FA1A S2_28_68 ( .A(\ab[28][68] ), .B(\CARRYB[27][68] ), .CI(\SUMB[27][69] ), 
        .CO(\CARRYB[28][68] ), .S(\SUMB[28][68] ) );
  FA1A S2_28_58 ( .A(\ab[28][58] ), .B(\CARRYB[27][58] ), .CI(\SUMB[27][59] ), 
        .CO(\CARRYB[28][58] ), .S(\SUMB[28][58] ) );
  FA1A S2_27_56 ( .A(\ab[27][56] ), .B(\CARRYB[26][56] ), .CI(\SUMB[26][57] ), 
        .CO(\CARRYB[27][56] ), .S(\SUMB[27][56] ) );
  FA1A S2_27_55 ( .A(\ab[27][55] ), .B(\CARRYB[26][55] ), .CI(\SUMB[26][56] ), 
        .CO(\CARRYB[27][55] ), .S(\SUMB[27][55] ) );
  FA1A S2_27_54 ( .A(\ab[27][54] ), .B(\CARRYB[26][54] ), .CI(\SUMB[26][55] ), 
        .CO(\CARRYB[27][54] ), .S(\SUMB[27][54] ) );
  FA1A S2_27_59 ( .A(\ab[27][59] ), .B(\CARRYB[26][59] ), .CI(\SUMB[26][60] ), 
        .CO(\CARRYB[27][59] ), .S(\SUMB[27][59] ) );
  FA1A S2_27_65 ( .A(\ab[27][65] ), .B(\CARRYB[26][65] ), .CI(\SUMB[26][66] ), 
        .CO(\CARRYB[27][65] ), .S(\SUMB[27][65] ) );
  FA1A S2_27_66 ( .A(\ab[27][66] ), .B(\CARRYB[26][66] ), .CI(\SUMB[26][67] ), 
        .CO(\CARRYB[27][66] ), .S(\SUMB[27][66] ) );
  FA1A S2_27_67 ( .A(\ab[27][67] ), .B(\CARRYB[26][67] ), .CI(\SUMB[26][68] ), 
        .CO(\CARRYB[27][67] ), .S(\SUMB[27][67] ) );
  FA1A S2_27_68 ( .A(\ab[27][68] ), .B(\CARRYB[26][68] ), .CI(\SUMB[26][69] ), 
        .CO(\CARRYB[27][68] ), .S(\SUMB[27][68] ) );
  FA1A S2_27_58 ( .A(\ab[27][58] ), .B(\CARRYB[26][58] ), .CI(\SUMB[26][59] ), 
        .CO(\CARRYB[27][58] ), .S(\SUMB[27][58] ) );
  FA1A S4_60 ( .A(\ab[29][60] ), .B(\CARRYB[28][60] ), .CI(\SUMB[28][61] ), 
        .CO(\CARRYB[29][60] ), .S(\SUMB[29][60] ) );
  FA1A S2_27_53 ( .A(\ab[27][53] ), .B(\CARRYB[26][53] ), .CI(\SUMB[26][54] ), 
        .CO(\CARRYB[27][53] ), .S(\SUMB[27][53] ) );
  FA1A S2_26_56 ( .A(\ab[26][56] ), .B(\CARRYB[25][56] ), .CI(\SUMB[25][57] ), 
        .CO(\CARRYB[26][56] ), .S(\SUMB[26][56] ) );
  FA1A S2_26_55 ( .A(\ab[26][55] ), .B(\CARRYB[25][55] ), .CI(\SUMB[25][56] ), 
        .CO(\CARRYB[26][55] ), .S(\SUMB[26][55] ) );
  FA1A S2_26_59 ( .A(\ab[26][59] ), .B(\CARRYB[25][59] ), .CI(\SUMB[25][60] ), 
        .CO(\CARRYB[26][59] ), .S(\SUMB[26][59] ) );
  FA1A S2_26_66 ( .A(\ab[26][66] ), .B(\CARRYB[25][66] ), .CI(\SUMB[25][67] ), 
        .CO(\CARRYB[26][66] ), .S(\SUMB[26][66] ) );
  FA1A S2_26_67 ( .A(\ab[26][67] ), .B(\CARRYB[25][67] ), .CI(\SUMB[25][68] ), 
        .CO(\CARRYB[26][67] ), .S(\SUMB[26][67] ) );
  FA1A S2_26_68 ( .A(\ab[26][68] ), .B(\CARRYB[25][68] ), .CI(\SUMB[25][69] ), 
        .CO(\CARRYB[26][68] ), .S(\SUMB[26][68] ) );
  FA1A S2_26_58 ( .A(\ab[26][58] ), .B(\CARRYB[25][58] ), .CI(\SUMB[25][59] ), 
        .CO(\CARRYB[26][58] ), .S(\SUMB[26][58] ) );
  FA1A S2_28_60 ( .A(\ab[28][60] ), .B(\CARRYB[27][60] ), .CI(\SUMB[27][61] ), 
        .CO(\CARRYB[28][60] ), .S(\SUMB[28][60] ) );
  FA1A S2_26_54 ( .A(\ab[26][54] ), .B(\CARRYB[25][54] ), .CI(\SUMB[25][55] ), 
        .CO(\CARRYB[26][54] ), .S(\SUMB[26][54] ) );
  FA1A S2_25_56 ( .A(\ab[25][56] ), .B(\CARRYB[24][56] ), .CI(\SUMB[24][57] ), 
        .CO(\CARRYB[25][56] ), .S(\SUMB[25][56] ) );
  FA1A S2_25_59 ( .A(\ab[25][59] ), .B(\CARRYB[24][59] ), .CI(\SUMB[24][60] ), 
        .CO(\CARRYB[25][59] ), .S(\SUMB[25][59] ) );
  FA1A S2_25_67 ( .A(\ab[25][67] ), .B(\CARRYB[24][67] ), .CI(\SUMB[24][68] ), 
        .CO(\CARRYB[25][67] ), .S(\SUMB[25][67] ) );
  FA1A S2_25_68 ( .A(\ab[25][68] ), .B(\CARRYB[24][68] ), .CI(\SUMB[24][69] ), 
        .CO(\CARRYB[25][68] ), .S(\SUMB[25][68] ) );
  FA1A S2_25_58 ( .A(\ab[25][58] ), .B(\CARRYB[24][58] ), .CI(\SUMB[24][59] ), 
        .CO(\CARRYB[25][58] ), .S(\SUMB[25][58] ) );
  FA1A S2_27_60 ( .A(\ab[27][60] ), .B(\CARRYB[26][60] ), .CI(\SUMB[26][61] ), 
        .CO(\CARRYB[27][60] ), .S(\SUMB[27][60] ) );
  FA1A S2_27_64 ( .A(\ab[27][64] ), .B(\CARRYB[26][64] ), .CI(\SUMB[26][65] ), 
        .CO(\CARRYB[27][64] ), .S(\SUMB[27][64] ) );
  FA1A S2_25_55 ( .A(\ab[25][55] ), .B(\CARRYB[24][55] ), .CI(\SUMB[24][56] ), 
        .CO(\CARRYB[25][55] ), .S(\SUMB[25][55] ) );
  FA1A S2_24_59 ( .A(\ab[24][59] ), .B(\CARRYB[23][59] ), .CI(\SUMB[23][60] ), 
        .CO(\CARRYB[24][59] ), .S(\SUMB[24][59] ) );
  FA1A S2_24_68 ( .A(\ab[24][68] ), .B(\CARRYB[23][68] ), .CI(\SUMB[23][69] ), 
        .CO(\CARRYB[24][68] ), .S(\SUMB[24][68] ) );
  FA1A S2_24_58 ( .A(\ab[24][58] ), .B(\CARRYB[23][58] ), .CI(\SUMB[23][59] ), 
        .CO(\CARRYB[24][58] ), .S(\SUMB[24][58] ) );
  FA1A S2_26_60 ( .A(\ab[26][60] ), .B(\CARRYB[25][60] ), .CI(\SUMB[25][61] ), 
        .CO(\CARRYB[26][60] ), .S(\SUMB[26][60] ) );
  FA1A S2_26_64 ( .A(\ab[26][64] ), .B(\CARRYB[25][64] ), .CI(\SUMB[25][65] ), 
        .CO(\CARRYB[26][64] ), .S(\SUMB[26][64] ) );
  FA1A S2_26_65 ( .A(\ab[26][65] ), .B(\CARRYB[25][65] ), .CI(\SUMB[25][66] ), 
        .CO(\CARRYB[26][65] ), .S(\SUMB[26][65] ) );
  FA1A S2_24_56 ( .A(\ab[24][56] ), .B(\CARRYB[23][56] ), .CI(\SUMB[23][57] ), 
        .CO(\CARRYB[24][56] ), .S(\SUMB[24][56] ) );
  FA1A S2_26_53 ( .A(\ab[26][53] ), .B(\CARRYB[25][53] ), .CI(\SUMB[25][54] ), 
        .CO(\CARRYB[26][53] ), .S(\SUMB[26][53] ) );
  FA1A S2_23_59 ( .A(\ab[23][59] ), .B(\CARRYB[22][59] ), .CI(\SUMB[22][60] ), 
        .CO(\CARRYB[23][59] ), .S(\SUMB[23][59] ) );
  FA1A S2_23_58 ( .A(\ab[23][58] ), .B(\CARRYB[22][58] ), .CI(\SUMB[22][59] ), 
        .CO(\CARRYB[23][58] ), .S(\SUMB[23][58] ) );
  FA1A S2_25_64 ( .A(\ab[25][64] ), .B(\CARRYB[24][64] ), .CI(\SUMB[24][65] ), 
        .CO(\CARRYB[25][64] ), .S(\SUMB[25][64] ) );
  FA1A S2_25_60 ( .A(\ab[25][60] ), .B(\CARRYB[24][60] ), .CI(\SUMB[24][61] ), 
        .CO(\CARRYB[25][60] ), .S(\SUMB[25][60] ) );
  FA1A S2_25_65 ( .A(\ab[25][65] ), .B(\CARRYB[24][65] ), .CI(\SUMB[24][66] ), 
        .CO(\CARRYB[25][65] ), .S(\SUMB[25][65] ) );
  FA1A S2_25_66 ( .A(\ab[25][66] ), .B(\CARRYB[24][66] ), .CI(\SUMB[24][67] ), 
        .CO(\CARRYB[25][66] ), .S(\SUMB[25][66] ) );
  FA1A S2_25_53 ( .A(\ab[25][53] ), .B(\CARRYB[24][53] ), .CI(\SUMB[24][54] ), 
        .CO(\CARRYB[25][53] ), .S(\SUMB[25][53] ) );
  FA1A S2_25_54 ( .A(\ab[25][54] ), .B(\CARRYB[24][54] ), .CI(\SUMB[24][55] ), 
        .CO(\CARRYB[25][54] ), .S(\SUMB[25][54] ) );
  FA1A S2_22_59 ( .A(\ab[22][59] ), .B(\CARRYB[21][59] ), .CI(\SUMB[21][60] ), 
        .CO(\CARRYB[22][59] ), .S(\SUMB[22][59] ) );
  FA1A S2_22_58 ( .A(\ab[22][58] ), .B(\CARRYB[21][58] ), .CI(\SUMB[21][59] ), 
        .CO(\CARRYB[22][58] ), .S(\SUMB[22][58] ) );
  FA1A S2_24_65 ( .A(\ab[24][65] ), .B(\CARRYB[23][65] ), .CI(\SUMB[23][66] ), 
        .CO(\CARRYB[24][65] ), .S(\SUMB[24][65] ) );
  FA1A S2_24_64 ( .A(\ab[24][64] ), .B(\CARRYB[23][64] ), .CI(\SUMB[23][65] ), 
        .CO(\CARRYB[24][64] ), .S(\SUMB[24][64] ) );
  FA1A S2_24_60 ( .A(\ab[24][60] ), .B(\CARRYB[23][60] ), .CI(\SUMB[23][61] ), 
        .CO(\CARRYB[24][60] ), .S(\SUMB[24][60] ) );
  FA1A S2_24_66 ( .A(\ab[24][66] ), .B(\CARRYB[23][66] ), .CI(\SUMB[23][67] ), 
        .CO(\CARRYB[24][66] ), .S(\SUMB[24][66] ) );
  FA1A S2_24_67 ( .A(\ab[24][67] ), .B(\CARRYB[23][67] ), .CI(\SUMB[23][68] ), 
        .CO(\CARRYB[24][67] ), .S(\SUMB[24][67] ) );
  FA1A S2_24_53 ( .A(\ab[24][53] ), .B(\CARRYB[23][53] ), .CI(\SUMB[23][54] ), 
        .CO(\CARRYB[24][53] ), .S(\SUMB[24][53] ) );
  FA1A S2_24_54 ( .A(\ab[24][54] ), .B(\CARRYB[23][54] ), .CI(\SUMB[23][55] ), 
        .CO(\CARRYB[24][54] ), .S(\SUMB[24][54] ) );
  FA1A S2_24_55 ( .A(\ab[24][55] ), .B(\CARRYB[23][55] ), .CI(\SUMB[23][56] ), 
        .CO(\CARRYB[24][55] ), .S(\SUMB[24][55] ) );
  FA1A S2_21_59 ( .A(\ab[21][59] ), .B(\CARRYB[20][59] ), .CI(\SUMB[20][60] ), 
        .CO(\CARRYB[21][59] ), .S(\SUMB[21][59] ) );
  FA1A S2_23_66 ( .A(\ab[23][66] ), .B(\CARRYB[22][66] ), .CI(\SUMB[22][67] ), 
        .CO(\CARRYB[23][66] ), .S(\SUMB[23][66] ) );
  FA1A S2_23_65 ( .A(\ab[23][65] ), .B(\CARRYB[22][65] ), .CI(\SUMB[22][66] ), 
        .CO(\CARRYB[23][65] ), .S(\SUMB[23][65] ) );
  FA1A S2_23_64 ( .A(\ab[23][64] ), .B(\CARRYB[22][64] ), .CI(\SUMB[22][65] ), 
        .CO(\CARRYB[23][64] ), .S(\SUMB[23][64] ) );
  FA1A S2_23_60 ( .A(\ab[23][60] ), .B(\CARRYB[22][60] ), .CI(\SUMB[22][61] ), 
        .CO(\CARRYB[23][60] ), .S(\SUMB[23][60] ) );
  FA1A S2_23_67 ( .A(\ab[23][67] ), .B(\CARRYB[22][67] ), .CI(\SUMB[22][68] ), 
        .CO(\CARRYB[23][67] ), .S(\SUMB[23][67] ) );
  FA1A S2_23_68 ( .A(\ab[23][68] ), .B(\CARRYB[22][68] ), .CI(\SUMB[22][69] ), 
        .CO(\CARRYB[23][68] ), .S(\SUMB[23][68] ) );
  FA1A S2_23_54 ( .A(\ab[23][54] ), .B(\CARRYB[22][54] ), .CI(\SUMB[22][55] ), 
        .CO(\CARRYB[23][54] ), .S(\SUMB[23][54] ) );
  FA1A S2_23_53 ( .A(\ab[23][53] ), .B(\CARRYB[22][53] ), .CI(\SUMB[22][54] ), 
        .CO(\CARRYB[23][53] ), .S(\SUMB[23][53] ) );
  FA1A S2_23_55 ( .A(\ab[23][55] ), .B(\CARRYB[22][55] ), .CI(\SUMB[22][56] ), 
        .CO(\CARRYB[23][55] ), .S(\SUMB[23][55] ) );
  FA1A S2_23_56 ( .A(\ab[23][56] ), .B(\CARRYB[22][56] ), .CI(\SUMB[22][57] ), 
        .CO(\CARRYB[23][56] ), .S(\SUMB[23][56] ) );
  FA1A S2_22_67 ( .A(\ab[22][67] ), .B(\CARRYB[21][67] ), .CI(\SUMB[21][68] ), 
        .CO(\CARRYB[22][67] ), .S(\SUMB[22][67] ) );
  FA1A S2_22_66 ( .A(\ab[22][66] ), .B(\CARRYB[21][66] ), .CI(\SUMB[21][67] ), 
        .CO(\CARRYB[22][66] ), .S(\SUMB[22][66] ) );
  FA1A S2_22_65 ( .A(\ab[22][65] ), .B(\CARRYB[21][65] ), .CI(\SUMB[21][66] ), 
        .CO(\CARRYB[22][65] ), .S(\SUMB[22][65] ) );
  FA1A S2_22_64 ( .A(\ab[22][64] ), .B(\CARRYB[21][64] ), .CI(\SUMB[21][65] ), 
        .CO(\CARRYB[22][64] ), .S(\SUMB[22][64] ) );
  FA1A S2_22_60 ( .A(\ab[22][60] ), .B(\CARRYB[21][60] ), .CI(\SUMB[21][61] ), 
        .CO(\CARRYB[22][60] ), .S(\SUMB[22][60] ) );
  FA1A S2_22_68 ( .A(\ab[22][68] ), .B(\CARRYB[21][68] ), .CI(\SUMB[21][69] ), 
        .CO(\CARRYB[22][68] ), .S(\SUMB[22][68] ) );
  FA1A S2_22_55 ( .A(\ab[22][55] ), .B(\CARRYB[21][55] ), .CI(\SUMB[21][56] ), 
        .CO(\CARRYB[22][55] ), .S(\SUMB[22][55] ) );
  FA1A S2_22_54 ( .A(\ab[22][54] ), .B(\CARRYB[21][54] ), .CI(\SUMB[21][55] ), 
        .CO(\CARRYB[22][54] ), .S(\SUMB[22][54] ) );
  FA1A S2_22_53 ( .A(\ab[22][53] ), .B(\CARRYB[21][53] ), .CI(\SUMB[21][54] ), 
        .CO(\CARRYB[22][53] ), .S(\SUMB[22][53] ) );
  FA1A S2_22_56 ( .A(\ab[22][56] ), .B(\CARRYB[21][56] ), .CI(\SUMB[21][57] ), 
        .CO(\CARRYB[22][56] ), .S(\SUMB[22][56] ) );
  FA1A S2_21_68 ( .A(\ab[21][68] ), .B(\CARRYB[20][68] ), .CI(\SUMB[20][69] ), 
        .CO(\CARRYB[21][68] ), .S(\SUMB[21][68] ) );
  FA1A S2_21_67 ( .A(\ab[21][67] ), .B(\CARRYB[20][67] ), .CI(\SUMB[20][68] ), 
        .CO(\CARRYB[21][67] ), .S(\SUMB[21][67] ) );
  FA1A S2_21_66 ( .A(\ab[21][66] ), .B(\CARRYB[20][66] ), .CI(\SUMB[20][67] ), 
        .CO(\CARRYB[21][66] ), .S(\SUMB[21][66] ) );
  FA1A S2_21_65 ( .A(\ab[21][65] ), .B(\CARRYB[20][65] ), .CI(\SUMB[20][66] ), 
        .CO(\CARRYB[21][65] ), .S(\SUMB[21][65] ) );
  FA1A S2_21_64 ( .A(\ab[21][64] ), .B(\CARRYB[20][64] ), .CI(\SUMB[20][65] ), 
        .CO(\CARRYB[21][64] ), .S(\SUMB[21][64] ) );
  FA1A S2_21_60 ( .A(\ab[21][60] ), .B(\CARRYB[20][60] ), .CI(\SUMB[20][61] ), 
        .CO(\CARRYB[21][60] ), .S(\SUMB[21][60] ) );
  FA1A S2_21_56 ( .A(\ab[21][56] ), .B(\CARRYB[20][56] ), .CI(\SUMB[20][57] ), 
        .CO(\CARRYB[21][56] ), .S(\SUMB[21][56] ) );
  FA1A S2_21_55 ( .A(\ab[21][55] ), .B(\CARRYB[20][55] ), .CI(\SUMB[20][56] ), 
        .CO(\CARRYB[21][55] ), .S(\SUMB[21][55] ) );
  FA1A S2_21_54 ( .A(\ab[21][54] ), .B(\CARRYB[20][54] ), .CI(\SUMB[20][55] ), 
        .CO(\CARRYB[21][54] ), .S(\SUMB[21][54] ) );
  FA1A S2_21_53 ( .A(\ab[21][53] ), .B(\CARRYB[20][53] ), .CI(\SUMB[20][54] ), 
        .CO(\CARRYB[21][53] ), .S(\SUMB[21][53] ) );
  FA1A S2_21_58 ( .A(\ab[21][58] ), .B(\CARRYB[20][58] ), .CI(\SUMB[20][59] ), 
        .CO(\CARRYB[21][58] ), .S(\SUMB[21][58] ) );
  FA1A S2_20_68 ( .A(\ab[20][68] ), .B(\CARRYB[19][68] ), .CI(\SUMB[19][69] ), 
        .CO(\CARRYB[20][68] ), .S(\SUMB[20][68] ) );
  FA1A S2_20_67 ( .A(\ab[20][67] ), .B(\CARRYB[19][67] ), .CI(\SUMB[19][68] ), 
        .CO(\CARRYB[20][67] ), .S(\SUMB[20][67] ) );
  FA1A S2_20_66 ( .A(\ab[20][66] ), .B(\CARRYB[19][66] ), .CI(\SUMB[19][67] ), 
        .CO(\CARRYB[20][66] ), .S(\SUMB[20][66] ) );
  FA1A S2_20_65 ( .A(\ab[20][65] ), .B(\CARRYB[19][65] ), .CI(\SUMB[19][66] ), 
        .CO(\CARRYB[20][65] ), .S(\SUMB[20][65] ) );
  FA1A S2_20_64 ( .A(\ab[20][64] ), .B(\CARRYB[19][64] ), .CI(\SUMB[19][65] ), 
        .CO(\CARRYB[20][64] ), .S(\SUMB[20][64] ) );
  FA1A S2_20_60 ( .A(\ab[20][60] ), .B(\CARRYB[19][60] ), .CI(\SUMB[19][61] ), 
        .CO(\CARRYB[20][60] ), .S(\SUMB[20][60] ) );
  FA1A S2_20_56 ( .A(\ab[20][56] ), .B(\CARRYB[19][56] ), .CI(\SUMB[19][57] ), 
        .CO(\CARRYB[20][56] ), .S(\SUMB[20][56] ) );
  FA1A S2_20_55 ( .A(\ab[20][55] ), .B(\CARRYB[19][55] ), .CI(\SUMB[19][56] ), 
        .CO(\CARRYB[20][55] ), .S(\SUMB[20][55] ) );
  FA1A S2_20_54 ( .A(\ab[20][54] ), .B(\CARRYB[19][54] ), .CI(\SUMB[19][55] ), 
        .CO(\CARRYB[20][54] ), .S(\SUMB[20][54] ) );
  FA1A S2_20_53 ( .A(\ab[20][53] ), .B(\CARRYB[19][53] ), .CI(\SUMB[19][54] ), 
        .CO(\CARRYB[20][53] ), .S(\SUMB[20][53] ) );
  FA1A S2_20_58 ( .A(\ab[20][58] ), .B(\CARRYB[19][58] ), .CI(\SUMB[19][59] ), 
        .CO(\CARRYB[20][58] ), .S(\SUMB[20][58] ) );
  FA1A S2_20_59 ( .A(\ab[20][59] ), .B(\CARRYB[19][59] ), .CI(\SUMB[19][60] ), 
        .CO(\CARRYB[20][59] ), .S(\SUMB[20][59] ) );
  FA1A S2_19_68 ( .A(\ab[19][68] ), .B(\CARRYB[18][68] ), .CI(\SUMB[18][69] ), 
        .CO(\CARRYB[19][68] ), .S(\SUMB[19][68] ) );
  FA1A S2_19_67 ( .A(\ab[19][67] ), .B(\CARRYB[18][67] ), .CI(\SUMB[18][68] ), 
        .CO(\CARRYB[19][67] ), .S(\SUMB[19][67] ) );
  FA1A S2_19_66 ( .A(\ab[19][66] ), .B(\CARRYB[18][66] ), .CI(\SUMB[18][67] ), 
        .CO(\CARRYB[19][66] ), .S(\SUMB[19][66] ) );
  FA1A S2_19_65 ( .A(\ab[19][65] ), .B(\CARRYB[18][65] ), .CI(\SUMB[18][66] ), 
        .CO(\CARRYB[19][65] ), .S(\SUMB[19][65] ) );
  FA1A S2_19_64 ( .A(\ab[19][64] ), .B(\CARRYB[18][64] ), .CI(\SUMB[18][65] ), 
        .CO(\CARRYB[19][64] ), .S(\SUMB[19][64] ) );
  FA1A S2_19_60 ( .A(\ab[19][60] ), .B(\CARRYB[18][60] ), .CI(\SUMB[18][61] ), 
        .CO(\CARRYB[19][60] ), .S(\SUMB[19][60] ) );
  FA1A S2_19_58 ( .A(\ab[19][58] ), .B(\CARRYB[18][58] ), .CI(\SUMB[18][59] ), 
        .CO(\CARRYB[19][58] ), .S(\SUMB[19][58] ) );
  FA1A S2_19_56 ( .A(\ab[19][56] ), .B(\CARRYB[18][56] ), .CI(\SUMB[18][57] ), 
        .CO(\CARRYB[19][56] ), .S(\SUMB[19][56] ) );
  FA1A S2_19_55 ( .A(\ab[19][55] ), .B(\CARRYB[18][55] ), .CI(\SUMB[18][56] ), 
        .CO(\CARRYB[19][55] ), .S(\SUMB[19][55] ) );
  FA1A S2_19_54 ( .A(\ab[19][54] ), .B(\CARRYB[18][54] ), .CI(\SUMB[18][55] ), 
        .CO(\CARRYB[19][54] ), .S(\SUMB[19][54] ) );
  FA1A S2_19_53 ( .A(\ab[19][53] ), .B(\CARRYB[18][53] ), .CI(\SUMB[18][54] ), 
        .CO(\CARRYB[19][53] ), .S(\SUMB[19][53] ) );
  FA1A S2_19_59 ( .A(\ab[19][59] ), .B(\CARRYB[18][59] ), .CI(\SUMB[18][60] ), 
        .CO(\CARRYB[19][59] ), .S(\SUMB[19][59] ) );
  FA1A S2_18_68 ( .A(\ab[18][68] ), .B(\CARRYB[17][68] ), .CI(\SUMB[17][69] ), 
        .CO(\CARRYB[18][68] ), .S(\SUMB[18][68] ) );
  FA1A S2_18_67 ( .A(\ab[18][67] ), .B(\CARRYB[17][67] ), .CI(\SUMB[17][68] ), 
        .CO(\CARRYB[18][67] ), .S(\SUMB[18][67] ) );
  FA1A S2_18_66 ( .A(\ab[18][66] ), .B(\CARRYB[17][66] ), .CI(\SUMB[17][67] ), 
        .CO(\CARRYB[18][66] ), .S(\SUMB[18][66] ) );
  FA1A S2_18_65 ( .A(\ab[18][65] ), .B(\CARRYB[17][65] ), .CI(\SUMB[17][66] ), 
        .CO(\CARRYB[18][65] ), .S(\SUMB[18][65] ) );
  FA1A S2_18_64 ( .A(\ab[18][64] ), .B(\CARRYB[17][64] ), .CI(\SUMB[17][65] ), 
        .CO(\CARRYB[18][64] ), .S(\SUMB[18][64] ) );
  FA1A S2_18_60 ( .A(\ab[18][60] ), .B(\CARRYB[17][60] ), .CI(\SUMB[17][61] ), 
        .CO(\CARRYB[18][60] ), .S(\SUMB[18][60] ) );
  FA1A S2_18_53 ( .A(\ab[18][53] ), .B(\CARRYB[17][53] ), .CI(\SUMB[17][54] ), 
        .CO(\CARRYB[18][53] ), .S(\SUMB[18][53] ) );
  FA1A S2_18_59 ( .A(\ab[18][59] ), .B(\CARRYB[17][59] ), .CI(\SUMB[17][60] ), 
        .CO(\CARRYB[18][59] ), .S(\SUMB[18][59] ) );
  FA1A S2_18_58 ( .A(\ab[18][58] ), .B(\CARRYB[17][58] ), .CI(\SUMB[17][59] ), 
        .CO(\CARRYB[18][58] ), .S(\SUMB[18][58] ) );
  FA1A S2_18_56 ( .A(\ab[18][56] ), .B(\CARRYB[17][56] ), .CI(\SUMB[17][57] ), 
        .CO(\CARRYB[18][56] ), .S(\SUMB[18][56] ) );
  FA1A S2_18_55 ( .A(\ab[18][55] ), .B(\CARRYB[17][55] ), .CI(\SUMB[17][56] ), 
        .CO(\CARRYB[18][55] ), .S(\SUMB[18][55] ) );
  FA1A S2_18_54 ( .A(\ab[18][54] ), .B(\CARRYB[17][54] ), .CI(\SUMB[17][55] ), 
        .CO(\CARRYB[18][54] ), .S(\SUMB[18][54] ) );
  FA1A S2_17_68 ( .A(\ab[17][68] ), .B(\CARRYB[16][68] ), .CI(\SUMB[16][69] ), 
        .CO(\CARRYB[17][68] ), .S(\SUMB[17][68] ) );
  FA1A S2_17_67 ( .A(\ab[17][67] ), .B(\CARRYB[16][67] ), .CI(\SUMB[16][68] ), 
        .CO(\CARRYB[17][67] ), .S(\SUMB[17][67] ) );
  FA1A S2_17_66 ( .A(\ab[17][66] ), .B(\CARRYB[16][66] ), .CI(\SUMB[16][67] ), 
        .CO(\CARRYB[17][66] ), .S(\SUMB[17][66] ) );
  FA1A S2_17_65 ( .A(\ab[17][65] ), .B(\CARRYB[16][65] ), .CI(\SUMB[16][66] ), 
        .CO(\CARRYB[17][65] ), .S(\SUMB[17][65] ) );
  FA1A S2_17_64 ( .A(\ab[17][64] ), .B(\CARRYB[16][64] ), .CI(\SUMB[16][65] ), 
        .CO(\CARRYB[17][64] ), .S(\SUMB[17][64] ) );
  FA1A S2_17_60 ( .A(\ab[17][60] ), .B(\CARRYB[16][60] ), .CI(\SUMB[16][61] ), 
        .CO(\CARRYB[17][60] ), .S(\SUMB[17][60] ) );
  FA1A S2_17_54 ( .A(\ab[17][54] ), .B(\CARRYB[16][54] ), .CI(\SUMB[16][55] ), 
        .CO(\CARRYB[17][54] ), .S(\SUMB[17][54] ) );
  FA1A S2_17_53 ( .A(\ab[17][53] ), .B(\CARRYB[16][53] ), .CI(\SUMB[16][54] ), 
        .CO(\CARRYB[17][53] ), .S(\SUMB[17][53] ) );
  FA1A S2_17_59 ( .A(\ab[17][59] ), .B(\CARRYB[16][59] ), .CI(\SUMB[16][60] ), 
        .CO(\CARRYB[17][59] ), .S(\SUMB[17][59] ) );
  FA1A S2_17_58 ( .A(\ab[17][58] ), .B(\CARRYB[16][58] ), .CI(\SUMB[16][59] ), 
        .CO(\CARRYB[17][58] ), .S(\SUMB[17][58] ) );
  FA1A S2_17_56 ( .A(\ab[17][56] ), .B(\CARRYB[16][56] ), .CI(\SUMB[16][57] ), 
        .CO(\CARRYB[17][56] ), .S(\SUMB[17][56] ) );
  FA1A S2_17_55 ( .A(\ab[17][55] ), .B(\CARRYB[16][55] ), .CI(\SUMB[16][56] ), 
        .CO(\CARRYB[17][55] ), .S(\SUMB[17][55] ) );
  FA1A S2_16_68 ( .A(\ab[16][68] ), .B(\CARRYB[15][68] ), .CI(\SUMB[15][69] ), 
        .CO(\CARRYB[16][68] ), .S(\SUMB[16][68] ) );
  FA1A S2_16_67 ( .A(\ab[16][67] ), .B(\CARRYB[15][67] ), .CI(\SUMB[15][68] ), 
        .CO(\CARRYB[16][67] ), .S(\SUMB[16][67] ) );
  FA1A S2_16_66 ( .A(\ab[16][66] ), .B(\CARRYB[15][66] ), .CI(\SUMB[15][67] ), 
        .CO(\CARRYB[16][66] ), .S(\SUMB[16][66] ) );
  FA1A S2_16_65 ( .A(\ab[16][65] ), .B(\CARRYB[15][65] ), .CI(\SUMB[15][66] ), 
        .CO(\CARRYB[16][65] ), .S(\SUMB[16][65] ) );
  FA1A S2_16_64 ( .A(\ab[16][64] ), .B(\CARRYB[15][64] ), .CI(\SUMB[15][65] ), 
        .CO(\CARRYB[16][64] ), .S(\SUMB[16][64] ) );
  FA1A S2_16_60 ( .A(\ab[16][60] ), .B(\CARRYB[15][60] ), .CI(\SUMB[15][61] ), 
        .CO(\CARRYB[16][60] ), .S(\SUMB[16][60] ) );
  FA1A S2_16_55 ( .A(\ab[16][55] ), .B(\CARRYB[15][55] ), .CI(\SUMB[15][56] ), 
        .CO(\CARRYB[16][55] ), .S(\SUMB[16][55] ) );
  FA1A S2_16_54 ( .A(\ab[16][54] ), .B(\CARRYB[15][54] ), .CI(\SUMB[15][55] ), 
        .CO(\CARRYB[16][54] ), .S(\SUMB[16][54] ) );
  FA1A S2_16_53 ( .A(\ab[16][53] ), .B(\CARRYB[15][53] ), .CI(\SUMB[15][54] ), 
        .CO(\CARRYB[16][53] ), .S(\SUMB[16][53] ) );
  FA1A S2_16_59 ( .A(\ab[16][59] ), .B(\CARRYB[15][59] ), .CI(\SUMB[15][60] ), 
        .CO(\CARRYB[16][59] ), .S(\SUMB[16][59] ) );
  FA1A S2_16_58 ( .A(\ab[16][58] ), .B(\CARRYB[15][58] ), .CI(\SUMB[15][59] ), 
        .CO(\CARRYB[16][58] ), .S(\SUMB[16][58] ) );
  FA1A S2_16_56 ( .A(\ab[16][56] ), .B(\CARRYB[15][56] ), .CI(\SUMB[15][57] ), 
        .CO(\CARRYB[16][56] ), .S(\SUMB[16][56] ) );
  FA1A S2_15_68 ( .A(\ab[15][68] ), .B(\CARRYB[14][68] ), .CI(\SUMB[14][69] ), 
        .CO(\CARRYB[15][68] ), .S(\SUMB[15][68] ) );
  FA1A S2_15_67 ( .A(\ab[15][67] ), .B(\CARRYB[14][67] ), .CI(\SUMB[14][68] ), 
        .CO(\CARRYB[15][67] ), .S(\SUMB[15][67] ) );
  FA1A S2_15_66 ( .A(\ab[15][66] ), .B(\CARRYB[14][66] ), .CI(\SUMB[14][67] ), 
        .CO(\CARRYB[15][66] ), .S(\SUMB[15][66] ) );
  FA1A S2_15_65 ( .A(\ab[15][65] ), .B(\CARRYB[14][65] ), .CI(\SUMB[14][66] ), 
        .CO(\CARRYB[15][65] ), .S(\SUMB[15][65] ) );
  FA1A S2_15_64 ( .A(\ab[15][64] ), .B(\CARRYB[14][64] ), .CI(\SUMB[14][65] ), 
        .CO(\CARRYB[15][64] ), .S(\SUMB[15][64] ) );
  FA1A S2_15_60 ( .A(\ab[15][60] ), .B(\CARRYB[14][60] ), .CI(\SUMB[14][61] ), 
        .CO(\CARRYB[15][60] ), .S(\SUMB[15][60] ) );
  FA1A S2_15_56 ( .A(\ab[15][56] ), .B(\CARRYB[14][56] ), .CI(\SUMB[14][57] ), 
        .CO(\CARRYB[15][56] ), .S(\SUMB[15][56] ) );
  FA1A S2_15_55 ( .A(\ab[15][55] ), .B(\CARRYB[14][55] ), .CI(\SUMB[14][56] ), 
        .CO(\CARRYB[15][55] ), .S(\SUMB[15][55] ) );
  FA1A S2_15_54 ( .A(\ab[15][54] ), .B(\CARRYB[14][54] ), .CI(\SUMB[14][55] ), 
        .CO(\CARRYB[15][54] ), .S(\SUMB[15][54] ) );
  FA1A S2_15_53 ( .A(\ab[15][53] ), .B(\CARRYB[14][53] ), .CI(\SUMB[14][54] ), 
        .CO(\CARRYB[15][53] ), .S(\SUMB[15][53] ) );
  FA1A S2_15_59 ( .A(\ab[15][59] ), .B(\CARRYB[14][59] ), .CI(\SUMB[14][60] ), 
        .CO(\CARRYB[15][59] ), .S(\SUMB[15][59] ) );
  FA1A S2_15_58 ( .A(\ab[15][58] ), .B(\CARRYB[14][58] ), .CI(\SUMB[14][59] ), 
        .CO(\CARRYB[15][58] ), .S(\SUMB[15][58] ) );
  FA1A S2_14_55 ( .A(\ab[14][55] ), .B(\CARRYB[13][55] ), .CI(\SUMB[13][56] ), 
        .CO(\CARRYB[14][55] ), .S(\SUMB[14][55] ) );
  FA1A S2_13_55 ( .A(\ab[13][55] ), .B(\CARRYB[12][55] ), .CI(\SUMB[12][56] ), 
        .CO(\CARRYB[13][55] ), .S(\SUMB[13][55] ) );
  FA1A S2_12_55 ( .A(\ab[12][55] ), .B(\CARRYB[11][55] ), .CI(\SUMB[11][56] ), 
        .CO(\CARRYB[12][55] ), .S(\SUMB[12][55] ) );
  FA1A S2_11_55 ( .A(\ab[11][55] ), .B(\CARRYB[10][55] ), .CI(\SUMB[10][56] ), 
        .CO(\CARRYB[11][55] ), .S(\SUMB[11][55] ) );
  FA1A S2_10_55 ( .A(\ab[10][55] ), .B(\CARRYB[9][55] ), .CI(\SUMB[9][56] ), 
        .CO(\CARRYB[10][55] ), .S(\SUMB[10][55] ) );
  FA1A S2_9_55 ( .A(\ab[9][55] ), .B(\CARRYB[8][55] ), .CI(\SUMB[8][56] ), 
        .CO(\CARRYB[9][55] ), .S(\SUMB[9][55] ) );
  FA1A S2_8_55 ( .A(\ab[8][55] ), .B(\CARRYB[7][55] ), .CI(\SUMB[7][56] ), 
        .CO(\CARRYB[8][55] ), .S(\SUMB[8][55] ) );
  FA1A S2_7_55 ( .A(\ab[7][55] ), .B(\CARRYB[6][55] ), .CI(\SUMB[6][56] ), 
        .CO(\CARRYB[7][55] ), .S(\SUMB[7][55] ) );
  FA1A S2_6_55 ( .A(\ab[6][55] ), .B(\CARRYB[5][55] ), .CI(\SUMB[5][56] ), 
        .CO(\CARRYB[6][55] ), .S(\SUMB[6][55] ) );
  FA1A S2_5_55 ( .A(\ab[5][55] ), .B(\CARRYB[4][55] ), .CI(\SUMB[4][56] ), 
        .CO(\CARRYB[5][55] ), .S(\SUMB[5][55] ) );
  FA1A S2_4_55 ( .A(\ab[4][55] ), .B(\CARRYB[3][55] ), .CI(\SUMB[3][56] ), 
        .CO(\CARRYB[4][55] ), .S(\SUMB[4][55] ) );
  FA1A S2_3_55 ( .A(\ab[3][55] ), .B(\CARRYB[2][55] ), .CI(\SUMB[2][56] ), 
        .CO(\CARRYB[3][55] ), .S(\SUMB[3][55] ) );
  FA1A S2_2_55 ( .A(\ab[2][55] ), .B(\CARRYB[1][55] ), .CI(\SUMB[1][56] ), 
        .CO(\CARRYB[2][55] ), .S(\SUMB[2][55] ) );
  FA1A S4_68 ( .A(\ab[29][68] ), .B(\CARRYB[28][68] ), .CI(\SUMB[28][69] ), 
        .CO(\CARRYB[29][68] ), .S(\SUMB[29][68] ) );
  FA1A S4_56 ( .A(\ab[29][56] ), .B(\CARRYB[28][56] ), .CI(\SUMB[28][57] ), 
        .CO(\CARRYB[29][56] ), .S(\SUMB[29][56] ) );
  FA1A S4_55 ( .A(\ab[29][55] ), .B(\CARRYB[28][55] ), .CI(\SUMB[28][56] ), 
        .CO(\CARRYB[29][55] ), .S(\SUMB[29][55] ) );
  FA1A S4_59 ( .A(\ab[29][59] ), .B(\CARRYB[28][59] ), .CI(\SUMB[28][60] ), 
        .CO(\CARRYB[29][59] ), .S(\SUMB[29][59] ) );
  FA1A S4_39 ( .A(\ab[29][39] ), .B(\CARRYB[28][39] ), .CI(\SUMB[28][40] ), 
        .CO(\CARRYB[29][39] ), .S(\SUMB[29][39] ) );
  FA1A S4_44 ( .A(\ab[29][44] ), .B(\CARRYB[28][44] ), .CI(\SUMB[28][45] ), 
        .CO(\CARRYB[29][44] ), .S(\SUMB[29][44] ) );
  FA1A S4_43 ( .A(\ab[29][43] ), .B(\CARRYB[28][43] ), .CI(\SUMB[28][44] ), 
        .CO(\CARRYB[29][43] ), .S(\SUMB[29][43] ) );
  FA1A S2_28_52 ( .A(\ab[28][52] ), .B(\CARRYB[27][52] ), .CI(\SUMB[27][53] ), 
        .CO(\CARRYB[28][52] ), .S(\SUMB[28][52] ) );
  FA1A S2_28_44 ( .A(\ab[28][44] ), .B(\CARRYB[27][44] ), .CI(\SUMB[27][45] ), 
        .CO(\CARRYB[28][44] ), .S(\SUMB[28][44] ) );
  FA1A S4_61 ( .A(\ab[29][61] ), .B(\CARRYB[28][61] ), .CI(\SUMB[28][62] ), 
        .CO(\CARRYB[29][61] ), .S(\SUMB[29][61] ) );
  FA1A S4_62 ( .A(\ab[29][62] ), .B(\CARRYB[28][62] ), .CI(\SUMB[28][63] ), 
        .CO(\CARRYB[29][62] ), .S(\SUMB[29][62] ) );
  FA1A S4_42 ( .A(\ab[29][42] ), .B(\CARRYB[28][42] ), .CI(\SUMB[28][43] ), 
        .CO(\CARRYB[29][42] ), .S(\SUMB[29][42] ) );
  FA1A S4_41 ( .A(\ab[29][41] ), .B(\CARRYB[28][41] ), .CI(\SUMB[28][42] ), 
        .CO(\CARRYB[29][41] ), .S(\SUMB[29][41] ) );
  FA1A S4_40 ( .A(\ab[29][40] ), .B(\CARRYB[28][40] ), .CI(\SUMB[28][41] ), 
        .CO(\CARRYB[29][40] ), .S(\SUMB[29][40] ) );
  FA1A S2_28_61 ( .A(\ab[28][61] ), .B(\CARRYB[27][61] ), .CI(\SUMB[27][62] ), 
        .CO(\CARRYB[28][61] ), .S(\SUMB[28][61] ) );
  FA1A S2_28_62 ( .A(\ab[28][62] ), .B(\CARRYB[27][62] ), .CI(\SUMB[27][63] ), 
        .CO(\CARRYB[28][62] ), .S(\SUMB[28][62] ) );
  FA1A S2_28_63 ( .A(\ab[28][63] ), .B(\CARRYB[27][63] ), .CI(\SUMB[27][64] ), 
        .CO(\CARRYB[28][63] ), .S(\SUMB[28][63] ) );
  FA1A S2_28_43 ( .A(\ab[28][43] ), .B(\CARRYB[27][43] ), .CI(\SUMB[27][44] ), 
        .CO(\CARRYB[28][43] ), .S(\SUMB[28][43] ) );
  FA1A S2_28_42 ( .A(\ab[28][42] ), .B(\CARRYB[27][42] ), .CI(\SUMB[27][43] ), 
        .CO(\CARRYB[28][42] ), .S(\SUMB[28][42] ) );
  FA1A S2_28_41 ( .A(\ab[28][41] ), .B(\CARRYB[27][41] ), .CI(\SUMB[27][42] ), 
        .CO(\CARRYB[28][41] ), .S(\SUMB[28][41] ) );
  FA1A S2_28_40 ( .A(\ab[28][40] ), .B(\CARRYB[27][40] ), .CI(\SUMB[27][41] ), 
        .CO(\CARRYB[28][40] ), .S(\SUMB[28][40] ) );
  FA1A S2_28_39 ( .A(\ab[28][39] ), .B(\CARRYB[27][39] ), .CI(\SUMB[27][40] ), 
        .CO(\CARRYB[28][39] ), .S(\SUMB[28][39] ) );
  FA1A S2_27_62 ( .A(\ab[27][62] ), .B(\CARRYB[26][62] ), .CI(\SUMB[26][63] ), 
        .CO(\CARRYB[27][62] ), .S(\SUMB[27][62] ) );
  FA1A S2_27_61 ( .A(\ab[27][61] ), .B(\CARRYB[26][61] ), .CI(\SUMB[26][62] ), 
        .CO(\CARRYB[27][61] ), .S(\SUMB[27][61] ) );
  FA1A S2_27_63 ( .A(\ab[27][63] ), .B(\CARRYB[26][63] ), .CI(\SUMB[26][64] ), 
        .CO(\CARRYB[27][63] ), .S(\SUMB[27][63] ) );
  FA1A S2_27_44 ( .A(\ab[27][44] ), .B(\CARRYB[26][44] ), .CI(\SUMB[26][45] ), 
        .CO(\CARRYB[27][44] ), .S(\SUMB[27][44] ) );
  FA1A S2_27_43 ( .A(\ab[27][43] ), .B(\CARRYB[26][43] ), .CI(\SUMB[26][44] ), 
        .CO(\CARRYB[27][43] ), .S(\SUMB[27][43] ) );
  FA1A S2_27_42 ( .A(\ab[27][42] ), .B(\CARRYB[26][42] ), .CI(\SUMB[26][43] ), 
        .CO(\CARRYB[27][42] ), .S(\SUMB[27][42] ) );
  FA1A S2_27_41 ( .A(\ab[27][41] ), .B(\CARRYB[26][41] ), .CI(\SUMB[26][42] ), 
        .CO(\CARRYB[27][41] ), .S(\SUMB[27][41] ) );
  FA1A S2_27_40 ( .A(\ab[27][40] ), .B(\CARRYB[26][40] ), .CI(\SUMB[26][41] ), 
        .CO(\CARRYB[27][40] ), .S(\SUMB[27][40] ) );
  FA1A S2_27_39 ( .A(\ab[27][39] ), .B(\CARRYB[26][39] ), .CI(\SUMB[26][40] ), 
        .CO(\CARRYB[27][39] ), .S(\SUMB[27][39] ) );
  FA1A S2_27_52 ( .A(\ab[27][52] ), .B(\CARRYB[26][52] ), .CI(\SUMB[26][53] ), 
        .CO(\CARRYB[27][52] ), .S(\SUMB[27][52] ) );
  FA1A S2_26_63 ( .A(\ab[26][63] ), .B(\CARRYB[25][63] ), .CI(\SUMB[25][64] ), 
        .CO(\CARRYB[26][63] ), .S(\SUMB[26][63] ) );
  FA1A S2_26_62 ( .A(\ab[26][62] ), .B(\CARRYB[25][62] ), .CI(\SUMB[25][63] ), 
        .CO(\CARRYB[26][62] ), .S(\SUMB[26][62] ) );
  FA1A S2_26_61 ( .A(\ab[26][61] ), .B(\CARRYB[25][61] ), .CI(\SUMB[25][62] ), 
        .CO(\CARRYB[26][61] ), .S(\SUMB[26][61] ) );
  FA1A S2_26_44 ( .A(\ab[26][44] ), .B(\CARRYB[25][44] ), .CI(\SUMB[25][45] ), 
        .CO(\CARRYB[26][44] ), .S(\SUMB[26][44] ) );
  FA1A S2_26_43 ( .A(\ab[26][43] ), .B(\CARRYB[25][43] ), .CI(\SUMB[25][44] ), 
        .CO(\CARRYB[26][43] ), .S(\SUMB[26][43] ) );
  FA1A S2_26_42 ( .A(\ab[26][42] ), .B(\CARRYB[25][42] ), .CI(\SUMB[25][43] ), 
        .CO(\CARRYB[26][42] ), .S(\SUMB[26][42] ) );
  FA1A S2_26_41 ( .A(\ab[26][41] ), .B(\CARRYB[25][41] ), .CI(\SUMB[25][42] ), 
        .CO(\CARRYB[26][41] ), .S(\SUMB[26][41] ) );
  FA1A S2_26_40 ( .A(\ab[26][40] ), .B(\CARRYB[25][40] ), .CI(\SUMB[25][41] ), 
        .CO(\CARRYB[26][40] ), .S(\SUMB[26][40] ) );
  FA1A S2_26_39 ( .A(\ab[26][39] ), .B(\CARRYB[25][39] ), .CI(\SUMB[25][40] ), 
        .CO(\CARRYB[26][39] ), .S(\SUMB[26][39] ) );
  FA1A S2_26_52 ( .A(\ab[26][52] ), .B(\CARRYB[25][52] ), .CI(\SUMB[25][53] ), 
        .CO(\CARRYB[26][52] ), .S(\SUMB[26][52] ) );
  FA1A S2_25_63 ( .A(\ab[25][63] ), .B(\CARRYB[24][63] ), .CI(\SUMB[24][64] ), 
        .CO(\CARRYB[25][63] ), .S(\SUMB[25][63] ) );
  FA1A S2_25_62 ( .A(\ab[25][62] ), .B(\CARRYB[24][62] ), .CI(\SUMB[24][63] ), 
        .CO(\CARRYB[25][62] ), .S(\SUMB[25][62] ) );
  FA1A S2_25_61 ( .A(\ab[25][61] ), .B(\CARRYB[24][61] ), .CI(\SUMB[24][62] ), 
        .CO(\CARRYB[25][61] ), .S(\SUMB[25][61] ) );
  FA1A S2_25_44 ( .A(\ab[25][44] ), .B(\CARRYB[24][44] ), .CI(\SUMB[24][45] ), 
        .CO(\CARRYB[25][44] ), .S(\SUMB[25][44] ) );
  FA1A S2_25_43 ( .A(\ab[25][43] ), .B(\CARRYB[24][43] ), .CI(\SUMB[24][44] ), 
        .CO(\CARRYB[25][43] ), .S(\SUMB[25][43] ) );
  FA1A S2_25_42 ( .A(\ab[25][42] ), .B(\CARRYB[24][42] ), .CI(\SUMB[24][43] ), 
        .CO(\CARRYB[25][42] ), .S(\SUMB[25][42] ) );
  FA1A S2_25_41 ( .A(\ab[25][41] ), .B(\CARRYB[24][41] ), .CI(\SUMB[24][42] ), 
        .CO(\CARRYB[25][41] ), .S(\SUMB[25][41] ) );
  FA1A S2_25_40 ( .A(\ab[25][40] ), .B(\CARRYB[24][40] ), .CI(\SUMB[24][41] ), 
        .CO(\CARRYB[25][40] ), .S(\SUMB[25][40] ) );
  FA1A S2_25_39 ( .A(\ab[25][39] ), .B(\CARRYB[24][39] ), .CI(\SUMB[24][40] ), 
        .CO(\CARRYB[25][39] ), .S(\SUMB[25][39] ) );
  FA1A S2_25_52 ( .A(\ab[25][52] ), .B(\CARRYB[24][52] ), .CI(\SUMB[24][53] ), 
        .CO(\CARRYB[25][52] ), .S(\SUMB[25][52] ) );
  FA1A S2_24_63 ( .A(\ab[24][63] ), .B(\CARRYB[23][63] ), .CI(\SUMB[23][64] ), 
        .CO(\CARRYB[24][63] ), .S(\SUMB[24][63] ) );
  FA1A S2_24_62 ( .A(\ab[24][62] ), .B(\CARRYB[23][62] ), .CI(\SUMB[23][63] ), 
        .CO(\CARRYB[24][62] ), .S(\SUMB[24][62] ) );
  FA1A S2_24_61 ( .A(\ab[24][61] ), .B(\CARRYB[23][61] ), .CI(\SUMB[23][62] ), 
        .CO(\CARRYB[24][61] ), .S(\SUMB[24][61] ) );
  FA1A S2_24_44 ( .A(\ab[24][44] ), .B(\CARRYB[23][44] ), .CI(\SUMB[23][45] ), 
        .CO(\CARRYB[24][44] ), .S(\SUMB[24][44] ) );
  FA1A S2_24_43 ( .A(\ab[24][43] ), .B(\CARRYB[23][43] ), .CI(\SUMB[23][44] ), 
        .CO(\CARRYB[24][43] ), .S(\SUMB[24][43] ) );
  FA1A S2_24_42 ( .A(\ab[24][42] ), .B(\CARRYB[23][42] ), .CI(\SUMB[23][43] ), 
        .CO(\CARRYB[24][42] ), .S(\SUMB[24][42] ) );
  FA1A S2_24_41 ( .A(\ab[24][41] ), .B(\CARRYB[23][41] ), .CI(\SUMB[23][42] ), 
        .CO(\CARRYB[24][41] ), .S(\SUMB[24][41] ) );
  FA1A S2_24_40 ( .A(\ab[24][40] ), .B(\CARRYB[23][40] ), .CI(\SUMB[23][41] ), 
        .CO(\CARRYB[24][40] ), .S(\SUMB[24][40] ) );
  FA1A S2_24_39 ( .A(\ab[24][39] ), .B(\CARRYB[23][39] ), .CI(\SUMB[23][40] ), 
        .CO(\CARRYB[24][39] ), .S(\SUMB[24][39] ) );
  FA1A S2_24_52 ( .A(\ab[24][52] ), .B(\CARRYB[23][52] ), .CI(\SUMB[23][53] ), 
        .CO(\CARRYB[24][52] ), .S(\SUMB[24][52] ) );
  FA1A S2_23_63 ( .A(\ab[23][63] ), .B(\CARRYB[22][63] ), .CI(\SUMB[22][64] ), 
        .CO(\CARRYB[23][63] ), .S(\SUMB[23][63] ) );
  FA1A S2_23_62 ( .A(\ab[23][62] ), .B(\CARRYB[22][62] ), .CI(\SUMB[22][63] ), 
        .CO(\CARRYB[23][62] ), .S(\SUMB[23][62] ) );
  FA1A S2_23_61 ( .A(\ab[23][61] ), .B(\CARRYB[22][61] ), .CI(\SUMB[22][62] ), 
        .CO(\CARRYB[23][61] ), .S(\SUMB[23][61] ) );
  FA1A S2_23_44 ( .A(\ab[23][44] ), .B(\CARRYB[22][44] ), .CI(\SUMB[22][45] ), 
        .CO(\CARRYB[23][44] ), .S(\SUMB[23][44] ) );
  FA1A S2_23_43 ( .A(\ab[23][43] ), .B(\CARRYB[22][43] ), .CI(\SUMB[22][44] ), 
        .CO(\CARRYB[23][43] ), .S(\SUMB[23][43] ) );
  FA1A S2_23_42 ( .A(\ab[23][42] ), .B(\CARRYB[22][42] ), .CI(\SUMB[22][43] ), 
        .CO(\CARRYB[23][42] ), .S(\SUMB[23][42] ) );
  FA1A S2_23_41 ( .A(\ab[23][41] ), .B(\CARRYB[22][41] ), .CI(\SUMB[22][42] ), 
        .CO(\CARRYB[23][41] ), .S(\SUMB[23][41] ) );
  FA1A S2_23_40 ( .A(\ab[23][40] ), .B(\CARRYB[22][40] ), .CI(\SUMB[22][41] ), 
        .CO(\CARRYB[23][40] ), .S(\SUMB[23][40] ) );
  FA1A S2_23_39 ( .A(\ab[23][39] ), .B(\CARRYB[22][39] ), .CI(\SUMB[22][40] ), 
        .CO(\CARRYB[23][39] ), .S(\SUMB[23][39] ) );
  FA1A S2_23_52 ( .A(\ab[23][52] ), .B(\CARRYB[22][52] ), .CI(\SUMB[22][53] ), 
        .CO(\CARRYB[23][52] ), .S(\SUMB[23][52] ) );
  FA1A S2_22_63 ( .A(\ab[22][63] ), .B(\CARRYB[21][63] ), .CI(\SUMB[21][64] ), 
        .CO(\CARRYB[22][63] ), .S(\SUMB[22][63] ) );
  FA1A S2_22_62 ( .A(\ab[22][62] ), .B(\CARRYB[21][62] ), .CI(\SUMB[21][63] ), 
        .CO(\CARRYB[22][62] ), .S(\SUMB[22][62] ) );
  FA1A S2_22_61 ( .A(\ab[22][61] ), .B(\CARRYB[21][61] ), .CI(\SUMB[21][62] ), 
        .CO(\CARRYB[22][61] ), .S(\SUMB[22][61] ) );
  FA1A S2_22_44 ( .A(\ab[22][44] ), .B(\CARRYB[21][44] ), .CI(\SUMB[21][45] ), 
        .CO(\CARRYB[22][44] ), .S(\SUMB[22][44] ) );
  FA1A S2_22_43 ( .A(\ab[22][43] ), .B(\CARRYB[21][43] ), .CI(\SUMB[21][44] ), 
        .CO(\CARRYB[22][43] ), .S(\SUMB[22][43] ) );
  FA1A S2_22_42 ( .A(\ab[22][42] ), .B(\CARRYB[21][42] ), .CI(\SUMB[21][43] ), 
        .CO(\CARRYB[22][42] ), .S(\SUMB[22][42] ) );
  FA1A S2_22_41 ( .A(\ab[22][41] ), .B(\CARRYB[21][41] ), .CI(\SUMB[21][42] ), 
        .CO(\CARRYB[22][41] ), .S(\SUMB[22][41] ) );
  FA1A S2_22_40 ( .A(\ab[22][40] ), .B(\CARRYB[21][40] ), .CI(\SUMB[21][41] ), 
        .CO(\CARRYB[22][40] ), .S(\SUMB[22][40] ) );
  FA1A S2_22_39 ( .A(\ab[22][39] ), .B(\CARRYB[21][39] ), .CI(\SUMB[21][40] ), 
        .CO(\CARRYB[22][39] ), .S(\SUMB[22][39] ) );
  FA1A S2_22_52 ( .A(\ab[22][52] ), .B(\CARRYB[21][52] ), .CI(\SUMB[21][53] ), 
        .CO(\CARRYB[22][52] ), .S(\SUMB[22][52] ) );
  FA1A S2_21_63 ( .A(\ab[21][63] ), .B(\CARRYB[20][63] ), .CI(\SUMB[20][64] ), 
        .CO(\CARRYB[21][63] ), .S(\SUMB[21][63] ) );
  FA1A S2_21_62 ( .A(\ab[21][62] ), .B(\CARRYB[20][62] ), .CI(\SUMB[20][63] ), 
        .CO(\CARRYB[21][62] ), .S(\SUMB[21][62] ) );
  FA1A S2_21_61 ( .A(\ab[21][61] ), .B(\CARRYB[20][61] ), .CI(\SUMB[20][62] ), 
        .CO(\CARRYB[21][61] ), .S(\SUMB[21][61] ) );
  FA1A S2_21_44 ( .A(\ab[21][44] ), .B(\CARRYB[20][44] ), .CI(\SUMB[20][45] ), 
        .CO(\CARRYB[21][44] ), .S(\SUMB[21][44] ) );
  FA1A S2_21_43 ( .A(\ab[21][43] ), .B(\CARRYB[20][43] ), .CI(\SUMB[20][44] ), 
        .CO(\CARRYB[21][43] ), .S(\SUMB[21][43] ) );
  FA1A S2_21_42 ( .A(\ab[21][42] ), .B(\CARRYB[20][42] ), .CI(\SUMB[20][43] ), 
        .CO(\CARRYB[21][42] ), .S(\SUMB[21][42] ) );
  FA1A S2_21_41 ( .A(\ab[21][41] ), .B(\CARRYB[20][41] ), .CI(\SUMB[20][42] ), 
        .CO(\CARRYB[21][41] ), .S(\SUMB[21][41] ) );
  FA1A S2_21_40 ( .A(\ab[21][40] ), .B(\CARRYB[20][40] ), .CI(\SUMB[20][41] ), 
        .CO(\CARRYB[21][40] ), .S(\SUMB[21][40] ) );
  FA1A S2_21_39 ( .A(\ab[21][39] ), .B(\CARRYB[20][39] ), .CI(\SUMB[20][40] ), 
        .CO(\CARRYB[21][39] ), .S(\SUMB[21][39] ) );
  FA1A S2_21_52 ( .A(\ab[21][52] ), .B(\CARRYB[20][52] ), .CI(\SUMB[20][53] ), 
        .CO(\CARRYB[21][52] ), .S(\SUMB[21][52] ) );
  FA1A S2_20_63 ( .A(\ab[20][63] ), .B(\CARRYB[19][63] ), .CI(\SUMB[19][64] ), 
        .CO(\CARRYB[20][63] ), .S(\SUMB[20][63] ) );
  FA1A S2_20_62 ( .A(\ab[20][62] ), .B(\CARRYB[19][62] ), .CI(\SUMB[19][63] ), 
        .CO(\CARRYB[20][62] ), .S(\SUMB[20][62] ) );
  FA1A S2_20_61 ( .A(\ab[20][61] ), .B(\CARRYB[19][61] ), .CI(\SUMB[19][62] ), 
        .CO(\CARRYB[20][61] ), .S(\SUMB[20][61] ) );
  FA1A S2_20_44 ( .A(\ab[20][44] ), .B(\CARRYB[19][44] ), .CI(\SUMB[19][45] ), 
        .CO(\CARRYB[20][44] ), .S(\SUMB[20][44] ) );
  FA1A S2_20_43 ( .A(\ab[20][43] ), .B(\CARRYB[19][43] ), .CI(\SUMB[19][44] ), 
        .CO(\CARRYB[20][43] ), .S(\SUMB[20][43] ) );
  FA1A S2_20_42 ( .A(\ab[20][42] ), .B(\CARRYB[19][42] ), .CI(\SUMB[19][43] ), 
        .CO(\CARRYB[20][42] ), .S(\SUMB[20][42] ) );
  FA1A S2_20_41 ( .A(\ab[20][41] ), .B(\CARRYB[19][41] ), .CI(\SUMB[19][42] ), 
        .CO(\CARRYB[20][41] ), .S(\SUMB[20][41] ) );
  FA1A S2_20_40 ( .A(\ab[20][40] ), .B(\CARRYB[19][40] ), .CI(\SUMB[19][41] ), 
        .CO(\CARRYB[20][40] ), .S(\SUMB[20][40] ) );
  FA1A S2_20_39 ( .A(\ab[20][39] ), .B(\CARRYB[19][39] ), .CI(\SUMB[19][40] ), 
        .CO(\CARRYB[20][39] ), .S(\SUMB[20][39] ) );
  FA1A S2_20_52 ( .A(\ab[20][52] ), .B(\CARRYB[19][52] ), .CI(\SUMB[19][53] ), 
        .CO(\CARRYB[20][52] ), .S(\SUMB[20][52] ) );
  FA1A S2_19_63 ( .A(\ab[19][63] ), .B(\CARRYB[18][63] ), .CI(\SUMB[18][64] ), 
        .CO(\CARRYB[19][63] ), .S(\SUMB[19][63] ) );
  FA1A S2_19_62 ( .A(\ab[19][62] ), .B(\CARRYB[18][62] ), .CI(\SUMB[18][63] ), 
        .CO(\CARRYB[19][62] ), .S(\SUMB[19][62] ) );
  FA1A S2_19_61 ( .A(\ab[19][61] ), .B(\CARRYB[18][61] ), .CI(\SUMB[18][62] ), 
        .CO(\CARRYB[19][61] ), .S(\SUMB[19][61] ) );
  FA1A S2_19_52 ( .A(\ab[19][52] ), .B(\CARRYB[18][52] ), .CI(\SUMB[18][53] ), 
        .CO(\CARRYB[19][52] ), .S(\SUMB[19][52] ) );
  FA1A S2_19_44 ( .A(\ab[19][44] ), .B(\CARRYB[18][44] ), .CI(\SUMB[18][45] ), 
        .CO(\CARRYB[19][44] ), .S(\SUMB[19][44] ) );
  FA1A S2_19_43 ( .A(\ab[19][43] ), .B(\CARRYB[18][43] ), .CI(\SUMB[18][44] ), 
        .CO(\CARRYB[19][43] ), .S(\SUMB[19][43] ) );
  FA1A S2_19_42 ( .A(\ab[19][42] ), .B(\CARRYB[18][42] ), .CI(\SUMB[18][43] ), 
        .CO(\CARRYB[19][42] ), .S(\SUMB[19][42] ) );
  FA1A S2_19_41 ( .A(\ab[19][41] ), .B(\CARRYB[18][41] ), .CI(\SUMB[18][42] ), 
        .CO(\CARRYB[19][41] ), .S(\SUMB[19][41] ) );
  FA1A S2_19_40 ( .A(\ab[19][40] ), .B(\CARRYB[18][40] ), .CI(\SUMB[18][41] ), 
        .CO(\CARRYB[19][40] ), .S(\SUMB[19][40] ) );
  FA1A S2_19_39 ( .A(\ab[19][39] ), .B(\CARRYB[18][39] ), .CI(\SUMB[18][40] ), 
        .CO(\CARRYB[19][39] ), .S(\SUMB[19][39] ) );
  FA1A S2_18_63 ( .A(\ab[18][63] ), .B(\CARRYB[17][63] ), .CI(\SUMB[17][64] ), 
        .CO(\CARRYB[18][63] ), .S(\SUMB[18][63] ) );
  FA1A S2_18_62 ( .A(\ab[18][62] ), .B(\CARRYB[17][62] ), .CI(\SUMB[17][63] ), 
        .CO(\CARRYB[18][62] ), .S(\SUMB[18][62] ) );
  FA1A S2_18_61 ( .A(\ab[18][61] ), .B(\CARRYB[17][61] ), .CI(\SUMB[17][62] ), 
        .CO(\CARRYB[18][61] ), .S(\SUMB[18][61] ) );
  FA1A S2_18_52 ( .A(\ab[18][52] ), .B(\CARRYB[17][52] ), .CI(\SUMB[17][53] ), 
        .CO(\CARRYB[18][52] ), .S(\SUMB[18][52] ) );
  FA1A S2_18_44 ( .A(\ab[18][44] ), .B(\CARRYB[17][44] ), .CI(\SUMB[17][45] ), 
        .CO(\CARRYB[18][44] ), .S(\SUMB[18][44] ) );
  FA1A S2_18_43 ( .A(\ab[18][43] ), .B(\CARRYB[17][43] ), .CI(\SUMB[17][44] ), 
        .CO(\CARRYB[18][43] ), .S(\SUMB[18][43] ) );
  FA1A S2_18_42 ( .A(\ab[18][42] ), .B(\CARRYB[17][42] ), .CI(\SUMB[17][43] ), 
        .CO(\CARRYB[18][42] ), .S(\SUMB[18][42] ) );
  FA1A S2_18_41 ( .A(\ab[18][41] ), .B(\CARRYB[17][41] ), .CI(\SUMB[17][42] ), 
        .CO(\CARRYB[18][41] ), .S(\SUMB[18][41] ) );
  FA1A S2_18_40 ( .A(\ab[18][40] ), .B(\CARRYB[17][40] ), .CI(\SUMB[17][41] ), 
        .CO(\CARRYB[18][40] ), .S(\SUMB[18][40] ) );
  FA1A S2_18_39 ( .A(\ab[18][39] ), .B(\CARRYB[17][39] ), .CI(\SUMB[17][40] ), 
        .CO(\CARRYB[18][39] ), .S(\SUMB[18][39] ) );
  FA1A S2_17_63 ( .A(\ab[17][63] ), .B(\CARRYB[16][63] ), .CI(\SUMB[16][64] ), 
        .CO(\CARRYB[17][63] ), .S(\SUMB[17][63] ) );
  FA1A S2_17_62 ( .A(\ab[17][62] ), .B(\CARRYB[16][62] ), .CI(\SUMB[16][63] ), 
        .CO(\CARRYB[17][62] ), .S(\SUMB[17][62] ) );
  FA1A S2_17_61 ( .A(\ab[17][61] ), .B(\CARRYB[16][61] ), .CI(\SUMB[16][62] ), 
        .CO(\CARRYB[17][61] ), .S(\SUMB[17][61] ) );
  FA1A S2_17_52 ( .A(\ab[17][52] ), .B(\CARRYB[16][52] ), .CI(\SUMB[16][53] ), 
        .CO(\CARRYB[17][52] ), .S(\SUMB[17][52] ) );
  FA1A S2_17_44 ( .A(\ab[17][44] ), .B(\CARRYB[16][44] ), .CI(\SUMB[16][45] ), 
        .CO(\CARRYB[17][44] ), .S(\SUMB[17][44] ) );
  FA1A S2_17_43 ( .A(\ab[17][43] ), .B(\CARRYB[16][43] ), .CI(\SUMB[16][44] ), 
        .CO(\CARRYB[17][43] ), .S(\SUMB[17][43] ) );
  FA1A S2_17_42 ( .A(\ab[17][42] ), .B(\CARRYB[16][42] ), .CI(\SUMB[16][43] ), 
        .CO(\CARRYB[17][42] ), .S(\SUMB[17][42] ) );
  FA1A S2_17_41 ( .A(\ab[17][41] ), .B(\CARRYB[16][41] ), .CI(\SUMB[16][42] ), 
        .CO(\CARRYB[17][41] ), .S(\SUMB[17][41] ) );
  FA1A S2_17_40 ( .A(\ab[17][40] ), .B(\CARRYB[16][40] ), .CI(\SUMB[16][41] ), 
        .CO(\CARRYB[17][40] ), .S(\SUMB[17][40] ) );
  FA1A S2_17_39 ( .A(\ab[17][39] ), .B(\CARRYB[16][39] ), .CI(\SUMB[16][40] ), 
        .CO(\CARRYB[17][39] ), .S(\SUMB[17][39] ) );
  FA1A S2_16_63 ( .A(\ab[16][63] ), .B(\CARRYB[15][63] ), .CI(\SUMB[15][64] ), 
        .CO(\CARRYB[16][63] ), .S(\SUMB[16][63] ) );
  FA1A S2_16_62 ( .A(\ab[16][62] ), .B(\CARRYB[15][62] ), .CI(\SUMB[15][63] ), 
        .CO(\CARRYB[16][62] ), .S(\SUMB[16][62] ) );
  FA1A S2_16_61 ( .A(\ab[16][61] ), .B(\CARRYB[15][61] ), .CI(\SUMB[15][62] ), 
        .CO(\CARRYB[16][61] ), .S(\SUMB[16][61] ) );
  FA1A S2_16_52 ( .A(\ab[16][52] ), .B(\CARRYB[15][52] ), .CI(\SUMB[15][53] ), 
        .CO(\CARRYB[16][52] ), .S(\SUMB[16][52] ) );
  FA1A S2_16_44 ( .A(\ab[16][44] ), .B(\CARRYB[15][44] ), .CI(\SUMB[15][45] ), 
        .CO(\CARRYB[16][44] ), .S(\SUMB[16][44] ) );
  FA1A S2_16_43 ( .A(\ab[16][43] ), .B(\CARRYB[15][43] ), .CI(\SUMB[15][44] ), 
        .CO(\CARRYB[16][43] ), .S(\SUMB[16][43] ) );
  FA1A S2_16_42 ( .A(\ab[16][42] ), .B(\CARRYB[15][42] ), .CI(\SUMB[15][43] ), 
        .CO(\CARRYB[16][42] ), .S(\SUMB[16][42] ) );
  FA1A S2_16_41 ( .A(\ab[16][41] ), .B(\CARRYB[15][41] ), .CI(\SUMB[15][42] ), 
        .CO(\CARRYB[16][41] ), .S(\SUMB[16][41] ) );
  FA1A S2_16_40 ( .A(\ab[16][40] ), .B(\CARRYB[15][40] ), .CI(\SUMB[15][41] ), 
        .CO(\CARRYB[16][40] ), .S(\SUMB[16][40] ) );
  FA1A S2_16_39 ( .A(\ab[16][39] ), .B(\CARRYB[15][39] ), .CI(\SUMB[15][40] ), 
        .CO(\CARRYB[16][39] ), .S(\SUMB[16][39] ) );
  FA1A S2_15_63 ( .A(\ab[15][63] ), .B(\CARRYB[14][63] ), .CI(\SUMB[14][64] ), 
        .CO(\CARRYB[15][63] ), .S(\SUMB[15][63] ) );
  FA1A S2_15_62 ( .A(\ab[15][62] ), .B(\CARRYB[14][62] ), .CI(\SUMB[14][63] ), 
        .CO(\CARRYB[15][62] ), .S(\SUMB[15][62] ) );
  FA1A S2_15_61 ( .A(\ab[15][61] ), .B(\CARRYB[14][61] ), .CI(\SUMB[14][62] ), 
        .CO(\CARRYB[15][61] ), .S(\SUMB[15][61] ) );
  FA1A S2_15_52 ( .A(\ab[15][52] ), .B(\CARRYB[14][52] ), .CI(\SUMB[14][53] ), 
        .CO(\CARRYB[15][52] ), .S(\SUMB[15][52] ) );
  FA1A S2_15_44 ( .A(\ab[15][44] ), .B(\CARRYB[14][44] ), .CI(\SUMB[14][45] ), 
        .CO(\CARRYB[15][44] ), .S(\SUMB[15][44] ) );
  FA1A S2_15_43 ( .A(\ab[15][43] ), .B(\CARRYB[14][43] ), .CI(\SUMB[14][44] ), 
        .CO(\CARRYB[15][43] ), .S(\SUMB[15][43] ) );
  FA1A S2_15_42 ( .A(\ab[15][42] ), .B(\CARRYB[14][42] ), .CI(\SUMB[14][43] ), 
        .CO(\CARRYB[15][42] ), .S(\SUMB[15][42] ) );
  FA1A S2_15_41 ( .A(\ab[15][41] ), .B(\CARRYB[14][41] ), .CI(\SUMB[14][42] ), 
        .CO(\CARRYB[15][41] ), .S(\SUMB[15][41] ) );
  FA1A S2_15_40 ( .A(\ab[15][40] ), .B(\CARRYB[14][40] ), .CI(\SUMB[14][41] ), 
        .CO(\CARRYB[15][40] ), .S(\SUMB[15][40] ) );
  FA1A S2_15_38 ( .A(\ab[15][38] ), .B(\CARRYB[14][38] ), .CI(\SUMB[14][39] ), 
        .CO(\CARRYB[15][38] ), .S(\SUMB[15][38] ) );
  FA1A S2_15_39 ( .A(\ab[15][39] ), .B(\CARRYB[14][39] ), .CI(\SUMB[14][40] ), 
        .CO(\CARRYB[15][39] ), .S(\SUMB[15][39] ) );
  FA1A S2_14_38 ( .A(\ab[14][38] ), .B(\CARRYB[13][38] ), .CI(\SUMB[13][39] ), 
        .CO(\CARRYB[14][38] ), .S(\SUMB[14][38] ) );
  FA1A S2_13_38 ( .A(\ab[13][38] ), .B(\CARRYB[12][38] ), .CI(\SUMB[12][39] ), 
        .CO(\CARRYB[13][38] ), .S(\SUMB[13][38] ) );
  FA1A S2_12_38 ( .A(\ab[12][38] ), .B(\CARRYB[11][38] ), .CI(\SUMB[11][39] ), 
        .CO(\CARRYB[12][38] ), .S(\SUMB[12][38] ) );
  FA1A S2_11_38 ( .A(\ab[11][38] ), .B(\CARRYB[10][38] ), .CI(\SUMB[10][39] ), 
        .CO(\CARRYB[11][38] ), .S(\SUMB[11][38] ) );
  FA1A S2_10_38 ( .A(\ab[10][38] ), .B(\CARRYB[9][38] ), .CI(\SUMB[9][39] ), 
        .CO(\CARRYB[10][38] ), .S(\SUMB[10][38] ) );
  FA1A S2_9_38 ( .A(\ab[9][38] ), .B(\CARRYB[8][38] ), .CI(\SUMB[8][39] ), 
        .CO(\CARRYB[9][38] ), .S(\SUMB[9][38] ) );
  FA1A S2_8_38 ( .A(\ab[8][38] ), .B(\CARRYB[7][38] ), .CI(\SUMB[7][39] ), 
        .CO(\CARRYB[8][38] ), .S(\SUMB[8][38] ) );
  FA1A S2_7_38 ( .A(\ab[7][38] ), .B(\CARRYB[6][38] ), .CI(\SUMB[6][39] ), 
        .CO(\CARRYB[7][38] ), .S(\SUMB[7][38] ) );
  FA1A S2_6_38 ( .A(\ab[6][38] ), .B(\CARRYB[5][38] ), .CI(\SUMB[5][39] ), 
        .CO(\CARRYB[6][38] ), .S(\SUMB[6][38] ) );
  FA1A S2_5_38 ( .A(\ab[5][38] ), .B(\CARRYB[4][38] ), .CI(\SUMB[4][39] ), 
        .CO(\CARRYB[5][38] ), .S(\SUMB[5][38] ) );
  FA1A S2_4_38 ( .A(\ab[4][38] ), .B(\CARRYB[3][38] ), .CI(\SUMB[3][39] ), 
        .CO(\CARRYB[4][38] ), .S(\SUMB[4][38] ) );
  FA1A S2_3_38 ( .A(\ab[3][38] ), .B(\CARRYB[2][38] ), .CI(\SUMB[2][39] ), 
        .CO(\CARRYB[3][38] ), .S(\SUMB[3][38] ) );
  FA1A S2_2_38 ( .A(\ab[2][38] ), .B(\CARRYB[1][38] ), .CI(\SUMB[1][39] ), 
        .CO(\CARRYB[2][38] ), .S(\SUMB[2][38] ) );
  FA1A S2_2_37 ( .A(\ab[2][37] ), .B(\CARRYB[1][37] ), .CI(\SUMB[1][38] ), 
        .CO(\CARRYB[2][37] ), .S(\SUMB[2][37] ) );
  FA1A S4_52 ( .A(\ab[29][52] ), .B(\CARRYB[28][52] ), .CI(\SUMB[28][53] ), 
        .CO(\CARRYB[29][52] ), .S(\SUMB[29][52] ) );
  FA1A S4_63 ( .A(\ab[29][63] ), .B(\CARRYB[28][63] ), .CI(\SUMB[28][64] ), 
        .CO(\CARRYB[29][63] ), .S(\SUMB[29][63] ) );
  FA1A S4_47 ( .A(\ab[29][47] ), .B(\CARRYB[28][47] ), .CI(\SUMB[28][48] ), 
        .CO(\CARRYB[29][47] ), .S(\SUMB[29][47] ) );
  FA1A S4_46 ( .A(\ab[29][46] ), .B(\CARRYB[28][46] ), .CI(\SUMB[28][47] ), 
        .CO(\CARRYB[29][46] ), .S(\SUMB[29][46] ) );
  FA1A S2_28_47 ( .A(\ab[28][47] ), .B(\CARRYB[27][47] ), .CI(\SUMB[27][48] ), 
        .CO(\CARRYB[28][47] ), .S(\SUMB[28][47] ) );
  FA1A S4_49 ( .A(\ab[29][49] ), .B(\CARRYB[28][49] ), .CI(\SUMB[28][50] ), 
        .CO(\CARRYB[29][49] ), .S(\SUMB[29][49] ) );
  FA1A S4_50 ( .A(\ab[29][50] ), .B(\CARRYB[28][50] ), .CI(\SUMB[28][51] ), 
        .CO(\CARRYB[29][50] ), .S(\SUMB[29][50] ) );
  FA1A S4_45 ( .A(\ab[29][45] ), .B(\CARRYB[28][45] ), .CI(\SUMB[28][46] ), 
        .CO(\CARRYB[29][45] ), .S(\SUMB[29][45] ) );
  FA1A S2_28_49 ( .A(\ab[28][49] ), .B(\CARRYB[27][49] ), .CI(\SUMB[27][50] ), 
        .CO(\CARRYB[28][49] ), .S(\SUMB[28][49] ) );
  FA1A S2_28_48 ( .A(\ab[28][48] ), .B(\CARRYB[27][48] ), .CI(\SUMB[27][49] ), 
        .CO(\CARRYB[28][48] ), .S(\SUMB[28][48] ) );
  FA1A S2_28_50 ( .A(\ab[28][50] ), .B(\CARRYB[27][50] ), .CI(\SUMB[27][51] ), 
        .CO(\CARRYB[28][50] ), .S(\SUMB[28][50] ) );
  FA1A S2_28_51 ( .A(\ab[28][51] ), .B(\CARRYB[27][51] ), .CI(\SUMB[27][52] ), 
        .CO(\CARRYB[28][51] ), .S(\SUMB[28][51] ) );
  FA1A S2_28_46 ( .A(\ab[28][46] ), .B(\CARRYB[27][46] ), .CI(\SUMB[27][47] ), 
        .CO(\CARRYB[28][46] ), .S(\SUMB[28][46] ) );
  FA1A S2_28_45 ( .A(\ab[28][45] ), .B(\CARRYB[27][45] ), .CI(\SUMB[27][46] ), 
        .CO(\CARRYB[28][45] ), .S(\SUMB[28][45] ) );
  FA1A S2_27_50 ( .A(\ab[27][50] ), .B(\CARRYB[26][50] ), .CI(\SUMB[26][51] ), 
        .CO(\CARRYB[27][50] ), .S(\SUMB[27][50] ) );
  FA1A S2_27_49 ( .A(\ab[27][49] ), .B(\CARRYB[26][49] ), .CI(\SUMB[26][50] ), 
        .CO(\CARRYB[27][49] ), .S(\SUMB[27][49] ) );
  FA1A S2_27_48 ( .A(\ab[27][48] ), .B(\CARRYB[26][48] ), .CI(\SUMB[26][49] ), 
        .CO(\CARRYB[27][48] ), .S(\SUMB[27][48] ) );
  FA1A S2_27_51 ( .A(\ab[27][51] ), .B(\CARRYB[26][51] ), .CI(\SUMB[26][52] ), 
        .CO(\CARRYB[27][51] ), .S(\SUMB[27][51] ) );
  FA1A S2_27_47 ( .A(\ab[27][47] ), .B(\CARRYB[26][47] ), .CI(\SUMB[26][48] ), 
        .CO(\CARRYB[27][47] ), .S(\SUMB[27][47] ) );
  FA1A S2_27_46 ( .A(\ab[27][46] ), .B(\CARRYB[26][46] ), .CI(\SUMB[26][47] ), 
        .CO(\CARRYB[27][46] ), .S(\SUMB[27][46] ) );
  FA1A S2_27_45 ( .A(\ab[27][45] ), .B(\CARRYB[26][45] ), .CI(\SUMB[26][46] ), 
        .CO(\CARRYB[27][45] ), .S(\SUMB[27][45] ) );
  FA1A S2_26_45 ( .A(\ab[26][45] ), .B(\CARRYB[25][45] ), .CI(\SUMB[25][46] ), 
        .CO(\CARRYB[26][45] ), .S(\SUMB[26][45] ) );
  FA1A S2_26_51 ( .A(\ab[26][51] ), .B(\CARRYB[25][51] ), .CI(\SUMB[25][52] ), 
        .CO(\CARRYB[26][51] ), .S(\SUMB[26][51] ) );
  FA1A S2_26_50 ( .A(\ab[26][50] ), .B(\CARRYB[25][50] ), .CI(\SUMB[25][51] ), 
        .CO(\CARRYB[26][50] ), .S(\SUMB[26][50] ) );
  FA1A S2_26_49 ( .A(\ab[26][49] ), .B(\CARRYB[25][49] ), .CI(\SUMB[25][50] ), 
        .CO(\CARRYB[26][49] ), .S(\SUMB[26][49] ) );
  FA1A S2_26_48 ( .A(\ab[26][48] ), .B(\CARRYB[25][48] ), .CI(\SUMB[25][49] ), 
        .CO(\CARRYB[26][48] ), .S(\SUMB[26][48] ) );
  FA1A S2_26_47 ( .A(\ab[26][47] ), .B(\CARRYB[25][47] ), .CI(\SUMB[25][48] ), 
        .CO(\CARRYB[26][47] ), .S(\SUMB[26][47] ) );
  FA1A S2_26_46 ( .A(\ab[26][46] ), .B(\CARRYB[25][46] ), .CI(\SUMB[25][47] ), 
        .CO(\CARRYB[26][46] ), .S(\SUMB[26][46] ) );
  FA1A S2_25_46 ( .A(\ab[25][46] ), .B(\CARRYB[24][46] ), .CI(\SUMB[24][47] ), 
        .CO(\CARRYB[25][46] ), .S(\SUMB[25][46] ) );
  FA1A S2_25_45 ( .A(\ab[25][45] ), .B(\CARRYB[24][45] ), .CI(\SUMB[24][46] ), 
        .CO(\CARRYB[25][45] ), .S(\SUMB[25][45] ) );
  FA1A S2_25_51 ( .A(\ab[25][51] ), .B(\CARRYB[24][51] ), .CI(\SUMB[24][52] ), 
        .CO(\CARRYB[25][51] ), .S(\SUMB[25][51] ) );
  FA1A S2_25_50 ( .A(\ab[25][50] ), .B(\CARRYB[24][50] ), .CI(\SUMB[24][51] ), 
        .CO(\CARRYB[25][50] ), .S(\SUMB[25][50] ) );
  FA1A S2_25_49 ( .A(\ab[25][49] ), .B(\CARRYB[24][49] ), .CI(\SUMB[24][50] ), 
        .CO(\CARRYB[25][49] ), .S(\SUMB[25][49] ) );
  FA1A S2_25_48 ( .A(\ab[25][48] ), .B(\CARRYB[24][48] ), .CI(\SUMB[24][49] ), 
        .CO(\CARRYB[25][48] ), .S(\SUMB[25][48] ) );
  FA1A S2_25_47 ( .A(\ab[25][47] ), .B(\CARRYB[24][47] ), .CI(\SUMB[24][48] ), 
        .CO(\CARRYB[25][47] ), .S(\SUMB[25][47] ) );
  FA1A S2_24_47 ( .A(\ab[24][47] ), .B(\CARRYB[23][47] ), .CI(\SUMB[23][48] ), 
        .CO(\CARRYB[24][47] ), .S(\SUMB[24][47] ) );
  FA1A S2_24_46 ( .A(\ab[24][46] ), .B(\CARRYB[23][46] ), .CI(\SUMB[23][47] ), 
        .CO(\CARRYB[24][46] ), .S(\SUMB[24][46] ) );
  FA1A S2_24_45 ( .A(\ab[24][45] ), .B(\CARRYB[23][45] ), .CI(\SUMB[23][46] ), 
        .CO(\CARRYB[24][45] ), .S(\SUMB[24][45] ) );
  FA1A S2_24_51 ( .A(\ab[24][51] ), .B(\CARRYB[23][51] ), .CI(\SUMB[23][52] ), 
        .CO(\CARRYB[24][51] ), .S(\SUMB[24][51] ) );
  FA1A S2_24_50 ( .A(\ab[24][50] ), .B(\CARRYB[23][50] ), .CI(\SUMB[23][51] ), 
        .CO(\CARRYB[24][50] ), .S(\SUMB[24][50] ) );
  FA1A S2_24_49 ( .A(\ab[24][49] ), .B(\CARRYB[23][49] ), .CI(\SUMB[23][50] ), 
        .CO(\CARRYB[24][49] ), .S(\SUMB[24][49] ) );
  FA1A S2_24_48 ( .A(\ab[24][48] ), .B(\CARRYB[23][48] ), .CI(\SUMB[23][49] ), 
        .CO(\CARRYB[24][48] ), .S(\SUMB[24][48] ) );
  FA1A S2_23_48 ( .A(\ab[23][48] ), .B(\CARRYB[22][48] ), .CI(\SUMB[22][49] ), 
        .CO(\CARRYB[23][48] ), .S(\SUMB[23][48] ) );
  FA1A S2_23_47 ( .A(\ab[23][47] ), .B(\CARRYB[22][47] ), .CI(\SUMB[22][48] ), 
        .CO(\CARRYB[23][47] ), .S(\SUMB[23][47] ) );
  FA1A S2_23_46 ( .A(\ab[23][46] ), .B(\CARRYB[22][46] ), .CI(\SUMB[22][47] ), 
        .CO(\CARRYB[23][46] ), .S(\SUMB[23][46] ) );
  FA1A S2_23_45 ( .A(\ab[23][45] ), .B(\CARRYB[22][45] ), .CI(\SUMB[22][46] ), 
        .CO(\CARRYB[23][45] ), .S(\SUMB[23][45] ) );
  FA1A S2_23_51 ( .A(\ab[23][51] ), .B(\CARRYB[22][51] ), .CI(\SUMB[22][52] ), 
        .CO(\CARRYB[23][51] ), .S(\SUMB[23][51] ) );
  FA1A S2_23_50 ( .A(\ab[23][50] ), .B(\CARRYB[22][50] ), .CI(\SUMB[22][51] ), 
        .CO(\CARRYB[23][50] ), .S(\SUMB[23][50] ) );
  FA1A S2_23_49 ( .A(\ab[23][49] ), .B(\CARRYB[22][49] ), .CI(\SUMB[22][50] ), 
        .CO(\CARRYB[23][49] ), .S(\SUMB[23][49] ) );
  FA1A S2_22_49 ( .A(\ab[22][49] ), .B(\CARRYB[21][49] ), .CI(\SUMB[21][50] ), 
        .CO(\CARRYB[22][49] ), .S(\SUMB[22][49] ) );
  FA1A S2_22_48 ( .A(\ab[22][48] ), .B(\CARRYB[21][48] ), .CI(\SUMB[21][49] ), 
        .CO(\CARRYB[22][48] ), .S(\SUMB[22][48] ) );
  FA1A S2_22_47 ( .A(\ab[22][47] ), .B(\CARRYB[21][47] ), .CI(\SUMB[21][48] ), 
        .CO(\CARRYB[22][47] ), .S(\SUMB[22][47] ) );
  FA1A S2_22_46 ( .A(\ab[22][46] ), .B(\CARRYB[21][46] ), .CI(\SUMB[21][47] ), 
        .CO(\CARRYB[22][46] ), .S(\SUMB[22][46] ) );
  FA1A S2_22_45 ( .A(\ab[22][45] ), .B(\CARRYB[21][45] ), .CI(\SUMB[21][46] ), 
        .CO(\CARRYB[22][45] ), .S(\SUMB[22][45] ) );
  FA1A S2_22_51 ( .A(\ab[22][51] ), .B(\CARRYB[21][51] ), .CI(\SUMB[21][52] ), 
        .CO(\CARRYB[22][51] ), .S(\SUMB[22][51] ) );
  FA1A S2_22_50 ( .A(\ab[22][50] ), .B(\CARRYB[21][50] ), .CI(\SUMB[21][51] ), 
        .CO(\CARRYB[22][50] ), .S(\SUMB[22][50] ) );
  FA1A S2_21_50 ( .A(\ab[21][50] ), .B(\CARRYB[20][50] ), .CI(\SUMB[20][51] ), 
        .CO(\CARRYB[21][50] ), .S(\SUMB[21][50] ) );
  FA1A S2_21_49 ( .A(\ab[21][49] ), .B(\CARRYB[20][49] ), .CI(\SUMB[20][50] ), 
        .CO(\CARRYB[21][49] ), .S(\SUMB[21][49] ) );
  FA1A S2_21_48 ( .A(\ab[21][48] ), .B(\CARRYB[20][48] ), .CI(\SUMB[20][49] ), 
        .CO(\CARRYB[21][48] ), .S(\SUMB[21][48] ) );
  FA1A S2_21_47 ( .A(\ab[21][47] ), .B(\CARRYB[20][47] ), .CI(\SUMB[20][48] ), 
        .CO(\CARRYB[21][47] ), .S(\SUMB[21][47] ) );
  FA1A S2_21_46 ( .A(\ab[21][46] ), .B(\CARRYB[20][46] ), .CI(\SUMB[20][47] ), 
        .CO(\CARRYB[21][46] ), .S(\SUMB[21][46] ) );
  FA1A S2_21_45 ( .A(\ab[21][45] ), .B(\CARRYB[20][45] ), .CI(\SUMB[20][46] ), 
        .CO(\CARRYB[21][45] ), .S(\SUMB[21][45] ) );
  FA1A S2_21_51 ( .A(\ab[21][51] ), .B(\CARRYB[20][51] ), .CI(\SUMB[20][52] ), 
        .CO(\CARRYB[21][51] ), .S(\SUMB[21][51] ) );
  FA1A S2_20_51 ( .A(\ab[20][51] ), .B(\CARRYB[19][51] ), .CI(\SUMB[19][52] ), 
        .CO(\CARRYB[20][51] ), .S(\SUMB[20][51] ) );
  FA1A S2_20_50 ( .A(\ab[20][50] ), .B(\CARRYB[19][50] ), .CI(\SUMB[19][51] ), 
        .CO(\CARRYB[20][50] ), .S(\SUMB[20][50] ) );
  FA1A S2_20_49 ( .A(\ab[20][49] ), .B(\CARRYB[19][49] ), .CI(\SUMB[19][50] ), 
        .CO(\CARRYB[20][49] ), .S(\SUMB[20][49] ) );
  FA1A S2_20_48 ( .A(\ab[20][48] ), .B(\CARRYB[19][48] ), .CI(\SUMB[19][49] ), 
        .CO(\CARRYB[20][48] ), .S(\SUMB[20][48] ) );
  FA1A S2_20_47 ( .A(\ab[20][47] ), .B(\CARRYB[19][47] ), .CI(\SUMB[19][48] ), 
        .CO(\CARRYB[20][47] ), .S(\SUMB[20][47] ) );
  FA1A S2_20_46 ( .A(\ab[20][46] ), .B(\CARRYB[19][46] ), .CI(\SUMB[19][47] ), 
        .CO(\CARRYB[20][46] ), .S(\SUMB[20][46] ) );
  FA1A S2_20_45 ( .A(\ab[20][45] ), .B(\CARRYB[19][45] ), .CI(\SUMB[19][46] ), 
        .CO(\CARRYB[20][45] ), .S(\SUMB[20][45] ) );
  FA1A S2_19_51 ( .A(\ab[19][51] ), .B(\CARRYB[18][51] ), .CI(\SUMB[18][52] ), 
        .CO(\CARRYB[19][51] ), .S(\SUMB[19][51] ) );
  FA1A S2_19_50 ( .A(\ab[19][50] ), .B(\CARRYB[18][50] ), .CI(\SUMB[18][51] ), 
        .CO(\CARRYB[19][50] ), .S(\SUMB[19][50] ) );
  FA1A S2_19_49 ( .A(\ab[19][49] ), .B(\CARRYB[18][49] ), .CI(\SUMB[18][50] ), 
        .CO(\CARRYB[19][49] ), .S(\SUMB[19][49] ) );
  FA1A S2_19_48 ( .A(\ab[19][48] ), .B(\CARRYB[18][48] ), .CI(\SUMB[18][49] ), 
        .CO(\CARRYB[19][48] ), .S(\SUMB[19][48] ) );
  FA1A S2_19_47 ( .A(\ab[19][47] ), .B(\CARRYB[18][47] ), .CI(\SUMB[18][48] ), 
        .CO(\CARRYB[19][47] ), .S(\SUMB[19][47] ) );
  FA1A S2_19_46 ( .A(\ab[19][46] ), .B(\CARRYB[18][46] ), .CI(\SUMB[18][47] ), 
        .CO(\CARRYB[19][46] ), .S(\SUMB[19][46] ) );
  FA1A S2_19_45 ( .A(\ab[19][45] ), .B(\CARRYB[18][45] ), .CI(\SUMB[18][46] ), 
        .CO(\CARRYB[19][45] ), .S(\SUMB[19][45] ) );
  FA1A S2_18_51 ( .A(\ab[18][51] ), .B(\CARRYB[17][51] ), .CI(\SUMB[17][52] ), 
        .CO(\CARRYB[18][51] ), .S(\SUMB[18][51] ) );
  FA1A S2_18_50 ( .A(\ab[18][50] ), .B(\CARRYB[17][50] ), .CI(\SUMB[17][51] ), 
        .CO(\CARRYB[18][50] ), .S(\SUMB[18][50] ) );
  FA1A S2_18_49 ( .A(\ab[18][49] ), .B(\CARRYB[17][49] ), .CI(\SUMB[17][50] ), 
        .CO(\CARRYB[18][49] ), .S(\SUMB[18][49] ) );
  FA1A S2_18_48 ( .A(\ab[18][48] ), .B(\CARRYB[17][48] ), .CI(\SUMB[17][49] ), 
        .CO(\CARRYB[18][48] ), .S(\SUMB[18][48] ) );
  FA1A S2_18_47 ( .A(\ab[18][47] ), .B(\CARRYB[17][47] ), .CI(\SUMB[17][48] ), 
        .CO(\CARRYB[18][47] ), .S(\SUMB[18][47] ) );
  FA1A S2_18_46 ( .A(\ab[18][46] ), .B(\CARRYB[17][46] ), .CI(\SUMB[17][47] ), 
        .CO(\CARRYB[18][46] ), .S(\SUMB[18][46] ) );
  FA1A S2_18_45 ( .A(\ab[18][45] ), .B(\CARRYB[17][45] ), .CI(\SUMB[17][46] ), 
        .CO(\CARRYB[18][45] ), .S(\SUMB[18][45] ) );
  FA1A S2_17_51 ( .A(\ab[17][51] ), .B(\CARRYB[16][51] ), .CI(\SUMB[16][52] ), 
        .CO(\CARRYB[17][51] ), .S(\SUMB[17][51] ) );
  FA1A S2_17_50 ( .A(\ab[17][50] ), .B(\CARRYB[16][50] ), .CI(\SUMB[16][51] ), 
        .CO(\CARRYB[17][50] ), .S(\SUMB[17][50] ) );
  FA1A S2_17_49 ( .A(\ab[17][49] ), .B(\CARRYB[16][49] ), .CI(\SUMB[16][50] ), 
        .CO(\CARRYB[17][49] ), .S(\SUMB[17][49] ) );
  FA1A S2_17_48 ( .A(\ab[17][48] ), .B(\CARRYB[16][48] ), .CI(\SUMB[16][49] ), 
        .CO(\CARRYB[17][48] ), .S(\SUMB[17][48] ) );
  FA1A S2_17_47 ( .A(\ab[17][47] ), .B(\CARRYB[16][47] ), .CI(\SUMB[16][48] ), 
        .CO(\CARRYB[17][47] ), .S(\SUMB[17][47] ) );
  FA1A S2_17_46 ( .A(\ab[17][46] ), .B(\CARRYB[16][46] ), .CI(\SUMB[16][47] ), 
        .CO(\CARRYB[17][46] ), .S(\SUMB[17][46] ) );
  FA1A S2_17_45 ( .A(\ab[17][45] ), .B(\CARRYB[16][45] ), .CI(\SUMB[16][46] ), 
        .CO(\CARRYB[17][45] ), .S(\SUMB[17][45] ) );
  FA1A S2_16_51 ( .A(\ab[16][51] ), .B(\CARRYB[15][51] ), .CI(\SUMB[15][52] ), 
        .CO(\CARRYB[16][51] ), .S(\SUMB[16][51] ) );
  FA1A S2_16_50 ( .A(\ab[16][50] ), .B(\CARRYB[15][50] ), .CI(\SUMB[15][51] ), 
        .CO(\CARRYB[16][50] ), .S(\SUMB[16][50] ) );
  FA1A S2_16_49 ( .A(\ab[16][49] ), .B(\CARRYB[15][49] ), .CI(\SUMB[15][50] ), 
        .CO(\CARRYB[16][49] ), .S(\SUMB[16][49] ) );
  FA1A S2_16_48 ( .A(\ab[16][48] ), .B(\CARRYB[15][48] ), .CI(\SUMB[15][49] ), 
        .CO(\CARRYB[16][48] ), .S(\SUMB[16][48] ) );
  FA1A S2_16_47 ( .A(\ab[16][47] ), .B(\CARRYB[15][47] ), .CI(\SUMB[15][48] ), 
        .CO(\CARRYB[16][47] ), .S(\SUMB[16][47] ) );
  FA1A S2_16_46 ( .A(\ab[16][46] ), .B(\CARRYB[15][46] ), .CI(\SUMB[15][47] ), 
        .CO(\CARRYB[16][46] ), .S(\SUMB[16][46] ) );
  FA1A S2_16_45 ( .A(\ab[16][45] ), .B(\CARRYB[15][45] ), .CI(\SUMB[15][46] ), 
        .CO(\CARRYB[16][45] ), .S(\SUMB[16][45] ) );
  FA1A S2_15_51 ( .A(\ab[15][51] ), .B(\CARRYB[14][51] ), .CI(\SUMB[14][52] ), 
        .CO(\CARRYB[15][51] ), .S(\SUMB[15][51] ) );
  FA1A S2_15_50 ( .A(\ab[15][50] ), .B(\CARRYB[14][50] ), .CI(\SUMB[14][51] ), 
        .CO(\CARRYB[15][50] ), .S(\SUMB[15][50] ) );
  FA1A S2_15_49 ( .A(\ab[15][49] ), .B(\CARRYB[14][49] ), .CI(\SUMB[14][50] ), 
        .CO(\CARRYB[15][49] ), .S(\SUMB[15][49] ) );
  FA1A S2_15_48 ( .A(\ab[15][48] ), .B(\CARRYB[14][48] ), .CI(\SUMB[14][49] ), 
        .CO(\CARRYB[15][48] ), .S(\SUMB[15][48] ) );
  FA1A S2_15_47 ( .A(\ab[15][47] ), .B(\CARRYB[14][47] ), .CI(\SUMB[14][48] ), 
        .CO(\CARRYB[15][47] ), .S(\SUMB[15][47] ) );
  FA1A S2_15_46 ( .A(\ab[15][46] ), .B(\CARRYB[14][46] ), .CI(\SUMB[14][47] ), 
        .CO(\CARRYB[15][46] ), .S(\SUMB[15][46] ) );
  FA1A S2_15_45 ( .A(\ab[15][45] ), .B(\CARRYB[14][45] ), .CI(\SUMB[14][46] ), 
        .CO(\CARRYB[15][45] ), .S(\SUMB[15][45] ) );
  FA1A S4_51 ( .A(\ab[29][51] ), .B(\CARRYB[28][51] ), .CI(\SUMB[28][52] ), 
        .CO(\CARRYB[29][51] ), .S(\SUMB[29][51] ) );
  FA1A S4_48 ( .A(\ab[29][48] ), .B(\CARRYB[28][48] ), .CI(\SUMB[28][49] ), 
        .CO(\CARRYB[29][48] ), .S(\SUMB[29][48] ) );
  FA1A S3_14_94 ( .A(\ab[14][94] ), .B(\CARRYB[13][94] ), .CI(\ab[13][95] ), 
        .CO(\CARRYB[14][94] ), .S(\SUMB[14][94] ) );
  FA1A S3_13_94 ( .A(\ab[13][94] ), .B(\CARRYB[12][94] ), .CI(\ab[12][95] ), 
        .CO(\CARRYB[13][94] ), .S(\SUMB[13][94] ) );
  FA1A S3_12_94 ( .A(\ab[12][94] ), .B(\CARRYB[11][94] ), .CI(\ab[11][95] ), 
        .CO(\CARRYB[12][94] ), .S(\SUMB[12][94] ) );
  FA1A S3_11_94 ( .A(\ab[11][94] ), .B(\CARRYB[10][94] ), .CI(\ab[10][95] ), 
        .CO(\CARRYB[11][94] ), .S(\SUMB[11][94] ) );
  FA1A S3_10_94 ( .A(\ab[10][94] ), .B(\CARRYB[9][94] ), .CI(\ab[9][95] ), 
        .CO(\CARRYB[10][94] ), .S(\SUMB[10][94] ) );
  FA1A S3_9_94 ( .A(\ab[9][94] ), .B(\CARRYB[8][94] ), .CI(\ab[8][95] ), .CO(
        \CARRYB[9][94] ), .S(\SUMB[9][94] ) );
  FA1A S3_8_94 ( .A(\ab[8][94] ), .B(\CARRYB[7][94] ), .CI(\ab[7][95] ), .CO(
        \CARRYB[8][94] ), .S(\SUMB[8][94] ) );
  FA1A S3_7_94 ( .A(\ab[7][94] ), .B(\CARRYB[6][94] ), .CI(\ab[6][95] ), .CO(
        \CARRYB[7][94] ), .S(\SUMB[7][94] ) );
  FA1A S3_6_94 ( .A(\ab[6][94] ), .B(\CARRYB[5][94] ), .CI(\ab[5][95] ), .CO(
        \CARRYB[6][94] ), .S(\SUMB[6][94] ) );
  FA1A S3_5_94 ( .A(\ab[5][94] ), .B(\CARRYB[4][94] ), .CI(\ab[4][95] ), .CO(
        \CARRYB[5][94] ), .S(\SUMB[5][94] ) );
  FA1A S3_4_94 ( .A(\ab[4][94] ), .B(\CARRYB[3][94] ), .CI(\ab[3][95] ), .CO(
        \CARRYB[4][94] ), .S(\SUMB[4][94] ) );
  FA1A S3_3_94 ( .A(\ab[3][94] ), .B(\CARRYB[2][94] ), .CI(\ab[2][95] ), .CO(
        \CARRYB[3][94] ), .S(\SUMB[3][94] ) );
  FA1A S3_2_94 ( .A(\ab[2][94] ), .B(\CARRYB[1][94] ), .CI(\ab[1][95] ), .CO(
        \CARRYB[2][94] ), .S(\SUMB[2][94] ) );
  FA1A S2_14_93 ( .A(\ab[14][93] ), .B(\CARRYB[13][93] ), .CI(\SUMB[13][94] ), 
        .CO(\CARRYB[14][93] ), .S(\SUMB[14][93] ) );
  FA1A S2_13_93 ( .A(\ab[13][93] ), .B(\CARRYB[12][93] ), .CI(\SUMB[12][94] ), 
        .CO(\CARRYB[13][93] ), .S(\SUMB[13][93] ) );
  FA1A S2_12_93 ( .A(\ab[12][93] ), .B(\CARRYB[11][93] ), .CI(\SUMB[11][94] ), 
        .CO(\CARRYB[12][93] ), .S(\SUMB[12][93] ) );
  FA1A S2_11_93 ( .A(\ab[11][93] ), .B(\CARRYB[10][93] ), .CI(\SUMB[10][94] ), 
        .CO(\CARRYB[11][93] ), .S(\SUMB[11][93] ) );
  FA1A S2_10_93 ( .A(\ab[10][93] ), .B(\CARRYB[9][93] ), .CI(\SUMB[9][94] ), 
        .CO(\CARRYB[10][93] ), .S(\SUMB[10][93] ) );
  FA1A S2_9_93 ( .A(\ab[9][93] ), .B(\CARRYB[8][93] ), .CI(\SUMB[8][94] ), 
        .CO(\CARRYB[9][93] ), .S(\SUMB[9][93] ) );
  FA1A S2_8_93 ( .A(\ab[8][93] ), .B(\CARRYB[7][93] ), .CI(\SUMB[7][94] ), 
        .CO(\CARRYB[8][93] ), .S(\SUMB[8][93] ) );
  FA1A S2_7_93 ( .A(\ab[7][93] ), .B(\CARRYB[6][93] ), .CI(\SUMB[6][94] ), 
        .CO(\CARRYB[7][93] ), .S(\SUMB[7][93] ) );
  FA1A S2_6_93 ( .A(\ab[6][93] ), .B(\CARRYB[5][93] ), .CI(\SUMB[5][94] ), 
        .CO(\CARRYB[6][93] ), .S(\SUMB[6][93] ) );
  FA1A S2_5_93 ( .A(\ab[5][93] ), .B(\CARRYB[4][93] ), .CI(\SUMB[4][94] ), 
        .CO(\CARRYB[5][93] ), .S(\SUMB[5][93] ) );
  FA1A S2_4_93 ( .A(\ab[4][93] ), .B(\CARRYB[3][93] ), .CI(\SUMB[3][94] ), 
        .CO(\CARRYB[4][93] ), .S(\SUMB[4][93] ) );
  FA1A S2_3_93 ( .A(\ab[3][93] ), .B(\CARRYB[2][93] ), .CI(\SUMB[2][94] ), 
        .CO(\CARRYB[3][93] ), .S(\SUMB[3][93] ) );
  FA1A S2_2_93 ( .A(\ab[2][93] ), .B(\CARRYB[1][93] ), .CI(\SUMB[1][94] ), 
        .CO(\CARRYB[2][93] ), .S(\SUMB[2][93] ) );
  FA1A S2_14_92 ( .A(\ab[14][92] ), .B(\CARRYB[13][92] ), .CI(\SUMB[13][93] ), 
        .CO(\CARRYB[14][92] ), .S(\SUMB[14][92] ) );
  FA1A S2_13_92 ( .A(\ab[13][92] ), .B(\CARRYB[12][92] ), .CI(\SUMB[12][93] ), 
        .CO(\CARRYB[13][92] ), .S(\SUMB[13][92] ) );
  FA1A S2_12_92 ( .A(\ab[12][92] ), .B(\CARRYB[11][92] ), .CI(\SUMB[11][93] ), 
        .CO(\CARRYB[12][92] ), .S(\SUMB[12][92] ) );
  FA1A S2_11_92 ( .A(\ab[11][92] ), .B(\CARRYB[10][92] ), .CI(\SUMB[10][93] ), 
        .CO(\CARRYB[11][92] ), .S(\SUMB[11][92] ) );
  FA1A S2_10_92 ( .A(\ab[10][92] ), .B(\CARRYB[9][92] ), .CI(\SUMB[9][93] ), 
        .CO(\CARRYB[10][92] ), .S(\SUMB[10][92] ) );
  FA1A S2_9_92 ( .A(\ab[9][92] ), .B(\CARRYB[8][92] ), .CI(\SUMB[8][93] ), 
        .CO(\CARRYB[9][92] ), .S(\SUMB[9][92] ) );
  FA1A S2_8_92 ( .A(\ab[8][92] ), .B(\CARRYB[7][92] ), .CI(\SUMB[7][93] ), 
        .CO(\CARRYB[8][92] ), .S(\SUMB[8][92] ) );
  FA1A S2_7_92 ( .A(\ab[7][92] ), .B(\CARRYB[6][92] ), .CI(\SUMB[6][93] ), 
        .CO(\CARRYB[7][92] ), .S(\SUMB[7][92] ) );
  FA1A S2_6_92 ( .A(\ab[6][92] ), .B(\CARRYB[5][92] ), .CI(\SUMB[5][93] ), 
        .CO(\CARRYB[6][92] ), .S(\SUMB[6][92] ) );
  FA1A S2_5_92 ( .A(\ab[5][92] ), .B(\CARRYB[4][92] ), .CI(\SUMB[4][93] ), 
        .CO(\CARRYB[5][92] ), .S(\SUMB[5][92] ) );
  FA1A S2_4_92 ( .A(\ab[4][92] ), .B(\CARRYB[3][92] ), .CI(\SUMB[3][93] ), 
        .CO(\CARRYB[4][92] ), .S(\SUMB[4][92] ) );
  FA1A S2_3_92 ( .A(\ab[3][92] ), .B(\CARRYB[2][92] ), .CI(\SUMB[2][93] ), 
        .CO(\CARRYB[3][92] ), .S(\SUMB[3][92] ) );
  FA1A S2_2_92 ( .A(\ab[2][92] ), .B(\CARRYB[1][92] ), .CI(\SUMB[1][93] ), 
        .CO(\CARRYB[2][92] ), .S(\SUMB[2][92] ) );
  FA1A S2_14_91 ( .A(\ab[14][91] ), .B(\CARRYB[13][91] ), .CI(\SUMB[13][92] ), 
        .CO(\CARRYB[14][91] ), .S(\SUMB[14][91] ) );
  FA1A S2_13_91 ( .A(\ab[13][91] ), .B(\CARRYB[12][91] ), .CI(\SUMB[12][92] ), 
        .CO(\CARRYB[13][91] ), .S(\SUMB[13][91] ) );
  FA1A S2_12_91 ( .A(\ab[12][91] ), .B(\CARRYB[11][91] ), .CI(\SUMB[11][92] ), 
        .CO(\CARRYB[12][91] ), .S(\SUMB[12][91] ) );
  FA1A S2_11_91 ( .A(\ab[11][91] ), .B(\CARRYB[10][91] ), .CI(\SUMB[10][92] ), 
        .CO(\CARRYB[11][91] ), .S(\SUMB[11][91] ) );
  FA1A S2_10_91 ( .A(\ab[10][91] ), .B(\CARRYB[9][91] ), .CI(\SUMB[9][92] ), 
        .CO(\CARRYB[10][91] ), .S(\SUMB[10][91] ) );
  FA1A S2_9_91 ( .A(\ab[9][91] ), .B(\CARRYB[8][91] ), .CI(\SUMB[8][92] ), 
        .CO(\CARRYB[9][91] ), .S(\SUMB[9][91] ) );
  FA1A S2_8_91 ( .A(\ab[8][91] ), .B(\CARRYB[7][91] ), .CI(\SUMB[7][92] ), 
        .CO(\CARRYB[8][91] ), .S(\SUMB[8][91] ) );
  FA1A S2_7_91 ( .A(\ab[7][91] ), .B(\CARRYB[6][91] ), .CI(\SUMB[6][92] ), 
        .CO(\CARRYB[7][91] ), .S(\SUMB[7][91] ) );
  FA1A S2_6_91 ( .A(\ab[6][91] ), .B(\CARRYB[5][91] ), .CI(\SUMB[5][92] ), 
        .CO(\CARRYB[6][91] ), .S(\SUMB[6][91] ) );
  FA1A S2_5_91 ( .A(\ab[5][91] ), .B(\CARRYB[4][91] ), .CI(\SUMB[4][92] ), 
        .CO(\CARRYB[5][91] ), .S(\SUMB[5][91] ) );
  FA1A S2_4_91 ( .A(\ab[4][91] ), .B(\CARRYB[3][91] ), .CI(\SUMB[3][92] ), 
        .CO(\CARRYB[4][91] ), .S(\SUMB[4][91] ) );
  FA1A S2_3_91 ( .A(\ab[3][91] ), .B(\CARRYB[2][91] ), .CI(\SUMB[2][92] ), 
        .CO(\CARRYB[3][91] ), .S(\SUMB[3][91] ) );
  FA1A S2_2_91 ( .A(\ab[2][91] ), .B(\CARRYB[1][91] ), .CI(\SUMB[1][92] ), 
        .CO(\CARRYB[2][91] ), .S(\SUMB[2][91] ) );
  FA1A S2_14_90 ( .A(\ab[14][90] ), .B(\CARRYB[13][90] ), .CI(\SUMB[13][91] ), 
        .CO(\CARRYB[14][90] ), .S(\SUMB[14][90] ) );
  FA1A S2_13_90 ( .A(\ab[13][90] ), .B(\CARRYB[12][90] ), .CI(\SUMB[12][91] ), 
        .CO(\CARRYB[13][90] ), .S(\SUMB[13][90] ) );
  FA1A S2_12_90 ( .A(\ab[12][90] ), .B(\CARRYB[11][90] ), .CI(\SUMB[11][91] ), 
        .CO(\CARRYB[12][90] ), .S(\SUMB[12][90] ) );
  FA1A S2_11_90 ( .A(\ab[11][90] ), .B(\CARRYB[10][90] ), .CI(\SUMB[10][91] ), 
        .CO(\CARRYB[11][90] ), .S(\SUMB[11][90] ) );
  FA1A S2_10_90 ( .A(\ab[10][90] ), .B(\CARRYB[9][90] ), .CI(\SUMB[9][91] ), 
        .CO(\CARRYB[10][90] ), .S(\SUMB[10][90] ) );
  FA1A S2_9_90 ( .A(\ab[9][90] ), .B(\CARRYB[8][90] ), .CI(\SUMB[8][91] ), 
        .CO(\CARRYB[9][90] ), .S(\SUMB[9][90] ) );
  FA1A S2_8_90 ( .A(\ab[8][90] ), .B(\CARRYB[7][90] ), .CI(\SUMB[7][91] ), 
        .CO(\CARRYB[8][90] ), .S(\SUMB[8][90] ) );
  FA1A S2_7_90 ( .A(\ab[7][90] ), .B(\CARRYB[6][90] ), .CI(\SUMB[6][91] ), 
        .CO(\CARRYB[7][90] ), .S(\SUMB[7][90] ) );
  FA1A S2_6_90 ( .A(\ab[6][90] ), .B(\CARRYB[5][90] ), .CI(\SUMB[5][91] ), 
        .CO(\CARRYB[6][90] ), .S(\SUMB[6][90] ) );
  FA1A S2_5_90 ( .A(\ab[5][90] ), .B(\CARRYB[4][90] ), .CI(\SUMB[4][91] ), 
        .CO(\CARRYB[5][90] ), .S(\SUMB[5][90] ) );
  FA1A S2_4_90 ( .A(\ab[4][90] ), .B(\CARRYB[3][90] ), .CI(\SUMB[3][91] ), 
        .CO(\CARRYB[4][90] ), .S(\SUMB[4][90] ) );
  FA1A S2_3_90 ( .A(\ab[3][90] ), .B(\CARRYB[2][90] ), .CI(\SUMB[2][91] ), 
        .CO(\CARRYB[3][90] ), .S(\SUMB[3][90] ) );
  FA1A S2_2_90 ( .A(\ab[2][90] ), .B(\CARRYB[1][90] ), .CI(\SUMB[1][91] ), 
        .CO(\CARRYB[2][90] ), .S(\SUMB[2][90] ) );
  FA1A S2_14_89 ( .A(\ab[14][89] ), .B(\CARRYB[13][89] ), .CI(\SUMB[13][90] ), 
        .CO(\CARRYB[14][89] ), .S(\SUMB[14][89] ) );
  FA1A S2_13_89 ( .A(\ab[13][89] ), .B(\CARRYB[12][89] ), .CI(\SUMB[12][90] ), 
        .CO(\CARRYB[13][89] ), .S(\SUMB[13][89] ) );
  FA1A S2_12_89 ( .A(\ab[12][89] ), .B(\CARRYB[11][89] ), .CI(\SUMB[11][90] ), 
        .CO(\CARRYB[12][89] ), .S(\SUMB[12][89] ) );
  FA1A S2_11_89 ( .A(\ab[11][89] ), .B(\CARRYB[10][89] ), .CI(\SUMB[10][90] ), 
        .CO(\CARRYB[11][89] ), .S(\SUMB[11][89] ) );
  FA1A S2_10_89 ( .A(\ab[10][89] ), .B(\CARRYB[9][89] ), .CI(\SUMB[9][90] ), 
        .CO(\CARRYB[10][89] ), .S(\SUMB[10][89] ) );
  FA1A S2_9_89 ( .A(\ab[9][89] ), .B(\CARRYB[8][89] ), .CI(\SUMB[8][90] ), 
        .CO(\CARRYB[9][89] ), .S(\SUMB[9][89] ) );
  FA1A S2_8_89 ( .A(\ab[8][89] ), .B(\CARRYB[7][89] ), .CI(\SUMB[7][90] ), 
        .CO(\CARRYB[8][89] ), .S(\SUMB[8][89] ) );
  FA1A S2_7_89 ( .A(\ab[7][89] ), .B(\CARRYB[6][89] ), .CI(\SUMB[6][90] ), 
        .CO(\CARRYB[7][89] ), .S(\SUMB[7][89] ) );
  FA1A S2_6_89 ( .A(\ab[6][89] ), .B(\CARRYB[5][89] ), .CI(\SUMB[5][90] ), 
        .CO(\CARRYB[6][89] ), .S(\SUMB[6][89] ) );
  FA1A S2_5_89 ( .A(\ab[5][89] ), .B(\CARRYB[4][89] ), .CI(\SUMB[4][90] ), 
        .CO(\CARRYB[5][89] ), .S(\SUMB[5][89] ) );
  FA1A S2_4_89 ( .A(\ab[4][89] ), .B(\CARRYB[3][89] ), .CI(\SUMB[3][90] ), 
        .CO(\CARRYB[4][89] ), .S(\SUMB[4][89] ) );
  FA1A S2_3_89 ( .A(\ab[3][89] ), .B(\CARRYB[2][89] ), .CI(\SUMB[2][90] ), 
        .CO(\CARRYB[3][89] ), .S(\SUMB[3][89] ) );
  FA1A S2_2_89 ( .A(\ab[2][89] ), .B(\CARRYB[1][89] ), .CI(\SUMB[1][90] ), 
        .CO(\CARRYB[2][89] ), .S(\SUMB[2][89] ) );
  FA1A S2_14_88 ( .A(\ab[14][88] ), .B(\CARRYB[13][88] ), .CI(\SUMB[13][89] ), 
        .CO(\CARRYB[14][88] ), .S(\SUMB[14][88] ) );
  FA1A S2_13_88 ( .A(\ab[13][88] ), .B(\CARRYB[12][88] ), .CI(\SUMB[12][89] ), 
        .CO(\CARRYB[13][88] ), .S(\SUMB[13][88] ) );
  FA1A S2_12_88 ( .A(\ab[12][88] ), .B(\CARRYB[11][88] ), .CI(\SUMB[11][89] ), 
        .CO(\CARRYB[12][88] ), .S(\SUMB[12][88] ) );
  FA1A S2_11_88 ( .A(\ab[11][88] ), .B(\CARRYB[10][88] ), .CI(\SUMB[10][89] ), 
        .CO(\CARRYB[11][88] ), .S(\SUMB[11][88] ) );
  FA1A S2_10_88 ( .A(\ab[10][88] ), .B(\CARRYB[9][88] ), .CI(\SUMB[9][89] ), 
        .CO(\CARRYB[10][88] ), .S(\SUMB[10][88] ) );
  FA1A S2_9_88 ( .A(\ab[9][88] ), .B(\CARRYB[8][88] ), .CI(\SUMB[8][89] ), 
        .CO(\CARRYB[9][88] ), .S(\SUMB[9][88] ) );
  FA1A S2_8_88 ( .A(\ab[8][88] ), .B(\CARRYB[7][88] ), .CI(\SUMB[7][89] ), 
        .CO(\CARRYB[8][88] ), .S(\SUMB[8][88] ) );
  FA1A S2_7_88 ( .A(\ab[7][88] ), .B(\CARRYB[6][88] ), .CI(\SUMB[6][89] ), 
        .CO(\CARRYB[7][88] ), .S(\SUMB[7][88] ) );
  FA1A S2_6_88 ( .A(\ab[6][88] ), .B(\CARRYB[5][88] ), .CI(\SUMB[5][89] ), 
        .CO(\CARRYB[6][88] ), .S(\SUMB[6][88] ) );
  FA1A S2_5_88 ( .A(\ab[5][88] ), .B(\CARRYB[4][88] ), .CI(\SUMB[4][89] ), 
        .CO(\CARRYB[5][88] ), .S(\SUMB[5][88] ) );
  FA1A S2_4_88 ( .A(\ab[4][88] ), .B(\CARRYB[3][88] ), .CI(\SUMB[3][89] ), 
        .CO(\CARRYB[4][88] ), .S(\SUMB[4][88] ) );
  FA1A S2_3_88 ( .A(\ab[3][88] ), .B(\CARRYB[2][88] ), .CI(\SUMB[2][89] ), 
        .CO(\CARRYB[3][88] ), .S(\SUMB[3][88] ) );
  FA1A S2_2_88 ( .A(\ab[2][88] ), .B(\CARRYB[1][88] ), .CI(\SUMB[1][89] ), 
        .CO(\CARRYB[2][88] ), .S(\SUMB[2][88] ) );
  FA1A S2_14_87 ( .A(\ab[14][87] ), .B(\CARRYB[13][87] ), .CI(\SUMB[13][88] ), 
        .CO(\CARRYB[14][87] ), .S(\SUMB[14][87] ) );
  FA1A S2_13_87 ( .A(\ab[13][87] ), .B(\CARRYB[12][87] ), .CI(\SUMB[12][88] ), 
        .CO(\CARRYB[13][87] ), .S(\SUMB[13][87] ) );
  FA1A S2_12_87 ( .A(\ab[12][87] ), .B(\CARRYB[11][87] ), .CI(\SUMB[11][88] ), 
        .CO(\CARRYB[12][87] ), .S(\SUMB[12][87] ) );
  FA1A S2_11_87 ( .A(\ab[11][87] ), .B(\CARRYB[10][87] ), .CI(\SUMB[10][88] ), 
        .CO(\CARRYB[11][87] ), .S(\SUMB[11][87] ) );
  FA1A S2_10_87 ( .A(\ab[10][87] ), .B(\CARRYB[9][87] ), .CI(\SUMB[9][88] ), 
        .CO(\CARRYB[10][87] ), .S(\SUMB[10][87] ) );
  FA1A S2_9_87 ( .A(\ab[9][87] ), .B(\CARRYB[8][87] ), .CI(\SUMB[8][88] ), 
        .CO(\CARRYB[9][87] ), .S(\SUMB[9][87] ) );
  FA1A S2_8_87 ( .A(\ab[8][87] ), .B(\CARRYB[7][87] ), .CI(\SUMB[7][88] ), 
        .CO(\CARRYB[8][87] ), .S(\SUMB[8][87] ) );
  FA1A S2_7_87 ( .A(\ab[7][87] ), .B(\CARRYB[6][87] ), .CI(\SUMB[6][88] ), 
        .CO(\CARRYB[7][87] ), .S(\SUMB[7][87] ) );
  FA1A S2_6_87 ( .A(\ab[6][87] ), .B(\CARRYB[5][87] ), .CI(\SUMB[5][88] ), 
        .CO(\CARRYB[6][87] ), .S(\SUMB[6][87] ) );
  FA1A S2_5_87 ( .A(\ab[5][87] ), .B(\CARRYB[4][87] ), .CI(\SUMB[4][88] ), 
        .CO(\CARRYB[5][87] ), .S(\SUMB[5][87] ) );
  FA1A S2_4_87 ( .A(\ab[4][87] ), .B(\CARRYB[3][87] ), .CI(\SUMB[3][88] ), 
        .CO(\CARRYB[4][87] ), .S(\SUMB[4][87] ) );
  FA1A S2_3_87 ( .A(\ab[3][87] ), .B(\CARRYB[2][87] ), .CI(\SUMB[2][88] ), 
        .CO(\CARRYB[3][87] ), .S(\SUMB[3][87] ) );
  FA1A S2_2_87 ( .A(\ab[2][87] ), .B(\CARRYB[1][87] ), .CI(\SUMB[1][88] ), 
        .CO(\CARRYB[2][87] ), .S(\SUMB[2][87] ) );
  FA1A S2_14_86 ( .A(\ab[14][86] ), .B(\CARRYB[13][86] ), .CI(\SUMB[13][87] ), 
        .CO(\CARRYB[14][86] ), .S(\SUMB[14][86] ) );
  FA1A S2_13_86 ( .A(\ab[13][86] ), .B(\CARRYB[12][86] ), .CI(\SUMB[12][87] ), 
        .CO(\CARRYB[13][86] ), .S(\SUMB[13][86] ) );
  FA1A S2_12_86 ( .A(\ab[12][86] ), .B(\CARRYB[11][86] ), .CI(\SUMB[11][87] ), 
        .CO(\CARRYB[12][86] ), .S(\SUMB[12][86] ) );
  FA1A S2_11_86 ( .A(\ab[11][86] ), .B(\CARRYB[10][86] ), .CI(\SUMB[10][87] ), 
        .CO(\CARRYB[11][86] ), .S(\SUMB[11][86] ) );
  FA1A S2_10_86 ( .A(\ab[10][86] ), .B(\CARRYB[9][86] ), .CI(\SUMB[9][87] ), 
        .CO(\CARRYB[10][86] ), .S(\SUMB[10][86] ) );
  FA1A S2_9_86 ( .A(\ab[9][86] ), .B(\CARRYB[8][86] ), .CI(\SUMB[8][87] ), 
        .CO(\CARRYB[9][86] ), .S(\SUMB[9][86] ) );
  FA1A S2_8_86 ( .A(\ab[8][86] ), .B(\CARRYB[7][86] ), .CI(\SUMB[7][87] ), 
        .CO(\CARRYB[8][86] ), .S(\SUMB[8][86] ) );
  FA1A S2_7_86 ( .A(\ab[7][86] ), .B(\CARRYB[6][86] ), .CI(\SUMB[6][87] ), 
        .CO(\CARRYB[7][86] ), .S(\SUMB[7][86] ) );
  FA1A S2_6_86 ( .A(\ab[6][86] ), .B(\CARRYB[5][86] ), .CI(\SUMB[5][87] ), 
        .CO(\CARRYB[6][86] ), .S(\SUMB[6][86] ) );
  FA1A S2_5_86 ( .A(\ab[5][86] ), .B(\CARRYB[4][86] ), .CI(\SUMB[4][87] ), 
        .CO(\CARRYB[5][86] ), .S(\SUMB[5][86] ) );
  FA1A S2_4_86 ( .A(\ab[4][86] ), .B(\CARRYB[3][86] ), .CI(\SUMB[3][87] ), 
        .CO(\CARRYB[4][86] ), .S(\SUMB[4][86] ) );
  FA1A S2_3_86 ( .A(\ab[3][86] ), .B(\CARRYB[2][86] ), .CI(\SUMB[2][87] ), 
        .CO(\CARRYB[3][86] ), .S(\SUMB[3][86] ) );
  FA1A S2_2_86 ( .A(\ab[2][86] ), .B(\CARRYB[1][86] ), .CI(\SUMB[1][87] ), 
        .CO(\CARRYB[2][86] ), .S(\SUMB[2][86] ) );
  FA1A S2_14_85 ( .A(\ab[14][85] ), .B(\CARRYB[13][85] ), .CI(\SUMB[13][86] ), 
        .CO(\CARRYB[14][85] ), .S(\SUMB[14][85] ) );
  FA1A S2_13_85 ( .A(\ab[13][85] ), .B(\CARRYB[12][85] ), .CI(\SUMB[12][86] ), 
        .CO(\CARRYB[13][85] ), .S(\SUMB[13][85] ) );
  FA1A S2_12_85 ( .A(\ab[12][85] ), .B(\CARRYB[11][85] ), .CI(\SUMB[11][86] ), 
        .CO(\CARRYB[12][85] ), .S(\SUMB[12][85] ) );
  FA1A S2_11_85 ( .A(\ab[11][85] ), .B(\CARRYB[10][85] ), .CI(\SUMB[10][86] ), 
        .CO(\CARRYB[11][85] ), .S(\SUMB[11][85] ) );
  FA1A S2_10_85 ( .A(\ab[10][85] ), .B(\CARRYB[9][85] ), .CI(\SUMB[9][86] ), 
        .CO(\CARRYB[10][85] ), .S(\SUMB[10][85] ) );
  FA1A S2_9_85 ( .A(\ab[9][85] ), .B(\CARRYB[8][85] ), .CI(\SUMB[8][86] ), 
        .CO(\CARRYB[9][85] ), .S(\SUMB[9][85] ) );
  FA1A S2_8_85 ( .A(\ab[8][85] ), .B(\CARRYB[7][85] ), .CI(\SUMB[7][86] ), 
        .CO(\CARRYB[8][85] ), .S(\SUMB[8][85] ) );
  FA1A S2_7_85 ( .A(\ab[7][85] ), .B(\CARRYB[6][85] ), .CI(\SUMB[6][86] ), 
        .CO(\CARRYB[7][85] ), .S(\SUMB[7][85] ) );
  FA1A S2_6_85 ( .A(\ab[6][85] ), .B(\CARRYB[5][85] ), .CI(\SUMB[5][86] ), 
        .CO(\CARRYB[6][85] ), .S(\SUMB[6][85] ) );
  FA1A S2_5_85 ( .A(\ab[5][85] ), .B(\CARRYB[4][85] ), .CI(\SUMB[4][86] ), 
        .CO(\CARRYB[5][85] ), .S(\SUMB[5][85] ) );
  FA1A S2_4_85 ( .A(\ab[4][85] ), .B(\CARRYB[3][85] ), .CI(\SUMB[3][86] ), 
        .CO(\CARRYB[4][85] ), .S(\SUMB[4][85] ) );
  FA1A S2_3_85 ( .A(\ab[3][85] ), .B(\CARRYB[2][85] ), .CI(\SUMB[2][86] ), 
        .CO(\CARRYB[3][85] ), .S(\SUMB[3][85] ) );
  FA1A S2_2_85 ( .A(\ab[2][85] ), .B(\CARRYB[1][85] ), .CI(\SUMB[1][86] ), 
        .CO(\CARRYB[2][85] ), .S(\SUMB[2][85] ) );
  FA1A S2_14_81 ( .A(\ab[14][81] ), .B(\CARRYB[13][81] ), .CI(\SUMB[13][82] ), 
        .CO(\CARRYB[14][81] ), .S(\SUMB[14][81] ) );
  FA1A S2_13_81 ( .A(\ab[13][81] ), .B(\CARRYB[12][81] ), .CI(\SUMB[12][82] ), 
        .CO(\CARRYB[13][81] ), .S(\SUMB[13][81] ) );
  FA1A S2_12_81 ( .A(\ab[12][81] ), .B(\CARRYB[11][81] ), .CI(\SUMB[11][82] ), 
        .CO(\CARRYB[12][81] ), .S(\SUMB[12][81] ) );
  FA1A S2_11_81 ( .A(\ab[11][81] ), .B(\CARRYB[10][81] ), .CI(\SUMB[10][82] ), 
        .CO(\CARRYB[11][81] ), .S(\SUMB[11][81] ) );
  FA1A S2_10_81 ( .A(\ab[10][81] ), .B(\CARRYB[9][81] ), .CI(\SUMB[9][82] ), 
        .CO(\CARRYB[10][81] ), .S(\SUMB[10][81] ) );
  FA1A S2_9_81 ( .A(\ab[9][81] ), .B(\CARRYB[8][81] ), .CI(\SUMB[8][82] ), 
        .CO(\CARRYB[9][81] ), .S(\SUMB[9][81] ) );
  FA1A S2_8_81 ( .A(\ab[8][81] ), .B(\CARRYB[7][81] ), .CI(\SUMB[7][82] ), 
        .CO(\CARRYB[8][81] ), .S(\SUMB[8][81] ) );
  FA1A S2_7_81 ( .A(\ab[7][81] ), .B(\CARRYB[6][81] ), .CI(\SUMB[6][82] ), 
        .CO(\CARRYB[7][81] ), .S(\SUMB[7][81] ) );
  FA1A S2_6_81 ( .A(\ab[6][81] ), .B(\CARRYB[5][81] ), .CI(\SUMB[5][82] ), 
        .CO(\CARRYB[6][81] ), .S(\SUMB[6][81] ) );
  FA1A S2_5_81 ( .A(\ab[5][81] ), .B(\CARRYB[4][81] ), .CI(\SUMB[4][82] ), 
        .CO(\CARRYB[5][81] ), .S(\SUMB[5][81] ) );
  FA1A S2_4_81 ( .A(\ab[4][81] ), .B(\CARRYB[3][81] ), .CI(\SUMB[3][82] ), 
        .CO(\CARRYB[4][81] ), .S(\SUMB[4][81] ) );
  FA1A S2_3_81 ( .A(\ab[3][81] ), .B(\CARRYB[2][81] ), .CI(\SUMB[2][82] ), 
        .CO(\CARRYB[3][81] ), .S(\SUMB[3][81] ) );
  FA1A S2_2_81 ( .A(\ab[2][81] ), .B(\CARRYB[1][81] ), .CI(\SUMB[1][82] ), 
        .CO(\CARRYB[2][81] ), .S(\SUMB[2][81] ) );
  FA1A S2_14_84 ( .A(\ab[14][84] ), .B(\CARRYB[13][84] ), .CI(\SUMB[13][85] ), 
        .CO(\CARRYB[14][84] ), .S(\SUMB[14][84] ) );
  FA1A S2_14_83 ( .A(\ab[14][83] ), .B(\CARRYB[13][83] ), .CI(\SUMB[13][84] ), 
        .CO(\CARRYB[14][83] ), .S(\SUMB[14][83] ) );
  FA1A S2_13_84 ( .A(\ab[13][84] ), .B(\CARRYB[12][84] ), .CI(\SUMB[12][85] ), 
        .CO(\CARRYB[13][84] ), .S(\SUMB[13][84] ) );
  FA1A S2_14_80 ( .A(\ab[14][80] ), .B(\CARRYB[13][80] ), .CI(\SUMB[13][81] ), 
        .CO(\CARRYB[14][80] ), .S(\SUMB[14][80] ) );
  FA1A S2_14_82 ( .A(\ab[14][82] ), .B(\CARRYB[13][82] ), .CI(\SUMB[13][83] ), 
        .CO(\CARRYB[14][82] ), .S(\SUMB[14][82] ) );
  FA1A S2_13_80 ( .A(\ab[13][80] ), .B(\CARRYB[12][80] ), .CI(\SUMB[12][81] ), 
        .CO(\CARRYB[13][80] ), .S(\SUMB[13][80] ) );
  FA1A S2_13_82 ( .A(\ab[13][82] ), .B(\CARRYB[12][82] ), .CI(\SUMB[12][83] ), 
        .CO(\CARRYB[13][82] ), .S(\SUMB[13][82] ) );
  FA1A S2_13_83 ( .A(\ab[13][83] ), .B(\CARRYB[12][83] ), .CI(\SUMB[12][84] ), 
        .CO(\CARRYB[13][83] ), .S(\SUMB[13][83] ) );
  FA1A S2_12_80 ( .A(\ab[12][80] ), .B(\CARRYB[11][80] ), .CI(\SUMB[11][81] ), 
        .CO(\CARRYB[12][80] ), .S(\SUMB[12][80] ) );
  FA1A S2_12_82 ( .A(\ab[12][82] ), .B(\CARRYB[11][82] ), .CI(\SUMB[11][83] ), 
        .CO(\CARRYB[12][82] ), .S(\SUMB[12][82] ) );
  FA1A S2_12_83 ( .A(\ab[12][83] ), .B(\CARRYB[11][83] ), .CI(\SUMB[11][84] ), 
        .CO(\CARRYB[12][83] ), .S(\SUMB[12][83] ) );
  FA1A S2_12_84 ( .A(\ab[12][84] ), .B(\CARRYB[11][84] ), .CI(\SUMB[11][85] ), 
        .CO(\CARRYB[12][84] ), .S(\SUMB[12][84] ) );
  FA1A S2_11_82 ( .A(\ab[11][82] ), .B(\CARRYB[10][82] ), .CI(\SUMB[10][83] ), 
        .CO(\CARRYB[11][82] ), .S(\SUMB[11][82] ) );
  FA1A S2_11_83 ( .A(\ab[11][83] ), .B(\CARRYB[10][83] ), .CI(\SUMB[10][84] ), 
        .CO(\CARRYB[11][83] ), .S(\SUMB[11][83] ) );
  FA1A S2_11_84 ( .A(\ab[11][84] ), .B(\CARRYB[10][84] ), .CI(\SUMB[10][85] ), 
        .CO(\CARRYB[11][84] ), .S(\SUMB[11][84] ) );
  FA1A S2_10_82 ( .A(\ab[10][82] ), .B(\CARRYB[9][82] ), .CI(\SUMB[9][83] ), 
        .CO(\CARRYB[10][82] ), .S(\SUMB[10][82] ) );
  FA1A S2_10_83 ( .A(\ab[10][83] ), .B(\CARRYB[9][83] ), .CI(\SUMB[9][84] ), 
        .CO(\CARRYB[10][83] ), .S(\SUMB[10][83] ) );
  FA1A S2_10_84 ( .A(\ab[10][84] ), .B(\CARRYB[9][84] ), .CI(\SUMB[9][85] ), 
        .CO(\CARRYB[10][84] ), .S(\SUMB[10][84] ) );
  FA1A S2_9_83 ( .A(\ab[9][83] ), .B(\CARRYB[8][83] ), .CI(\SUMB[8][84] ), 
        .CO(\CARRYB[9][83] ), .S(\SUMB[9][83] ) );
  FA1A S2_9_84 ( .A(\ab[9][84] ), .B(\CARRYB[8][84] ), .CI(\SUMB[8][85] ), 
        .CO(\CARRYB[9][84] ), .S(\SUMB[9][84] ) );
  FA1A S2_11_80 ( .A(\ab[11][80] ), .B(\CARRYB[10][80] ), .CI(\SUMB[10][81] ), 
        .CO(\CARRYB[11][80] ), .S(\SUMB[11][80] ) );
  FA1A S2_8_84 ( .A(\ab[8][84] ), .B(\CARRYB[7][84] ), .CI(\SUMB[7][85] ), 
        .CO(\CARRYB[8][84] ), .S(\SUMB[8][84] ) );
  FA1A S2_10_80 ( .A(\ab[10][80] ), .B(\CARRYB[9][80] ), .CI(\SUMB[9][81] ), 
        .CO(\CARRYB[10][80] ), .S(\SUMB[10][80] ) );
  FA1A S2_9_80 ( .A(\ab[9][80] ), .B(\CARRYB[8][80] ), .CI(\SUMB[8][81] ), 
        .CO(\CARRYB[9][80] ), .S(\SUMB[9][80] ) );
  FA1A S2_9_82 ( .A(\ab[9][82] ), .B(\CARRYB[8][82] ), .CI(\SUMB[8][83] ), 
        .CO(\CARRYB[9][82] ), .S(\SUMB[9][82] ) );
  FA1A S2_8_80 ( .A(\ab[8][80] ), .B(\CARRYB[7][80] ), .CI(\SUMB[7][81] ), 
        .CO(\CARRYB[8][80] ), .S(\SUMB[8][80] ) );
  FA1A S2_8_82 ( .A(\ab[8][82] ), .B(\CARRYB[7][82] ), .CI(\SUMB[7][83] ), 
        .CO(\CARRYB[8][82] ), .S(\SUMB[8][82] ) );
  FA1A S2_8_83 ( .A(\ab[8][83] ), .B(\CARRYB[7][83] ), .CI(\SUMB[7][84] ), 
        .CO(\CARRYB[8][83] ), .S(\SUMB[8][83] ) );
  FA1A S2_7_82 ( .A(\ab[7][82] ), .B(\CARRYB[6][82] ), .CI(\SUMB[6][83] ), 
        .CO(\CARRYB[7][82] ), .S(\SUMB[7][82] ) );
  FA1A S2_7_80 ( .A(\ab[7][80] ), .B(\CARRYB[6][80] ), .CI(\SUMB[6][81] ), 
        .CO(\CARRYB[7][80] ), .S(\SUMB[7][80] ) );
  FA1A S2_7_83 ( .A(\ab[7][83] ), .B(\CARRYB[6][83] ), .CI(\SUMB[6][84] ), 
        .CO(\CARRYB[7][83] ), .S(\SUMB[7][83] ) );
  FA1A S2_7_84 ( .A(\ab[7][84] ), .B(\CARRYB[6][84] ), .CI(\SUMB[6][85] ), 
        .CO(\CARRYB[7][84] ), .S(\SUMB[7][84] ) );
  FA1A S2_6_83 ( .A(\ab[6][83] ), .B(\CARRYB[5][83] ), .CI(\SUMB[5][84] ), 
        .CO(\CARRYB[6][83] ), .S(\SUMB[6][83] ) );
  FA1A S2_6_82 ( .A(\ab[6][82] ), .B(\CARRYB[5][82] ), .CI(\SUMB[5][83] ), 
        .CO(\CARRYB[6][82] ), .S(\SUMB[6][82] ) );
  FA1A S2_6_80 ( .A(\ab[6][80] ), .B(\CARRYB[5][80] ), .CI(\SUMB[5][81] ), 
        .CO(\CARRYB[6][80] ), .S(\SUMB[6][80] ) );
  FA1A S2_6_84 ( .A(\ab[6][84] ), .B(\CARRYB[5][84] ), .CI(\SUMB[5][85] ), 
        .CO(\CARRYB[6][84] ), .S(\SUMB[6][84] ) );
  FA1A S2_5_84 ( .A(\ab[5][84] ), .B(\CARRYB[4][84] ), .CI(\SUMB[4][85] ), 
        .CO(\CARRYB[5][84] ), .S(\SUMB[5][84] ) );
  FA1A S2_5_83 ( .A(\ab[5][83] ), .B(\CARRYB[4][83] ), .CI(\SUMB[4][84] ), 
        .CO(\CARRYB[5][83] ), .S(\SUMB[5][83] ) );
  FA1A S2_5_82 ( .A(\ab[5][82] ), .B(\CARRYB[4][82] ), .CI(\SUMB[4][83] ), 
        .CO(\CARRYB[5][82] ), .S(\SUMB[5][82] ) );
  FA1A S2_5_80 ( .A(\ab[5][80] ), .B(\CARRYB[4][80] ), .CI(\SUMB[4][81] ), 
        .CO(\CARRYB[5][80] ), .S(\SUMB[5][80] ) );
  FA1A S2_4_84 ( .A(\ab[4][84] ), .B(\CARRYB[3][84] ), .CI(\SUMB[3][85] ), 
        .CO(\CARRYB[4][84] ), .S(\SUMB[4][84] ) );
  FA1A S2_4_83 ( .A(\ab[4][83] ), .B(\CARRYB[3][83] ), .CI(\SUMB[3][84] ), 
        .CO(\CARRYB[4][83] ), .S(\SUMB[4][83] ) );
  FA1A S2_4_82 ( .A(\ab[4][82] ), .B(\CARRYB[3][82] ), .CI(\SUMB[3][83] ), 
        .CO(\CARRYB[4][82] ), .S(\SUMB[4][82] ) );
  FA1A S2_4_80 ( .A(\ab[4][80] ), .B(\CARRYB[3][80] ), .CI(\SUMB[3][81] ), 
        .CO(\CARRYB[4][80] ), .S(\SUMB[4][80] ) );
  FA1A S2_3_84 ( .A(\ab[3][84] ), .B(\CARRYB[2][84] ), .CI(\SUMB[2][85] ), 
        .CO(\CARRYB[3][84] ), .S(\SUMB[3][84] ) );
  FA1A S2_3_83 ( .A(\ab[3][83] ), .B(\CARRYB[2][83] ), .CI(\SUMB[2][84] ), 
        .CO(\CARRYB[3][83] ), .S(\SUMB[3][83] ) );
  FA1A S2_3_82 ( .A(\ab[3][82] ), .B(\CARRYB[2][82] ), .CI(\SUMB[2][83] ), 
        .CO(\CARRYB[3][82] ), .S(\SUMB[3][82] ) );
  FA1A S2_3_80 ( .A(\ab[3][80] ), .B(\CARRYB[2][80] ), .CI(\SUMB[2][81] ), 
        .CO(\CARRYB[3][80] ), .S(\SUMB[3][80] ) );
  FA1A S2_2_84 ( .A(\ab[2][84] ), .B(\CARRYB[1][84] ), .CI(\SUMB[1][85] ), 
        .CO(\CARRYB[2][84] ), .S(\SUMB[2][84] ) );
  FA1A S2_2_83 ( .A(\ab[2][83] ), .B(\CARRYB[1][83] ), .CI(\SUMB[1][84] ), 
        .CO(\CARRYB[2][83] ), .S(\SUMB[2][83] ) );
  FA1A S2_2_82 ( .A(\ab[2][82] ), .B(\CARRYB[1][82] ), .CI(\SUMB[1][83] ), 
        .CO(\CARRYB[2][82] ), .S(\SUMB[2][82] ) );
  FA1A S2_2_80 ( .A(\ab[2][80] ), .B(\CARRYB[1][80] ), .CI(\SUMB[1][81] ), 
        .CO(\CARRYB[2][80] ), .S(\SUMB[2][80] ) );
  FA1A S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FA1A S4_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), .CO(
        \CARRYB[29][0] ), .S(\SUMB[29][0] ) );
  FA1A S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FA1A S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FA1A S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(\A1[22] ) );
  FA1A S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FA1A S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA1A S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\A1[21] ) );
  FA1A S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA1A S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FA1A S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA1A S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA1A S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA1A S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S2_14_78 ( .A(\ab[14][78] ), .B(\CARRYB[13][78] ), .CI(\SUMB[13][79] ), 
        .CO(\CARRYB[14][78] ), .S(\SUMB[14][78] ) );
  FA1A S2_14_79 ( .A(\ab[14][79] ), .B(\CARRYB[13][79] ), .CI(\SUMB[13][80] ), 
        .CO(\CARRYB[14][79] ), .S(\SUMB[14][79] ) );
  FA1A S2_13_79 ( .A(\ab[13][79] ), .B(\CARRYB[12][79] ), .CI(\SUMB[12][80] ), 
        .CO(\CARRYB[13][79] ), .S(\SUMB[13][79] ) );
  FA1A S2_14_75 ( .A(\ab[14][75] ), .B(\CARRYB[13][75] ), .CI(\SUMB[13][76] ), 
        .CO(\CARRYB[14][75] ), .S(\SUMB[14][75] ) );
  FA1A S2_14_74 ( .A(\ab[14][74] ), .B(\CARRYB[13][74] ), .CI(\SUMB[13][75] ), 
        .CO(\CARRYB[14][74] ), .S(\SUMB[14][74] ) );
  FA1A S2_14_73 ( .A(\ab[14][73] ), .B(\CARRYB[13][73] ), .CI(\SUMB[13][74] ), 
        .CO(\CARRYB[14][73] ), .S(\SUMB[14][73] ) );
  FA1A S2_14_72 ( .A(\ab[14][72] ), .B(\CARRYB[13][72] ), .CI(\SUMB[13][73] ), 
        .CO(\CARRYB[14][72] ), .S(\SUMB[14][72] ) );
  FA1A S2_14_71 ( .A(\ab[14][71] ), .B(\CARRYB[13][71] ), .CI(\SUMB[13][72] ), 
        .CO(\CARRYB[14][71] ), .S(\SUMB[14][71] ) );
  FA1A S2_14_70 ( .A(\ab[14][70] ), .B(\CARRYB[13][70] ), .CI(\SUMB[13][71] ), 
        .CO(\CARRYB[14][70] ), .S(\SUMB[14][70] ) );
  FA1A S2_14_69 ( .A(\ab[14][69] ), .B(\CARRYB[13][69] ), .CI(\SUMB[13][70] ), 
        .CO(\CARRYB[14][69] ), .S(\SUMB[14][69] ) );
  FA1A S2_14_76 ( .A(\ab[14][76] ), .B(\CARRYB[13][76] ), .CI(\SUMB[13][77] ), 
        .CO(\CARRYB[14][76] ), .S(\SUMB[14][76] ) );
  FA1A S2_14_77 ( .A(\ab[14][77] ), .B(\CARRYB[13][77] ), .CI(\SUMB[13][78] ), 
        .CO(\CARRYB[14][77] ), .S(\SUMB[14][77] ) );
  FA1A S2_13_76 ( .A(\ab[13][76] ), .B(\CARRYB[12][76] ), .CI(\SUMB[12][77] ), 
        .CO(\CARRYB[13][76] ), .S(\SUMB[13][76] ) );
  FA1A S2_13_75 ( .A(\ab[13][75] ), .B(\CARRYB[12][75] ), .CI(\SUMB[12][76] ), 
        .CO(\CARRYB[13][75] ), .S(\SUMB[13][75] ) );
  FA1A S2_13_74 ( .A(\ab[13][74] ), .B(\CARRYB[12][74] ), .CI(\SUMB[12][75] ), 
        .CO(\CARRYB[13][74] ), .S(\SUMB[13][74] ) );
  FA1A S2_13_73 ( .A(\ab[13][73] ), .B(\CARRYB[12][73] ), .CI(\SUMB[12][74] ), 
        .CO(\CARRYB[13][73] ), .S(\SUMB[13][73] ) );
  FA1A S2_13_72 ( .A(\ab[13][72] ), .B(\CARRYB[12][72] ), .CI(\SUMB[12][73] ), 
        .CO(\CARRYB[13][72] ), .S(\SUMB[13][72] ) );
  FA1A S2_13_71 ( .A(\ab[13][71] ), .B(\CARRYB[12][71] ), .CI(\SUMB[12][72] ), 
        .CO(\CARRYB[13][71] ), .S(\SUMB[13][71] ) );
  FA1A S2_13_70 ( .A(\ab[13][70] ), .B(\CARRYB[12][70] ), .CI(\SUMB[12][71] ), 
        .CO(\CARRYB[13][70] ), .S(\SUMB[13][70] ) );
  FA1A S2_13_69 ( .A(\ab[13][69] ), .B(\CARRYB[12][69] ), .CI(\SUMB[12][70] ), 
        .CO(\CARRYB[13][69] ), .S(\SUMB[13][69] ) );
  FA1A S2_13_77 ( .A(\ab[13][77] ), .B(\CARRYB[12][77] ), .CI(\SUMB[12][78] ), 
        .CO(\CARRYB[13][77] ), .S(\SUMB[13][77] ) );
  FA1A S2_13_78 ( .A(\ab[13][78] ), .B(\CARRYB[12][78] ), .CI(\SUMB[12][79] ), 
        .CO(\CARRYB[13][78] ), .S(\SUMB[13][78] ) );
  FA1A S2_12_77 ( .A(\ab[12][77] ), .B(\CARRYB[11][77] ), .CI(\SUMB[11][78] ), 
        .CO(\CARRYB[12][77] ), .S(\SUMB[12][77] ) );
  FA1A S2_12_76 ( .A(\ab[12][76] ), .B(\CARRYB[11][76] ), .CI(\SUMB[11][77] ), 
        .CO(\CARRYB[12][76] ), .S(\SUMB[12][76] ) );
  FA1A S2_12_75 ( .A(\ab[12][75] ), .B(\CARRYB[11][75] ), .CI(\SUMB[11][76] ), 
        .CO(\CARRYB[12][75] ), .S(\SUMB[12][75] ) );
  FA1A S2_12_74 ( .A(\ab[12][74] ), .B(\CARRYB[11][74] ), .CI(\SUMB[11][75] ), 
        .CO(\CARRYB[12][74] ), .S(\SUMB[12][74] ) );
  FA1A S2_12_73 ( .A(\ab[12][73] ), .B(\CARRYB[11][73] ), .CI(\SUMB[11][74] ), 
        .CO(\CARRYB[12][73] ), .S(\SUMB[12][73] ) );
  FA1A S2_12_72 ( .A(\ab[12][72] ), .B(\CARRYB[11][72] ), .CI(\SUMB[11][73] ), 
        .CO(\CARRYB[12][72] ), .S(\SUMB[12][72] ) );
  FA1A S2_12_71 ( .A(\ab[12][71] ), .B(\CARRYB[11][71] ), .CI(\SUMB[11][72] ), 
        .CO(\CARRYB[12][71] ), .S(\SUMB[12][71] ) );
  FA1A S2_12_70 ( .A(\ab[12][70] ), .B(\CARRYB[11][70] ), .CI(\SUMB[11][71] ), 
        .CO(\CARRYB[12][70] ), .S(\SUMB[12][70] ) );
  FA1A S2_12_69 ( .A(\ab[12][69] ), .B(\CARRYB[11][69] ), .CI(\SUMB[11][70] ), 
        .CO(\CARRYB[12][69] ), .S(\SUMB[12][69] ) );
  FA1A S2_12_78 ( .A(\ab[12][78] ), .B(\CARRYB[11][78] ), .CI(\SUMB[11][79] ), 
        .CO(\CARRYB[12][78] ), .S(\SUMB[12][78] ) );
  FA1A S2_12_79 ( .A(\ab[12][79] ), .B(\CARRYB[11][79] ), .CI(\SUMB[11][80] ), 
        .CO(\CARRYB[12][79] ), .S(\SUMB[12][79] ) );
  FA1A S2_11_78 ( .A(\ab[11][78] ), .B(\CARRYB[10][78] ), .CI(\SUMB[10][79] ), 
        .CO(\CARRYB[11][78] ), .S(\SUMB[11][78] ) );
  FA1A S2_11_77 ( .A(\ab[11][77] ), .B(\CARRYB[10][77] ), .CI(\SUMB[10][78] ), 
        .CO(\CARRYB[11][77] ), .S(\SUMB[11][77] ) );
  FA1A S2_11_76 ( .A(\ab[11][76] ), .B(\CARRYB[10][76] ), .CI(\SUMB[10][77] ), 
        .CO(\CARRYB[11][76] ), .S(\SUMB[11][76] ) );
  FA1A S2_11_75 ( .A(\ab[11][75] ), .B(\CARRYB[10][75] ), .CI(\SUMB[10][76] ), 
        .CO(\CARRYB[11][75] ), .S(\SUMB[11][75] ) );
  FA1A S2_11_74 ( .A(\ab[11][74] ), .B(\CARRYB[10][74] ), .CI(\SUMB[10][75] ), 
        .CO(\CARRYB[11][74] ), .S(\SUMB[11][74] ) );
  FA1A S2_11_73 ( .A(\ab[11][73] ), .B(\CARRYB[10][73] ), .CI(\SUMB[10][74] ), 
        .CO(\CARRYB[11][73] ), .S(\SUMB[11][73] ) );
  FA1A S2_11_72 ( .A(\ab[11][72] ), .B(\CARRYB[10][72] ), .CI(\SUMB[10][73] ), 
        .CO(\CARRYB[11][72] ), .S(\SUMB[11][72] ) );
  FA1A S2_11_71 ( .A(\ab[11][71] ), .B(\CARRYB[10][71] ), .CI(\SUMB[10][72] ), 
        .CO(\CARRYB[11][71] ), .S(\SUMB[11][71] ) );
  FA1A S2_11_70 ( .A(\ab[11][70] ), .B(\CARRYB[10][70] ), .CI(\SUMB[10][71] ), 
        .CO(\CARRYB[11][70] ), .S(\SUMB[11][70] ) );
  FA1A S2_11_69 ( .A(\ab[11][69] ), .B(\CARRYB[10][69] ), .CI(\SUMB[10][70] ), 
        .CO(\CARRYB[11][69] ), .S(\SUMB[11][69] ) );
  FA1A S2_11_79 ( .A(\ab[11][79] ), .B(\CARRYB[10][79] ), .CI(\SUMB[10][80] ), 
        .CO(\CARRYB[11][79] ), .S(\SUMB[11][79] ) );
  FA1A S2_10_79 ( .A(\ab[10][79] ), .B(\CARRYB[9][79] ), .CI(\SUMB[9][80] ), 
        .CO(\CARRYB[10][79] ), .S(\SUMB[10][79] ) );
  FA1A S2_10_78 ( .A(\ab[10][78] ), .B(\CARRYB[9][78] ), .CI(\SUMB[9][79] ), 
        .CO(\CARRYB[10][78] ), .S(\SUMB[10][78] ) );
  FA1A S2_10_77 ( .A(\ab[10][77] ), .B(\CARRYB[9][77] ), .CI(\SUMB[9][78] ), 
        .CO(\CARRYB[10][77] ), .S(\SUMB[10][77] ) );
  FA1A S2_10_76 ( .A(\ab[10][76] ), .B(\CARRYB[9][76] ), .CI(\SUMB[9][77] ), 
        .CO(\CARRYB[10][76] ), .S(\SUMB[10][76] ) );
  FA1A S2_10_75 ( .A(\ab[10][75] ), .B(\CARRYB[9][75] ), .CI(\SUMB[9][76] ), 
        .CO(\CARRYB[10][75] ), .S(\SUMB[10][75] ) );
  FA1A S2_10_74 ( .A(\ab[10][74] ), .B(\CARRYB[9][74] ), .CI(\SUMB[9][75] ), 
        .CO(\CARRYB[10][74] ), .S(\SUMB[10][74] ) );
  FA1A S2_10_73 ( .A(\ab[10][73] ), .B(\CARRYB[9][73] ), .CI(\SUMB[9][74] ), 
        .CO(\CARRYB[10][73] ), .S(\SUMB[10][73] ) );
  FA1A S2_10_72 ( .A(\ab[10][72] ), .B(\CARRYB[9][72] ), .CI(\SUMB[9][73] ), 
        .CO(\CARRYB[10][72] ), .S(\SUMB[10][72] ) );
  FA1A S2_10_71 ( .A(\ab[10][71] ), .B(\CARRYB[9][71] ), .CI(\SUMB[9][72] ), 
        .CO(\CARRYB[10][71] ), .S(\SUMB[10][71] ) );
  FA1A S2_10_70 ( .A(\ab[10][70] ), .B(\CARRYB[9][70] ), .CI(\SUMB[9][71] ), 
        .CO(\CARRYB[10][70] ), .S(\SUMB[10][70] ) );
  FA1A S2_10_69 ( .A(\ab[10][69] ), .B(\CARRYB[9][69] ), .CI(\SUMB[9][70] ), 
        .CO(\CARRYB[10][69] ), .S(\SUMB[10][69] ) );
  FA1A S2_9_79 ( .A(\ab[9][79] ), .B(\CARRYB[8][79] ), .CI(\SUMB[8][80] ), 
        .CO(\CARRYB[9][79] ), .S(\SUMB[9][79] ) );
  FA1A S2_9_78 ( .A(\ab[9][78] ), .B(\CARRYB[8][78] ), .CI(\SUMB[8][79] ), 
        .CO(\CARRYB[9][78] ), .S(\SUMB[9][78] ) );
  FA1A S2_9_77 ( .A(\ab[9][77] ), .B(\CARRYB[8][77] ), .CI(\SUMB[8][78] ), 
        .CO(\CARRYB[9][77] ), .S(\SUMB[9][77] ) );
  FA1A S2_9_76 ( .A(\ab[9][76] ), .B(\CARRYB[8][76] ), .CI(\SUMB[8][77] ), 
        .CO(\CARRYB[9][76] ), .S(\SUMB[9][76] ) );
  FA1A S2_9_75 ( .A(\ab[9][75] ), .B(\CARRYB[8][75] ), .CI(\SUMB[8][76] ), 
        .CO(\CARRYB[9][75] ), .S(\SUMB[9][75] ) );
  FA1A S2_9_74 ( .A(\ab[9][74] ), .B(\CARRYB[8][74] ), .CI(\SUMB[8][75] ), 
        .CO(\CARRYB[9][74] ), .S(\SUMB[9][74] ) );
  FA1A S2_9_73 ( .A(\ab[9][73] ), .B(\CARRYB[8][73] ), .CI(\SUMB[8][74] ), 
        .CO(\CARRYB[9][73] ), .S(\SUMB[9][73] ) );
  FA1A S2_9_72 ( .A(\ab[9][72] ), .B(\CARRYB[8][72] ), .CI(\SUMB[8][73] ), 
        .CO(\CARRYB[9][72] ), .S(\SUMB[9][72] ) );
  FA1A S2_9_71 ( .A(\ab[9][71] ), .B(\CARRYB[8][71] ), .CI(\SUMB[8][72] ), 
        .CO(\CARRYB[9][71] ), .S(\SUMB[9][71] ) );
  FA1A S2_9_70 ( .A(\ab[9][70] ), .B(\CARRYB[8][70] ), .CI(\SUMB[8][71] ), 
        .CO(\CARRYB[9][70] ), .S(\SUMB[9][70] ) );
  FA1A S2_9_69 ( .A(\ab[9][69] ), .B(\CARRYB[8][69] ), .CI(\SUMB[8][70] ), 
        .CO(\CARRYB[9][69] ), .S(\SUMB[9][69] ) );
  FA1A S2_8_79 ( .A(\ab[8][79] ), .B(\CARRYB[7][79] ), .CI(\SUMB[7][80] ), 
        .CO(\CARRYB[8][79] ), .S(\SUMB[8][79] ) );
  FA1A S2_8_78 ( .A(\ab[8][78] ), .B(\CARRYB[7][78] ), .CI(\SUMB[7][79] ), 
        .CO(\CARRYB[8][78] ), .S(\SUMB[8][78] ) );
  FA1A S2_8_77 ( .A(\ab[8][77] ), .B(\CARRYB[7][77] ), .CI(\SUMB[7][78] ), 
        .CO(\CARRYB[8][77] ), .S(\SUMB[8][77] ) );
  FA1A S2_8_76 ( .A(\ab[8][76] ), .B(\CARRYB[7][76] ), .CI(\SUMB[7][77] ), 
        .CO(\CARRYB[8][76] ), .S(\SUMB[8][76] ) );
  FA1A S2_8_75 ( .A(\ab[8][75] ), .B(\CARRYB[7][75] ), .CI(\SUMB[7][76] ), 
        .CO(\CARRYB[8][75] ), .S(\SUMB[8][75] ) );
  FA1A S2_8_74 ( .A(\ab[8][74] ), .B(\CARRYB[7][74] ), .CI(\SUMB[7][75] ), 
        .CO(\CARRYB[8][74] ), .S(\SUMB[8][74] ) );
  FA1A S2_8_73 ( .A(\ab[8][73] ), .B(\CARRYB[7][73] ), .CI(\SUMB[7][74] ), 
        .CO(\CARRYB[8][73] ), .S(\SUMB[8][73] ) );
  FA1A S2_8_72 ( .A(\ab[8][72] ), .B(\CARRYB[7][72] ), .CI(\SUMB[7][73] ), 
        .CO(\CARRYB[8][72] ), .S(\SUMB[8][72] ) );
  FA1A S2_8_71 ( .A(\ab[8][71] ), .B(\CARRYB[7][71] ), .CI(\SUMB[7][72] ), 
        .CO(\CARRYB[8][71] ), .S(\SUMB[8][71] ) );
  FA1A S2_8_70 ( .A(\ab[8][70] ), .B(\CARRYB[7][70] ), .CI(\SUMB[7][71] ), 
        .CO(\CARRYB[8][70] ), .S(\SUMB[8][70] ) );
  FA1A S2_8_69 ( .A(\ab[8][69] ), .B(\CARRYB[7][69] ), .CI(\SUMB[7][70] ), 
        .CO(\CARRYB[8][69] ), .S(\SUMB[8][69] ) );
  FA1A S2_7_79 ( .A(\ab[7][79] ), .B(\CARRYB[6][79] ), .CI(\SUMB[6][80] ), 
        .CO(\CARRYB[7][79] ), .S(\SUMB[7][79] ) );
  FA1A S2_7_78 ( .A(\ab[7][78] ), .B(\CARRYB[6][78] ), .CI(\SUMB[6][79] ), 
        .CO(\CARRYB[7][78] ), .S(\SUMB[7][78] ) );
  FA1A S2_7_77 ( .A(\ab[7][77] ), .B(\CARRYB[6][77] ), .CI(\SUMB[6][78] ), 
        .CO(\CARRYB[7][77] ), .S(\SUMB[7][77] ) );
  FA1A S2_7_76 ( .A(\ab[7][76] ), .B(\CARRYB[6][76] ), .CI(\SUMB[6][77] ), 
        .CO(\CARRYB[7][76] ), .S(\SUMB[7][76] ) );
  FA1A S2_7_75 ( .A(\ab[7][75] ), .B(\CARRYB[6][75] ), .CI(\SUMB[6][76] ), 
        .CO(\CARRYB[7][75] ), .S(\SUMB[7][75] ) );
  FA1A S2_7_74 ( .A(\ab[7][74] ), .B(\CARRYB[6][74] ), .CI(\SUMB[6][75] ), 
        .CO(\CARRYB[7][74] ), .S(\SUMB[7][74] ) );
  FA1A S2_7_73 ( .A(\ab[7][73] ), .B(\CARRYB[6][73] ), .CI(\SUMB[6][74] ), 
        .CO(\CARRYB[7][73] ), .S(\SUMB[7][73] ) );
  FA1A S2_7_72 ( .A(\ab[7][72] ), .B(\CARRYB[6][72] ), .CI(\SUMB[6][73] ), 
        .CO(\CARRYB[7][72] ), .S(\SUMB[7][72] ) );
  FA1A S2_7_71 ( .A(\ab[7][71] ), .B(\CARRYB[6][71] ), .CI(\SUMB[6][72] ), 
        .CO(\CARRYB[7][71] ), .S(\SUMB[7][71] ) );
  FA1A S2_7_70 ( .A(\ab[7][70] ), .B(\CARRYB[6][70] ), .CI(\SUMB[6][71] ), 
        .CO(\CARRYB[7][70] ), .S(\SUMB[7][70] ) );
  FA1A S2_7_69 ( .A(\ab[7][69] ), .B(\CARRYB[6][69] ), .CI(\SUMB[6][70] ), 
        .CO(\CARRYB[7][69] ), .S(\SUMB[7][69] ) );
  FA1A S2_6_79 ( .A(\ab[6][79] ), .B(\CARRYB[5][79] ), .CI(\SUMB[5][80] ), 
        .CO(\CARRYB[6][79] ), .S(\SUMB[6][79] ) );
  FA1A S2_6_78 ( .A(\ab[6][78] ), .B(\CARRYB[5][78] ), .CI(\SUMB[5][79] ), 
        .CO(\CARRYB[6][78] ), .S(\SUMB[6][78] ) );
  FA1A S2_6_77 ( .A(\ab[6][77] ), .B(\CARRYB[5][77] ), .CI(\SUMB[5][78] ), 
        .CO(\CARRYB[6][77] ), .S(\SUMB[6][77] ) );
  FA1A S2_6_76 ( .A(\ab[6][76] ), .B(\CARRYB[5][76] ), .CI(\SUMB[5][77] ), 
        .CO(\CARRYB[6][76] ), .S(\SUMB[6][76] ) );
  FA1A S2_6_75 ( .A(\ab[6][75] ), .B(\CARRYB[5][75] ), .CI(\SUMB[5][76] ), 
        .CO(\CARRYB[6][75] ), .S(\SUMB[6][75] ) );
  FA1A S2_6_74 ( .A(\ab[6][74] ), .B(\CARRYB[5][74] ), .CI(\SUMB[5][75] ), 
        .CO(\CARRYB[6][74] ), .S(\SUMB[6][74] ) );
  FA1A S2_6_73 ( .A(\ab[6][73] ), .B(\CARRYB[5][73] ), .CI(\SUMB[5][74] ), 
        .CO(\CARRYB[6][73] ), .S(\SUMB[6][73] ) );
  FA1A S2_6_72 ( .A(\ab[6][72] ), .B(\CARRYB[5][72] ), .CI(\SUMB[5][73] ), 
        .CO(\CARRYB[6][72] ), .S(\SUMB[6][72] ) );
  FA1A S2_6_71 ( .A(\ab[6][71] ), .B(\CARRYB[5][71] ), .CI(\SUMB[5][72] ), 
        .CO(\CARRYB[6][71] ), .S(\SUMB[6][71] ) );
  FA1A S2_6_70 ( .A(\ab[6][70] ), .B(\CARRYB[5][70] ), .CI(\SUMB[5][71] ), 
        .CO(\CARRYB[6][70] ), .S(\SUMB[6][70] ) );
  FA1A S2_6_69 ( .A(\ab[6][69] ), .B(\CARRYB[5][69] ), .CI(\SUMB[5][70] ), 
        .CO(\CARRYB[6][69] ), .S(\SUMB[6][69] ) );
  FA1A S2_5_79 ( .A(\ab[5][79] ), .B(\CARRYB[4][79] ), .CI(\SUMB[4][80] ), 
        .CO(\CARRYB[5][79] ), .S(\SUMB[5][79] ) );
  FA1A S2_5_78 ( .A(\ab[5][78] ), .B(\CARRYB[4][78] ), .CI(\SUMB[4][79] ), 
        .CO(\CARRYB[5][78] ), .S(\SUMB[5][78] ) );
  FA1A S2_5_77 ( .A(\ab[5][77] ), .B(\CARRYB[4][77] ), .CI(\SUMB[4][78] ), 
        .CO(\CARRYB[5][77] ), .S(\SUMB[5][77] ) );
  FA1A S2_5_76 ( .A(\ab[5][76] ), .B(\CARRYB[4][76] ), .CI(\SUMB[4][77] ), 
        .CO(\CARRYB[5][76] ), .S(\SUMB[5][76] ) );
  FA1A S2_5_75 ( .A(\ab[5][75] ), .B(\CARRYB[4][75] ), .CI(\SUMB[4][76] ), 
        .CO(\CARRYB[5][75] ), .S(\SUMB[5][75] ) );
  FA1A S2_5_74 ( .A(\ab[5][74] ), .B(\CARRYB[4][74] ), .CI(\SUMB[4][75] ), 
        .CO(\CARRYB[5][74] ), .S(\SUMB[5][74] ) );
  FA1A S2_5_73 ( .A(\ab[5][73] ), .B(\CARRYB[4][73] ), .CI(\SUMB[4][74] ), 
        .CO(\CARRYB[5][73] ), .S(\SUMB[5][73] ) );
  FA1A S2_5_72 ( .A(\ab[5][72] ), .B(\CARRYB[4][72] ), .CI(\SUMB[4][73] ), 
        .CO(\CARRYB[5][72] ), .S(\SUMB[5][72] ) );
  FA1A S2_5_71 ( .A(\ab[5][71] ), .B(\CARRYB[4][71] ), .CI(\SUMB[4][72] ), 
        .CO(\CARRYB[5][71] ), .S(\SUMB[5][71] ) );
  FA1A S2_5_70 ( .A(\ab[5][70] ), .B(\CARRYB[4][70] ), .CI(\SUMB[4][71] ), 
        .CO(\CARRYB[5][70] ), .S(\SUMB[5][70] ) );
  FA1A S2_5_69 ( .A(\ab[5][69] ), .B(\CARRYB[4][69] ), .CI(\SUMB[4][70] ), 
        .CO(\CARRYB[5][69] ), .S(\SUMB[5][69] ) );
  FA1A S2_4_79 ( .A(\ab[4][79] ), .B(\CARRYB[3][79] ), .CI(\SUMB[3][80] ), 
        .CO(\CARRYB[4][79] ), .S(\SUMB[4][79] ) );
  FA1A S2_4_78 ( .A(\ab[4][78] ), .B(\CARRYB[3][78] ), .CI(\SUMB[3][79] ), 
        .CO(\CARRYB[4][78] ), .S(\SUMB[4][78] ) );
  FA1A S2_4_77 ( .A(\ab[4][77] ), .B(\CARRYB[3][77] ), .CI(\SUMB[3][78] ), 
        .CO(\CARRYB[4][77] ), .S(\SUMB[4][77] ) );
  FA1A S2_4_76 ( .A(\ab[4][76] ), .B(\CARRYB[3][76] ), .CI(\SUMB[3][77] ), 
        .CO(\CARRYB[4][76] ), .S(\SUMB[4][76] ) );
  FA1A S2_4_75 ( .A(\ab[4][75] ), .B(\CARRYB[3][75] ), .CI(\SUMB[3][76] ), 
        .CO(\CARRYB[4][75] ), .S(\SUMB[4][75] ) );
  FA1A S2_4_74 ( .A(\ab[4][74] ), .B(\CARRYB[3][74] ), .CI(\SUMB[3][75] ), 
        .CO(\CARRYB[4][74] ), .S(\SUMB[4][74] ) );
  FA1A S2_4_73 ( .A(\ab[4][73] ), .B(\CARRYB[3][73] ), .CI(\SUMB[3][74] ), 
        .CO(\CARRYB[4][73] ), .S(\SUMB[4][73] ) );
  FA1A S2_4_72 ( .A(\ab[4][72] ), .B(\CARRYB[3][72] ), .CI(\SUMB[3][73] ), 
        .CO(\CARRYB[4][72] ), .S(\SUMB[4][72] ) );
  FA1A S2_4_71 ( .A(\ab[4][71] ), .B(\CARRYB[3][71] ), .CI(\SUMB[3][72] ), 
        .CO(\CARRYB[4][71] ), .S(\SUMB[4][71] ) );
  FA1A S2_4_70 ( .A(\ab[4][70] ), .B(\CARRYB[3][70] ), .CI(\SUMB[3][71] ), 
        .CO(\CARRYB[4][70] ), .S(\SUMB[4][70] ) );
  FA1A S2_4_69 ( .A(\ab[4][69] ), .B(\CARRYB[3][69] ), .CI(\SUMB[3][70] ), 
        .CO(\CARRYB[4][69] ), .S(\SUMB[4][69] ) );
  FA1A S2_3_79 ( .A(\ab[3][79] ), .B(\CARRYB[2][79] ), .CI(\SUMB[2][80] ), 
        .CO(\CARRYB[3][79] ), .S(\SUMB[3][79] ) );
  FA1A S2_3_78 ( .A(\ab[3][78] ), .B(\CARRYB[2][78] ), .CI(\SUMB[2][79] ), 
        .CO(\CARRYB[3][78] ), .S(\SUMB[3][78] ) );
  FA1A S2_3_77 ( .A(\ab[3][77] ), .B(\CARRYB[2][77] ), .CI(\SUMB[2][78] ), 
        .CO(\CARRYB[3][77] ), .S(\SUMB[3][77] ) );
  FA1A S2_3_76 ( .A(\ab[3][76] ), .B(\CARRYB[2][76] ), .CI(\SUMB[2][77] ), 
        .CO(\CARRYB[3][76] ), .S(\SUMB[3][76] ) );
  FA1A S2_3_75 ( .A(\ab[3][75] ), .B(\CARRYB[2][75] ), .CI(\SUMB[2][76] ), 
        .CO(\CARRYB[3][75] ), .S(\SUMB[3][75] ) );
  FA1A S2_3_74 ( .A(\ab[3][74] ), .B(\CARRYB[2][74] ), .CI(\SUMB[2][75] ), 
        .CO(\CARRYB[3][74] ), .S(\SUMB[3][74] ) );
  FA1A S2_3_73 ( .A(\ab[3][73] ), .B(\CARRYB[2][73] ), .CI(\SUMB[2][74] ), 
        .CO(\CARRYB[3][73] ), .S(\SUMB[3][73] ) );
  FA1A S2_3_72 ( .A(\ab[3][72] ), .B(\CARRYB[2][72] ), .CI(\SUMB[2][73] ), 
        .CO(\CARRYB[3][72] ), .S(\SUMB[3][72] ) );
  FA1A S2_3_71 ( .A(\ab[3][71] ), .B(\CARRYB[2][71] ), .CI(\SUMB[2][72] ), 
        .CO(\CARRYB[3][71] ), .S(\SUMB[3][71] ) );
  FA1A S2_3_70 ( .A(\ab[3][70] ), .B(\CARRYB[2][70] ), .CI(\SUMB[2][71] ), 
        .CO(\CARRYB[3][70] ), .S(\SUMB[3][70] ) );
  FA1A S2_3_69 ( .A(\ab[3][69] ), .B(\CARRYB[2][69] ), .CI(\SUMB[2][70] ), 
        .CO(\CARRYB[3][69] ), .S(\SUMB[3][69] ) );
  FA1A S2_2_79 ( .A(\ab[2][79] ), .B(\CARRYB[1][79] ), .CI(\SUMB[1][80] ), 
        .CO(\CARRYB[2][79] ), .S(\SUMB[2][79] ) );
  FA1A S2_2_78 ( .A(\ab[2][78] ), .B(\CARRYB[1][78] ), .CI(\SUMB[1][79] ), 
        .CO(\CARRYB[2][78] ), .S(\SUMB[2][78] ) );
  FA1A S2_2_77 ( .A(\ab[2][77] ), .B(\CARRYB[1][77] ), .CI(\SUMB[1][78] ), 
        .CO(\CARRYB[2][77] ), .S(\SUMB[2][77] ) );
  FA1A S2_2_76 ( .A(\ab[2][76] ), .B(\CARRYB[1][76] ), .CI(\SUMB[1][77] ), 
        .CO(\CARRYB[2][76] ), .S(\SUMB[2][76] ) );
  FA1A S2_2_75 ( .A(\ab[2][75] ), .B(\CARRYB[1][75] ), .CI(\SUMB[1][76] ), 
        .CO(\CARRYB[2][75] ), .S(\SUMB[2][75] ) );
  FA1A S2_2_74 ( .A(\ab[2][74] ), .B(\CARRYB[1][74] ), .CI(\SUMB[1][75] ), 
        .CO(\CARRYB[2][74] ), .S(\SUMB[2][74] ) );
  FA1A S2_2_73 ( .A(\ab[2][73] ), .B(\CARRYB[1][73] ), .CI(\SUMB[1][74] ), 
        .CO(\CARRYB[2][73] ), .S(\SUMB[2][73] ) );
  FA1A S2_2_72 ( .A(\ab[2][72] ), .B(\CARRYB[1][72] ), .CI(\SUMB[1][73] ), 
        .CO(\CARRYB[2][72] ), .S(\SUMB[2][72] ) );
  FA1A S2_2_71 ( .A(\ab[2][71] ), .B(\CARRYB[1][71] ), .CI(\SUMB[1][72] ), 
        .CO(\CARRYB[2][71] ), .S(\SUMB[2][71] ) );
  FA1A S2_2_70 ( .A(\ab[2][70] ), .B(\CARRYB[1][70] ), .CI(\SUMB[1][71] ), 
        .CO(\CARRYB[2][70] ), .S(\SUMB[2][70] ) );
  FA1A S2_2_69 ( .A(\ab[2][69] ), .B(\CARRYB[1][69] ), .CI(\SUMB[1][70] ), 
        .CO(\CARRYB[2][69] ), .S(\SUMB[2][69] ) );
  FA1A S4_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), .CO(
        \CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA1A S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA1A S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA1A S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA1A S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA1A S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA1A S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA1A S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA1A S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1A S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1A S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA1A S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1A S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1A S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1A S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S4_30 ( .A(\ab[29][30] ), .B(\CARRYB[28][30] ), .CI(\SUMB[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FA1A S4_29 ( .A(\ab[29][29] ), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), 
        .CO(\CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_28_30 ( .A(\ab[28][30] ), .B(\CARRYB[27][30] ), .CI(\SUMB[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA1A S2_28_29 ( .A(\ab[28][29] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_27_30 ( .A(\ab[27][30] ), .B(\CARRYB[26][30] ), .CI(\SUMB[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_27_29 ( .A(\ab[27][29] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_26_29 ( .A(\ab[26][29] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA1A S2_26_30 ( .A(\ab[26][30] ), .B(\CARRYB[25][30] ), .CI(\SUMB[25][31] ), 
        .CO(\CARRYB[26][30] ), .S(\SUMB[26][30] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_25_30 ( .A(\ab[25][30] ), .B(\CARRYB[24][30] ), .CI(\SUMB[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_25_29 ( .A(\ab[25][29] ), .B(\CARRYB[24][29] ), .CI(\SUMB[24][30] ), 
        .CO(\CARRYB[25][29] ), .S(\SUMB[25][29] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_24_29 ( .A(\ab[24][29] ), .B(\CARRYB[23][29] ), .CI(\SUMB[23][30] ), 
        .CO(\CARRYB[24][29] ), .S(\SUMB[24][29] ) );
  FA1A S2_24_30 ( .A(\ab[24][30] ), .B(\CARRYB[23][30] ), .CI(\SUMB[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_23_30 ( .A(\ab[23][30] ), .B(\CARRYB[22][30] ), .CI(\SUMB[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_23_29 ( .A(\ab[23][29] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA1A S2_22_30 ( .A(\ab[22][30] ), .B(\CARRYB[21][30] ), .CI(\SUMB[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA1A S2_22_29 ( .A(\ab[22][29] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA1A S2_21_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\SUMB[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA1A S2_21_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA1A S2_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\SUMB[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA1A S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA1A S2_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\SUMB[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA1A S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA1A S2_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\SUMB[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA1A S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA1A S2_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\SUMB[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA1A S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA1A S2_14_68 ( .A(\ab[14][68] ), .B(\CARRYB[13][68] ), .CI(\SUMB[13][69] ), 
        .CO(\CARRYB[14][68] ), .S(\SUMB[14][68] ) );
  FA1A S2_14_67 ( .A(\ab[14][67] ), .B(\CARRYB[13][67] ), .CI(\SUMB[13][68] ), 
        .CO(\CARRYB[14][67] ), .S(\SUMB[14][67] ) );
  FA1A S2_14_66 ( .A(\ab[14][66] ), .B(\CARRYB[13][66] ), .CI(\SUMB[13][67] ), 
        .CO(\CARRYB[14][66] ), .S(\SUMB[14][66] ) );
  FA1A S2_14_65 ( .A(\ab[14][65] ), .B(\CARRYB[13][65] ), .CI(\SUMB[13][66] ), 
        .CO(\CARRYB[14][65] ), .S(\SUMB[14][65] ) );
  FA1A S2_14_64 ( .A(\ab[14][64] ), .B(\CARRYB[13][64] ), .CI(\SUMB[13][65] ), 
        .CO(\CARRYB[14][64] ), .S(\SUMB[14][64] ) );
  FA1A S2_14_60 ( .A(\ab[14][60] ), .B(\CARRYB[13][60] ), .CI(\SUMB[13][61] ), 
        .CO(\CARRYB[14][60] ), .S(\SUMB[14][60] ) );
  FA1A S2_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\SUMB[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA1A S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA1A S2_13_68 ( .A(\ab[13][68] ), .B(\CARRYB[12][68] ), .CI(\SUMB[12][69] ), 
        .CO(\CARRYB[13][68] ), .S(\SUMB[13][68] ) );
  FA1A S2_13_67 ( .A(\ab[13][67] ), .B(\CARRYB[12][67] ), .CI(\SUMB[12][68] ), 
        .CO(\CARRYB[13][67] ), .S(\SUMB[13][67] ) );
  FA1A S2_13_66 ( .A(\ab[13][66] ), .B(\CARRYB[12][66] ), .CI(\SUMB[12][67] ), 
        .CO(\CARRYB[13][66] ), .S(\SUMB[13][66] ) );
  FA1A S2_13_65 ( .A(\ab[13][65] ), .B(\CARRYB[12][65] ), .CI(\SUMB[12][66] ), 
        .CO(\CARRYB[13][65] ), .S(\SUMB[13][65] ) );
  FA1A S2_13_64 ( .A(\ab[13][64] ), .B(\CARRYB[12][64] ), .CI(\SUMB[12][65] ), 
        .CO(\CARRYB[13][64] ), .S(\SUMB[13][64] ) );
  FA1A S2_13_60 ( .A(\ab[13][60] ), .B(\CARRYB[12][60] ), .CI(\SUMB[12][61] ), 
        .CO(\CARRYB[13][60] ), .S(\SUMB[13][60] ) );
  FA1A S2_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\SUMB[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA1A S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA1A S2_12_68 ( .A(\ab[12][68] ), .B(\CARRYB[11][68] ), .CI(\SUMB[11][69] ), 
        .CO(\CARRYB[12][68] ), .S(\SUMB[12][68] ) );
  FA1A S2_12_67 ( .A(\ab[12][67] ), .B(\CARRYB[11][67] ), .CI(\SUMB[11][68] ), 
        .CO(\CARRYB[12][67] ), .S(\SUMB[12][67] ) );
  FA1A S2_12_66 ( .A(\ab[12][66] ), .B(\CARRYB[11][66] ), .CI(\SUMB[11][67] ), 
        .CO(\CARRYB[12][66] ), .S(\SUMB[12][66] ) );
  FA1A S2_12_65 ( .A(\ab[12][65] ), .B(\CARRYB[11][65] ), .CI(\SUMB[11][66] ), 
        .CO(\CARRYB[12][65] ), .S(\SUMB[12][65] ) );
  FA1A S2_12_64 ( .A(\ab[12][64] ), .B(\CARRYB[11][64] ), .CI(\SUMB[11][65] ), 
        .CO(\CARRYB[12][64] ), .S(\SUMB[12][64] ) );
  FA1A S2_12_60 ( .A(\ab[12][60] ), .B(\CARRYB[11][60] ), .CI(\SUMB[11][61] ), 
        .CO(\CARRYB[12][60] ), .S(\SUMB[12][60] ) );
  FA1A S2_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\SUMB[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA1A S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA1A S2_11_68 ( .A(\ab[11][68] ), .B(\CARRYB[10][68] ), .CI(\SUMB[10][69] ), 
        .CO(\CARRYB[11][68] ), .S(\SUMB[11][68] ) );
  FA1A S2_11_67 ( .A(\ab[11][67] ), .B(\CARRYB[10][67] ), .CI(\SUMB[10][68] ), 
        .CO(\CARRYB[11][67] ), .S(\SUMB[11][67] ) );
  FA1A S2_11_66 ( .A(\ab[11][66] ), .B(\CARRYB[10][66] ), .CI(\SUMB[10][67] ), 
        .CO(\CARRYB[11][66] ), .S(\SUMB[11][66] ) );
  FA1A S2_11_65 ( .A(\ab[11][65] ), .B(\CARRYB[10][65] ), .CI(\SUMB[10][66] ), 
        .CO(\CARRYB[11][65] ), .S(\SUMB[11][65] ) );
  FA1A S2_11_64 ( .A(\ab[11][64] ), .B(\CARRYB[10][64] ), .CI(\SUMB[10][65] ), 
        .CO(\CARRYB[11][64] ), .S(\SUMB[11][64] ) );
  FA1A S2_11_60 ( .A(\ab[11][60] ), .B(\CARRYB[10][60] ), .CI(\SUMB[10][61] ), 
        .CO(\CARRYB[11][60] ), .S(\SUMB[11][60] ) );
  FA1A S2_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\SUMB[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA1A S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA1A S2_10_68 ( .A(\ab[10][68] ), .B(\CARRYB[9][68] ), .CI(\SUMB[9][69] ), 
        .CO(\CARRYB[10][68] ), .S(\SUMB[10][68] ) );
  FA1A S2_10_67 ( .A(\ab[10][67] ), .B(\CARRYB[9][67] ), .CI(\SUMB[9][68] ), 
        .CO(\CARRYB[10][67] ), .S(\SUMB[10][67] ) );
  FA1A S2_10_66 ( .A(\ab[10][66] ), .B(\CARRYB[9][66] ), .CI(\SUMB[9][67] ), 
        .CO(\CARRYB[10][66] ), .S(\SUMB[10][66] ) );
  FA1A S2_10_65 ( .A(\ab[10][65] ), .B(\CARRYB[9][65] ), .CI(\SUMB[9][66] ), 
        .CO(\CARRYB[10][65] ), .S(\SUMB[10][65] ) );
  FA1A S2_10_64 ( .A(\ab[10][64] ), .B(\CARRYB[9][64] ), .CI(\SUMB[9][65] ), 
        .CO(\CARRYB[10][64] ), .S(\SUMB[10][64] ) );
  FA1A S2_10_60 ( .A(\ab[10][60] ), .B(\CARRYB[9][60] ), .CI(\SUMB[9][61] ), 
        .CO(\CARRYB[10][60] ), .S(\SUMB[10][60] ) );
  FA1A S2_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\SUMB[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA1A S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA1A S2_9_68 ( .A(\ab[9][68] ), .B(\CARRYB[8][68] ), .CI(\SUMB[8][69] ), 
        .CO(\CARRYB[9][68] ), .S(\SUMB[9][68] ) );
  FA1A S2_9_67 ( .A(\ab[9][67] ), .B(\CARRYB[8][67] ), .CI(\SUMB[8][68] ), 
        .CO(\CARRYB[9][67] ), .S(\SUMB[9][67] ) );
  FA1A S2_9_66 ( .A(\ab[9][66] ), .B(\CARRYB[8][66] ), .CI(\SUMB[8][67] ), 
        .CO(\CARRYB[9][66] ), .S(\SUMB[9][66] ) );
  FA1A S2_9_65 ( .A(\ab[9][65] ), .B(\CARRYB[8][65] ), .CI(\SUMB[8][66] ), 
        .CO(\CARRYB[9][65] ), .S(\SUMB[9][65] ) );
  FA1A S2_9_64 ( .A(\ab[9][64] ), .B(\CARRYB[8][64] ), .CI(\SUMB[8][65] ), 
        .CO(\CARRYB[9][64] ), .S(\SUMB[9][64] ) );
  FA1A S2_9_60 ( .A(\ab[9][60] ), .B(\CARRYB[8][60] ), .CI(\SUMB[8][61] ), 
        .CO(\CARRYB[9][60] ), .S(\SUMB[9][60] ) );
  FA1A S2_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\SUMB[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA1A S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1A S2_8_68 ( .A(\ab[8][68] ), .B(\CARRYB[7][68] ), .CI(\SUMB[7][69] ), 
        .CO(\CARRYB[8][68] ), .S(\SUMB[8][68] ) );
  FA1A S2_8_67 ( .A(\ab[8][67] ), .B(\CARRYB[7][67] ), .CI(\SUMB[7][68] ), 
        .CO(\CARRYB[8][67] ), .S(\SUMB[8][67] ) );
  FA1A S2_8_66 ( .A(\ab[8][66] ), .B(\CARRYB[7][66] ), .CI(\SUMB[7][67] ), 
        .CO(\CARRYB[8][66] ), .S(\SUMB[8][66] ) );
  FA1A S2_8_65 ( .A(\ab[8][65] ), .B(\CARRYB[7][65] ), .CI(\SUMB[7][66] ), 
        .CO(\CARRYB[8][65] ), .S(\SUMB[8][65] ) );
  FA1A S2_8_64 ( .A(\ab[8][64] ), .B(\CARRYB[7][64] ), .CI(\SUMB[7][65] ), 
        .CO(\CARRYB[8][64] ), .S(\SUMB[8][64] ) );
  FA1A S2_8_60 ( .A(\ab[8][60] ), .B(\CARRYB[7][60] ), .CI(\SUMB[7][61] ), 
        .CO(\CARRYB[8][60] ), .S(\SUMB[8][60] ) );
  FA1A S2_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\SUMB[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA1A S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1A S2_7_68 ( .A(\ab[7][68] ), .B(\CARRYB[6][68] ), .CI(\SUMB[6][69] ), 
        .CO(\CARRYB[7][68] ), .S(\SUMB[7][68] ) );
  FA1A S2_7_67 ( .A(\ab[7][67] ), .B(\CARRYB[6][67] ), .CI(\SUMB[6][68] ), 
        .CO(\CARRYB[7][67] ), .S(\SUMB[7][67] ) );
  FA1A S2_7_66 ( .A(\ab[7][66] ), .B(\CARRYB[6][66] ), .CI(\SUMB[6][67] ), 
        .CO(\CARRYB[7][66] ), .S(\SUMB[7][66] ) );
  FA1A S2_7_65 ( .A(\ab[7][65] ), .B(\CARRYB[6][65] ), .CI(\SUMB[6][66] ), 
        .CO(\CARRYB[7][65] ), .S(\SUMB[7][65] ) );
  FA1A S2_7_64 ( .A(\ab[7][64] ), .B(\CARRYB[6][64] ), .CI(\SUMB[6][65] ), 
        .CO(\CARRYB[7][64] ), .S(\SUMB[7][64] ) );
  FA1A S2_7_60 ( .A(\ab[7][60] ), .B(\CARRYB[6][60] ), .CI(\SUMB[6][61] ), 
        .CO(\CARRYB[7][60] ), .S(\SUMB[7][60] ) );
  FA1A S2_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\SUMB[8][31] ), 
        .CO(\CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA1A S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1A S2_6_68 ( .A(\ab[6][68] ), .B(\CARRYB[5][68] ), .CI(\SUMB[5][69] ), 
        .CO(\CARRYB[6][68] ), .S(\SUMB[6][68] ) );
  FA1A S2_6_67 ( .A(\ab[6][67] ), .B(\CARRYB[5][67] ), .CI(\SUMB[5][68] ), 
        .CO(\CARRYB[6][67] ), .S(\SUMB[6][67] ) );
  FA1A S2_6_66 ( .A(\ab[6][66] ), .B(\CARRYB[5][66] ), .CI(\SUMB[5][67] ), 
        .CO(\CARRYB[6][66] ), .S(\SUMB[6][66] ) );
  FA1A S2_6_65 ( .A(\ab[6][65] ), .B(\CARRYB[5][65] ), .CI(\SUMB[5][66] ), 
        .CO(\CARRYB[6][65] ), .S(\SUMB[6][65] ) );
  FA1A S2_6_64 ( .A(\ab[6][64] ), .B(\CARRYB[5][64] ), .CI(\SUMB[5][65] ), 
        .CO(\CARRYB[6][64] ), .S(\SUMB[6][64] ) );
  FA1A S2_6_60 ( .A(\ab[6][60] ), .B(\CARRYB[5][60] ), .CI(\SUMB[5][61] ), 
        .CO(\CARRYB[6][60] ), .S(\SUMB[6][60] ) );
  FA1A S2_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\SUMB[7][31] ), 
        .CO(\CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA1A S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1A S2_5_68 ( .A(\ab[5][68] ), .B(\CARRYB[4][68] ), .CI(\SUMB[4][69] ), 
        .CO(\CARRYB[5][68] ), .S(\SUMB[5][68] ) );
  FA1A S2_5_67 ( .A(\ab[5][67] ), .B(\CARRYB[4][67] ), .CI(\SUMB[4][68] ), 
        .CO(\CARRYB[5][67] ), .S(\SUMB[5][67] ) );
  FA1A S2_5_66 ( .A(\ab[5][66] ), .B(\CARRYB[4][66] ), .CI(\SUMB[4][67] ), 
        .CO(\CARRYB[5][66] ), .S(\SUMB[5][66] ) );
  FA1A S2_5_65 ( .A(\ab[5][65] ), .B(\CARRYB[4][65] ), .CI(\SUMB[4][66] ), 
        .CO(\CARRYB[5][65] ), .S(\SUMB[5][65] ) );
  FA1A S2_5_64 ( .A(\ab[5][64] ), .B(\CARRYB[4][64] ), .CI(\SUMB[4][65] ), 
        .CO(\CARRYB[5][64] ), .S(\SUMB[5][64] ) );
  FA1A S2_5_60 ( .A(\ab[5][60] ), .B(\CARRYB[4][60] ), .CI(\SUMB[4][61] ), 
        .CO(\CARRYB[5][60] ), .S(\SUMB[5][60] ) );
  FA1A S2_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\SUMB[6][31] ), 
        .CO(\CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA1A S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1A S2_4_68 ( .A(\ab[4][68] ), .B(\CARRYB[3][68] ), .CI(\SUMB[3][69] ), 
        .CO(\CARRYB[4][68] ), .S(\SUMB[4][68] ) );
  FA1A S2_4_67 ( .A(\ab[4][67] ), .B(\CARRYB[3][67] ), .CI(\SUMB[3][68] ), 
        .CO(\CARRYB[4][67] ), .S(\SUMB[4][67] ) );
  FA1A S2_4_66 ( .A(\ab[4][66] ), .B(\CARRYB[3][66] ), .CI(\SUMB[3][67] ), 
        .CO(\CARRYB[4][66] ), .S(\SUMB[4][66] ) );
  FA1A S2_4_65 ( .A(\ab[4][65] ), .B(\CARRYB[3][65] ), .CI(\SUMB[3][66] ), 
        .CO(\CARRYB[4][65] ), .S(\SUMB[4][65] ) );
  FA1A S2_4_64 ( .A(\ab[4][64] ), .B(\CARRYB[3][64] ), .CI(\SUMB[3][65] ), 
        .CO(\CARRYB[4][64] ), .S(\SUMB[4][64] ) );
  FA1A S2_4_60 ( .A(\ab[4][60] ), .B(\CARRYB[3][60] ), .CI(\SUMB[3][61] ), 
        .CO(\CARRYB[4][60] ), .S(\SUMB[4][60] ) );
  FA1A S2_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\SUMB[5][31] ), 
        .CO(\CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA1A S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA1A S2_3_68 ( .A(\ab[3][68] ), .B(\CARRYB[2][68] ), .CI(\SUMB[2][69] ), 
        .CO(\CARRYB[3][68] ), .S(\SUMB[3][68] ) );
  FA1A S2_3_67 ( .A(\ab[3][67] ), .B(\CARRYB[2][67] ), .CI(\SUMB[2][68] ), 
        .CO(\CARRYB[3][67] ), .S(\SUMB[3][67] ) );
  FA1A S2_3_66 ( .A(\ab[3][66] ), .B(\CARRYB[2][66] ), .CI(\SUMB[2][67] ), 
        .CO(\CARRYB[3][66] ), .S(\SUMB[3][66] ) );
  FA1A S2_3_65 ( .A(\ab[3][65] ), .B(\CARRYB[2][65] ), .CI(\SUMB[2][66] ), 
        .CO(\CARRYB[3][65] ), .S(\SUMB[3][65] ) );
  FA1A S2_3_64 ( .A(\ab[3][64] ), .B(\CARRYB[2][64] ), .CI(\SUMB[2][65] ), 
        .CO(\CARRYB[3][64] ), .S(\SUMB[3][64] ) );
  FA1A S2_3_60 ( .A(\ab[3][60] ), .B(\CARRYB[2][60] ), .CI(\SUMB[2][61] ), 
        .CO(\CARRYB[3][60] ), .S(\SUMB[3][60] ) );
  FA1A S2_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\SUMB[4][31] ), 
        .CO(\CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA1A S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA1A S2_2_68 ( .A(\ab[2][68] ), .B(\CARRYB[1][68] ), .CI(\SUMB[1][69] ), 
        .CO(\CARRYB[2][68] ), .S(\SUMB[2][68] ) );
  FA1A S2_2_67 ( .A(\ab[2][67] ), .B(\CARRYB[1][67] ), .CI(\SUMB[1][68] ), 
        .CO(\CARRYB[2][67] ), .S(\SUMB[2][67] ) );
  FA1A S2_2_66 ( .A(\ab[2][66] ), .B(\CARRYB[1][66] ), .CI(\SUMB[1][67] ), 
        .CO(\CARRYB[2][66] ), .S(\SUMB[2][66] ) );
  FA1A S2_2_65 ( .A(\ab[2][65] ), .B(\CARRYB[1][65] ), .CI(\SUMB[1][66] ), 
        .CO(\CARRYB[2][65] ), .S(\SUMB[2][65] ) );
  FA1A S2_2_64 ( .A(\ab[2][64] ), .B(\CARRYB[1][64] ), .CI(\SUMB[1][65] ), 
        .CO(\CARRYB[2][64] ), .S(\SUMB[2][64] ) );
  FA1A S2_2_60 ( .A(\ab[2][60] ), .B(\CARRYB[1][60] ), .CI(\SUMB[1][61] ), 
        .CO(\CARRYB[2][60] ), .S(\SUMB[2][60] ) );
  FA1A S2_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\SUMB[3][31] ), 
        .CO(\CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA1A S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\SUMB[3][30] ), 
        .CO(\CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1A S2_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .CI(\SUMB[2][31] ), 
        .CO(\CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA1A S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1A S2_2_30 ( .A(\ab[2][30] ), .B(\CARRYB[1][30] ), .CI(\SUMB[1][31] ), 
        .CO(\CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  FA1A S2_2_29 ( .A(\ab[2][29] ), .B(\CARRYB[1][29] ), .CI(\SUMB[1][30] ), 
        .CO(\CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1A S4_33 ( .A(\ab[29][33] ), .B(\CARRYB[28][33] ), .CI(\SUMB[28][34] ), 
        .CO(\CARRYB[29][33] ), .S(\SUMB[29][33] ) );
  FA1A S4_34 ( .A(\ab[29][34] ), .B(\CARRYB[28][34] ), .CI(\SUMB[28][35] ), 
        .CO(\CARRYB[29][34] ), .S(\SUMB[29][34] ) );
  FA1A S4_31 ( .A(\ab[29][31] ), .B(\CARRYB[28][31] ), .CI(\SUMB[28][32] ), 
        .CO(\CARRYB[29][31] ), .S(\SUMB[29][31] ) );
  FA1A S2_28_33 ( .A(\ab[28][33] ), .B(\CARRYB[27][33] ), .CI(\SUMB[27][34] ), 
        .CO(\CARRYB[28][33] ), .S(\SUMB[28][33] ) );
  FA1A S2_28_32 ( .A(\ab[28][32] ), .B(\CARRYB[27][32] ), .CI(\SUMB[27][33] ), 
        .CO(\CARRYB[28][32] ), .S(\SUMB[28][32] ) );
  FA1A S2_28_34 ( .A(\ab[28][34] ), .B(\CARRYB[27][34] ), .CI(\SUMB[27][35] ), 
        .CO(\CARRYB[28][34] ), .S(\SUMB[28][34] ) );
  FA1A S4_37 ( .A(\ab[29][37] ), .B(\CARRYB[28][37] ), .CI(\SUMB[28][38] ), 
        .CO(\CARRYB[29][37] ), .S(\SUMB[29][37] ) );
  FA1A S2_27_34 ( .A(\ab[27][34] ), .B(\CARRYB[26][34] ), .CI(\SUMB[26][35] ), 
        .CO(\CARRYB[27][34] ), .S(\SUMB[27][34] ) );
  FA1A S2_27_33 ( .A(\ab[27][33] ), .B(\CARRYB[26][33] ), .CI(\SUMB[26][34] ), 
        .CO(\CARRYB[27][33] ), .S(\SUMB[27][33] ) );
  FA1A S2_28_37 ( .A(\ab[28][37] ), .B(\CARRYB[27][37] ), .CI(\SUMB[27][38] ), 
        .CO(\CARRYB[28][37] ), .S(\SUMB[28][37] ) );
  FA1A S2_28_36 ( .A(\ab[28][36] ), .B(\CARRYB[27][36] ), .CI(\SUMB[27][37] ), 
        .CO(\CARRYB[28][36] ), .S(\SUMB[28][36] ) );
  FA1A S2_28_35 ( .A(\ab[28][35] ), .B(\CARRYB[27][35] ), .CI(\SUMB[27][36] ), 
        .CO(\CARRYB[28][35] ), .S(\SUMB[28][35] ) );
  FA1A S2_26_34 ( .A(\ab[26][34] ), .B(\CARRYB[25][34] ), .CI(\SUMB[25][35] ), 
        .CO(\CARRYB[26][34] ), .S(\SUMB[26][34] ) );
  FA1A S2_28_31 ( .A(\ab[28][31] ), .B(\CARRYB[27][31] ), .CI(\SUMB[27][32] ), 
        .CO(\CARRYB[28][31] ), .S(\SUMB[28][31] ) );
  FA1A S4_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), .CO(
        \CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA1A S2_27_37 ( .A(\ab[27][37] ), .B(\CARRYB[26][37] ), .CI(\SUMB[26][38] ), 
        .CO(\CARRYB[27][37] ), .S(\SUMB[27][37] ) );
  FA1A S2_27_36 ( .A(\ab[27][36] ), .B(\CARRYB[26][36] ), .CI(\SUMB[26][37] ), 
        .CO(\CARRYB[27][36] ), .S(\SUMB[27][36] ) );
  FA1A S2_27_35 ( .A(\ab[27][35] ), .B(\CARRYB[26][35] ), .CI(\SUMB[26][36] ), 
        .CO(\CARRYB[27][35] ), .S(\SUMB[27][35] ) );
  FA1A S2_27_32 ( .A(\ab[27][32] ), .B(\CARRYB[26][32] ), .CI(\SUMB[26][33] ), 
        .CO(\CARRYB[27][32] ), .S(\SUMB[27][32] ) );
  FA1A S2_27_31 ( .A(\ab[27][31] ), .B(\CARRYB[26][31] ), .CI(\SUMB[26][32] ), 
        .CO(\CARRYB[27][31] ), .S(\SUMB[27][31] ) );
  FA1A S4_27 ( .A(\ab[29][27] ), .B(\CARRYB[28][27] ), .CI(\SUMB[28][28] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA1A S4_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), .CO(
        \CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA1A S4_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), .CO(
        \CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA1A S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA1A S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA1A S2_26_37 ( .A(\ab[26][37] ), .B(\CARRYB[25][37] ), .CI(\SUMB[25][38] ), 
        .CO(\CARRYB[26][37] ), .S(\SUMB[26][37] ) );
  FA1A S2_26_36 ( .A(\ab[26][36] ), .B(\CARRYB[25][36] ), .CI(\SUMB[25][37] ), 
        .CO(\CARRYB[26][36] ), .S(\SUMB[26][36] ) );
  FA1A S2_28_38 ( .A(\ab[28][38] ), .B(\CARRYB[27][38] ), .CI(\SUMB[27][39] ), 
        .CO(\CARRYB[28][38] ), .S(\SUMB[28][38] ) );
  FA1A S2_26_35 ( .A(\ab[26][35] ), .B(\CARRYB[25][35] ), .CI(\SUMB[25][36] ), 
        .CO(\CARRYB[26][35] ), .S(\SUMB[26][35] ) );
  FA1A S2_26_33 ( .A(\ab[26][33] ), .B(\CARRYB[25][33] ), .CI(\SUMB[25][34] ), 
        .CO(\CARRYB[26][33] ), .S(\SUMB[26][33] ) );
  FA1A S2_26_32 ( .A(\ab[26][32] ), .B(\CARRYB[25][32] ), .CI(\SUMB[25][33] ), 
        .CO(\CARRYB[26][32] ), .S(\SUMB[26][32] ) );
  FA1A S2_26_31 ( .A(\ab[26][31] ), .B(\CARRYB[25][31] ), .CI(\SUMB[25][32] ), 
        .CO(\CARRYB[26][31] ), .S(\SUMB[26][31] ) );
  FA1A S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA1A S2_28_28 ( .A(\ab[28][28] ), .B(\CARRYB[27][28] ), .CI(\SUMB[27][29] ), 
        .CO(\CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA1A S4_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA1A S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA1A S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA1A S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA1A S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA1A S2_25_37 ( .A(\ab[25][37] ), .B(\CARRYB[24][37] ), .CI(\SUMB[24][38] ), 
        .CO(\CARRYB[25][37] ), .S(\SUMB[25][37] ) );
  FA1A S2_25_36 ( .A(\ab[25][36] ), .B(\CARRYB[24][36] ), .CI(\SUMB[24][37] ), 
        .CO(\CARRYB[25][36] ), .S(\SUMB[25][36] ) );
  FA1A S2_27_38 ( .A(\ab[27][38] ), .B(\CARRYB[26][38] ), .CI(\SUMB[26][39] ), 
        .CO(\CARRYB[27][38] ), .S(\SUMB[27][38] ) );
  FA1A S2_25_35 ( .A(\ab[25][35] ), .B(\CARRYB[24][35] ), .CI(\SUMB[24][36] ), 
        .CO(\CARRYB[25][35] ), .S(\SUMB[25][35] ) );
  FA1A S2_25_34 ( .A(\ab[25][34] ), .B(\CARRYB[24][34] ), .CI(\SUMB[24][35] ), 
        .CO(\CARRYB[25][34] ), .S(\SUMB[25][34] ) );
  FA1A S2_25_33 ( .A(\ab[25][33] ), .B(\CARRYB[24][33] ), .CI(\SUMB[24][34] ), 
        .CO(\CARRYB[25][33] ), .S(\SUMB[25][33] ) );
  FA1A S2_25_32 ( .A(\ab[25][32] ), .B(\CARRYB[24][32] ), .CI(\SUMB[24][33] ), 
        .CO(\CARRYB[25][32] ), .S(\SUMB[25][32] ) );
  FA1A S2_27_28 ( .A(\ab[27][28] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), 
        .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FA1A S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA1A S2_28_26 ( .A(\ab[28][26] ), .B(\CARRYB[27][26] ), .CI(\SUMB[27][27] ), 
        .CO(\CARRYB[28][26] ), .S(\SUMB[28][26] ) );
  FA1A S4_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA1A S4_22 ( .A(\ab[29][22] ), .B(\CARRYB[28][22] ), .CI(\SUMB[28][23] ), 
        .CO(\CARRYB[29][22] ), .S(\SUMB[29][22] ) );
  FA1A S4_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA1A S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA1A S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA1A S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA1A S2_28_7 ( .A(\ab[28][7] ), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA1A S2_28_6 ( .A(\ab[28][6] ), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA1A S2_24_37 ( .A(\ab[24][37] ), .B(\CARRYB[23][37] ), .CI(\SUMB[23][38] ), 
        .CO(\CARRYB[24][37] ), .S(\SUMB[24][37] ) );
  FA1A S2_24_36 ( .A(\ab[24][36] ), .B(\CARRYB[23][36] ), .CI(\SUMB[23][37] ), 
        .CO(\CARRYB[24][36] ), .S(\SUMB[24][36] ) );
  FA1A S2_26_38 ( .A(\ab[26][38] ), .B(\CARRYB[25][38] ), .CI(\SUMB[25][39] ), 
        .CO(\CARRYB[26][38] ), .S(\SUMB[26][38] ) );
  FA1A S2_24_35 ( .A(\ab[24][35] ), .B(\CARRYB[23][35] ), .CI(\SUMB[23][36] ), 
        .CO(\CARRYB[24][35] ), .S(\SUMB[24][35] ) );
  FA1A S2_24_34 ( .A(\ab[24][34] ), .B(\CARRYB[23][34] ), .CI(\SUMB[23][35] ), 
        .CO(\CARRYB[24][34] ), .S(\SUMB[24][34] ) );
  FA1A S2_24_33 ( .A(\ab[24][33] ), .B(\CARRYB[23][33] ), .CI(\SUMB[23][34] ), 
        .CO(\CARRYB[24][33] ), .S(\SUMB[24][33] ) );
  FA1A S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA1A S2_27_27 ( .A(\ab[27][27] ), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), 
        .CO(\CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA1A S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA1A S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA1A S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA1A S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA1A S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA1A S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA1A S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA1A S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA1A S2_27_7 ( .A(\ab[27][7] ), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA1A S2_27_6 ( .A(\ab[27][6] ), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA1A S2_23_37 ( .A(\ab[23][37] ), .B(\CARRYB[22][37] ), .CI(\SUMB[22][38] ), 
        .CO(\CARRYB[23][37] ), .S(\SUMB[23][37] ) );
  FA1A S2_23_36 ( .A(\ab[23][36] ), .B(\CARRYB[22][36] ), .CI(\SUMB[22][37] ), 
        .CO(\CARRYB[23][36] ), .S(\SUMB[23][36] ) );
  FA1A S2_25_38 ( .A(\ab[25][38] ), .B(\CARRYB[24][38] ), .CI(\SUMB[24][39] ), 
        .CO(\CARRYB[25][38] ), .S(\SUMB[25][38] ) );
  FA1A S2_23_35 ( .A(\ab[23][35] ), .B(\CARRYB[22][35] ), .CI(\SUMB[22][36] ), 
        .CO(\CARRYB[23][35] ), .S(\SUMB[23][35] ) );
  FA1A S2_23_34 ( .A(\ab[23][34] ), .B(\CARRYB[22][34] ), .CI(\SUMB[22][35] ), 
        .CO(\CARRYB[23][34] ), .S(\SUMB[23][34] ) );
  FA1A S2_25_31 ( .A(\ab[25][31] ), .B(\CARRYB[24][31] ), .CI(\SUMB[24][32] ), 
        .CO(\CARRYB[25][31] ), .S(\SUMB[25][31] ) );
  FA1A S2_26_27 ( .A(\ab[26][27] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), 
        .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FA1A S2_26_28 ( .A(\ab[26][28] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), 
        .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FA1A S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA1A S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA1A S2_27_23 ( .A(\ab[27][23] ), .B(\CARRYB[26][23] ), .CI(\SUMB[26][24] ), 
        .CO(\CARRYB[27][23] ), .S(\SUMB[27][23] ) );
  FA1A S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), 
        .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FA1A S2_27_21 ( .A(\ab[27][21] ), .B(\CARRYB[26][21] ), .CI(\SUMB[26][22] ), 
        .CO(\CARRYB[27][21] ), .S(\SUMB[27][21] ) );
  FA1A S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA1A S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA1A S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA1A S2_26_8 ( .A(\ab[26][8] ), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA1A S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA1A S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA1A S2_22_37 ( .A(\ab[22][37] ), .B(\CARRYB[21][37] ), .CI(\SUMB[21][38] ), 
        .CO(\CARRYB[22][37] ), .S(\SUMB[22][37] ) );
  FA1A S2_22_36 ( .A(\ab[22][36] ), .B(\CARRYB[21][36] ), .CI(\SUMB[21][37] ), 
        .CO(\CARRYB[22][36] ), .S(\SUMB[22][36] ) );
  FA1A S2_24_38 ( .A(\ab[24][38] ), .B(\CARRYB[23][38] ), .CI(\SUMB[23][39] ), 
        .CO(\CARRYB[24][38] ), .S(\SUMB[24][38] ) );
  FA1A S2_22_35 ( .A(\ab[22][35] ), .B(\CARRYB[21][35] ), .CI(\SUMB[21][36] ), 
        .CO(\CARRYB[22][35] ), .S(\SUMB[22][35] ) );
  FA1A S2_24_31 ( .A(\ab[24][31] ), .B(\CARRYB[23][31] ), .CI(\SUMB[23][32] ), 
        .CO(\CARRYB[24][31] ), .S(\SUMB[24][31] ) );
  FA1A S2_24_32 ( .A(\ab[24][32] ), .B(\CARRYB[23][32] ), .CI(\SUMB[23][33] ), 
        .CO(\CARRYB[24][32] ), .S(\SUMB[24][32] ) );
  FA1A S2_25_28 ( .A(\ab[25][28] ), .B(\CARRYB[24][28] ), .CI(\SUMB[24][29] ), 
        .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FA1A S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), 
        .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA1A S2_26_25 ( .A(\ab[26][25] ), .B(\CARRYB[25][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA1A S2_26_24 ( .A(\ab[26][24] ), .B(\CARRYB[25][24] ), .CI(\SUMB[25][25] ), 
        .CO(\CARRYB[26][24] ), .S(\SUMB[26][24] ) );
  FA1A S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA1A S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA1A S2_26_21 ( .A(\ab[26][21] ), .B(\CARRYB[25][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA1A S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA1A S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA1A S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA1A S2_25_8 ( .A(\ab[25][8] ), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA1A S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA1A S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA1A S2_21_37 ( .A(\ab[21][37] ), .B(\CARRYB[20][37] ), .CI(\SUMB[20][38] ), 
        .CO(\CARRYB[21][37] ), .S(\SUMB[21][37] ) );
  FA1A S2_21_36 ( .A(\ab[21][36] ), .B(\CARRYB[20][36] ), .CI(\SUMB[20][37] ), 
        .CO(\CARRYB[21][36] ), .S(\SUMB[21][36] ) );
  FA1A S2_23_38 ( .A(\ab[23][38] ), .B(\CARRYB[22][38] ), .CI(\SUMB[22][39] ), 
        .CO(\CARRYB[23][38] ), .S(\SUMB[23][38] ) );
  FA1A S2_23_32 ( .A(\ab[23][32] ), .B(\CARRYB[22][32] ), .CI(\SUMB[22][33] ), 
        .CO(\CARRYB[23][32] ), .S(\SUMB[23][32] ) );
  FA1A S2_23_33 ( .A(\ab[23][33] ), .B(\CARRYB[22][33] ), .CI(\SUMB[22][34] ), 
        .CO(\CARRYB[23][33] ), .S(\SUMB[23][33] ) );
  FA1A S2_25_27 ( .A(\ab[25][27] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA1A S2_25_26 ( .A(\ab[25][26] ), .B(\CARRYB[24][26] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA1A S2_25_25 ( .A(\ab[25][25] ), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), 
        .CO(\CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA1A S2_25_24 ( .A(\ab[25][24] ), .B(\CARRYB[24][24] ), .CI(\SUMB[24][25] ), 
        .CO(\CARRYB[25][24] ), .S(\SUMB[25][24] ) );
  FA1A S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA1A S2_25_22 ( .A(\ab[25][22] ), .B(\CARRYB[24][22] ), .CI(\SUMB[24][23] ), 
        .CO(\CARRYB[25][22] ), .S(\SUMB[25][22] ) );
  FA1A S2_25_21 ( .A(\ab[25][21] ), .B(\CARRYB[24][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA1A S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA1A S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA1A S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA1A S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA1A S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA1A S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA1A S2_20_37 ( .A(\ab[20][37] ), .B(\CARRYB[19][37] ), .CI(\SUMB[19][38] ), 
        .CO(\CARRYB[20][37] ), .S(\SUMB[20][37] ) );
  FA1A S2_22_38 ( .A(\ab[22][38] ), .B(\CARRYB[21][38] ), .CI(\SUMB[21][39] ), 
        .CO(\CARRYB[22][38] ), .S(\SUMB[22][38] ) );
  FA1A S2_22_33 ( .A(\ab[22][33] ), .B(\CARRYB[21][33] ), .CI(\SUMB[21][34] ), 
        .CO(\CARRYB[22][33] ), .S(\SUMB[22][33] ) );
  FA1A S2_22_34 ( .A(\ab[22][34] ), .B(\CARRYB[21][34] ), .CI(\SUMB[21][35] ), 
        .CO(\CARRYB[22][34] ), .S(\SUMB[22][34] ) );
  FA1A S2_23_31 ( .A(\ab[23][31] ), .B(\CARRYB[22][31] ), .CI(\SUMB[22][32] ), 
        .CO(\CARRYB[23][31] ), .S(\SUMB[23][31] ) );
  FA1A S2_24_28 ( .A(\ab[24][28] ), .B(\CARRYB[23][28] ), .CI(\SUMB[23][29] ), 
        .CO(\CARRYB[24][28] ), .S(\SUMB[24][28] ) );
  FA1A S2_24_27 ( .A(\ab[24][27] ), .B(\CARRYB[23][27] ), .CI(\SUMB[23][28] ), 
        .CO(\CARRYB[24][27] ), .S(\SUMB[24][27] ) );
  FA1A S2_24_26 ( .A(\ab[24][26] ), .B(\CARRYB[23][26] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA1A S2_24_25 ( .A(\ab[24][25] ), .B(\CARRYB[23][25] ), .CI(\SUMB[23][26] ), 
        .CO(\CARRYB[24][25] ), .S(\SUMB[24][25] ) );
  FA1A S2_24_24 ( .A(\ab[24][24] ), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), 
        .CO(\CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA1A S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA1A S2_24_22 ( .A(\ab[24][22] ), .B(\CARRYB[23][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA1A S2_24_21 ( .A(\ab[24][21] ), .B(\CARRYB[23][21] ), .CI(\SUMB[23][22] ), 
        .CO(\CARRYB[24][21] ), .S(\SUMB[24][21] ) );
  FA1A S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA1A S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1A S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1A S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA1A S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA1A S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA1A S2_21_38 ( .A(\ab[21][38] ), .B(\CARRYB[20][38] ), .CI(\SUMB[20][39] ), 
        .CO(\CARRYB[21][38] ), .S(\SUMB[21][38] ) );
  FA1A S2_21_34 ( .A(\ab[21][34] ), .B(\CARRYB[20][34] ), .CI(\SUMB[20][35] ), 
        .CO(\CARRYB[21][34] ), .S(\SUMB[21][34] ) );
  FA1A S2_21_35 ( .A(\ab[21][35] ), .B(\CARRYB[20][35] ), .CI(\SUMB[20][36] ), 
        .CO(\CARRYB[21][35] ), .S(\SUMB[21][35] ) );
  FA1A S2_22_31 ( .A(\ab[22][31] ), .B(\CARRYB[21][31] ), .CI(\SUMB[21][32] ), 
        .CO(\CARRYB[22][31] ), .S(\SUMB[22][31] ) );
  FA1A S2_22_32 ( .A(\ab[22][32] ), .B(\CARRYB[21][32] ), .CI(\SUMB[21][33] ), 
        .CO(\CARRYB[22][32] ), .S(\SUMB[22][32] ) );
  FA1A S2_23_28 ( .A(\ab[23][28] ), .B(\CARRYB[22][28] ), .CI(\SUMB[22][29] ), 
        .CO(\CARRYB[23][28] ), .S(\SUMB[23][28] ) );
  FA1A S2_23_27 ( .A(\ab[23][27] ), .B(\CARRYB[22][27] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA1A S2_23_26 ( .A(\ab[23][26] ), .B(\CARRYB[22][26] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA1A S2_23_25 ( .A(\ab[23][25] ), .B(\CARRYB[22][25] ), .CI(\SUMB[22][26] ), 
        .CO(\CARRYB[23][25] ), .S(\SUMB[23][25] ) );
  FA1A S2_23_24 ( .A(\ab[23][24] ), .B(\CARRYB[22][24] ), .CI(\SUMB[22][25] ), 
        .CO(\CARRYB[23][24] ), .S(\SUMB[23][24] ) );
  FA1A S2_23_23 ( .A(\ab[23][23] ), .B(\CARRYB[22][23] ), .CI(\SUMB[22][24] ), 
        .CO(\CARRYB[23][23] ), .S(\SUMB[23][23] ) );
  FA1A S2_23_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA1A S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA1A S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1A S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1A S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA1A S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA1A S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA1A S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA1A S2_20_38 ( .A(\ab[20][38] ), .B(\CARRYB[19][38] ), .CI(\SUMB[19][39] ), 
        .CO(\CARRYB[20][38] ), .S(\SUMB[20][38] ) );
  FA1A S2_20_35 ( .A(\ab[20][35] ), .B(\CARRYB[19][35] ), .CI(\SUMB[19][36] ), 
        .CO(\CARRYB[20][35] ), .S(\SUMB[20][35] ) );
  FA1A S2_20_36 ( .A(\ab[20][36] ), .B(\CARRYB[19][36] ), .CI(\SUMB[19][37] ), 
        .CO(\CARRYB[20][36] ), .S(\SUMB[20][36] ) );
  FA1A S2_21_32 ( .A(\ab[21][32] ), .B(\CARRYB[20][32] ), .CI(\SUMB[20][33] ), 
        .CO(\CARRYB[21][32] ), .S(\SUMB[21][32] ) );
  FA1A S2_21_33 ( .A(\ab[21][33] ), .B(\CARRYB[20][33] ), .CI(\SUMB[20][34] ), 
        .CO(\CARRYB[21][33] ), .S(\SUMB[21][33] ) );
  FA1A S2_22_28 ( .A(\ab[22][28] ), .B(\CARRYB[21][28] ), .CI(\SUMB[21][29] ), 
        .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FA1A S2_22_27 ( .A(\ab[22][27] ), .B(\CARRYB[21][27] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA1A S2_22_26 ( .A(\ab[22][26] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA1A S2_22_25 ( .A(\ab[22][25] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA1A S2_22_24 ( .A(\ab[22][24] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA1A S2_22_23 ( .A(\ab[22][23] ), .B(\CARRYB[21][23] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA1A S2_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA1A S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA1A S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA1A S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1A S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1A S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1A S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA1A S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA1A S2_19_38 ( .A(\ab[19][38] ), .B(\CARRYB[18][38] ), .CI(\SUMB[18][39] ), 
        .CO(\CARRYB[19][38] ), .S(\SUMB[19][38] ) );
  FA1A S2_19_36 ( .A(\ab[19][36] ), .B(\CARRYB[18][36] ), .CI(\SUMB[18][37] ), 
        .CO(\CARRYB[19][36] ), .S(\SUMB[19][36] ) );
  FA1A S2_19_37 ( .A(\ab[19][37] ), .B(\CARRYB[18][37] ), .CI(\SUMB[18][38] ), 
        .CO(\CARRYB[19][37] ), .S(\SUMB[19][37] ) );
  FA1A S2_20_33 ( .A(\ab[20][33] ), .B(\CARRYB[19][33] ), .CI(\SUMB[19][34] ), 
        .CO(\CARRYB[20][33] ), .S(\SUMB[20][33] ) );
  FA1A S2_20_34 ( .A(\ab[20][34] ), .B(\CARRYB[19][34] ), .CI(\SUMB[19][35] ), 
        .CO(\CARRYB[20][34] ), .S(\SUMB[20][34] ) );
  FA1A S2_21_31 ( .A(\ab[21][31] ), .B(\CARRYB[20][31] ), .CI(\SUMB[20][32] ), 
        .CO(\CARRYB[21][31] ), .S(\SUMB[21][31] ) );
  FA1A S2_21_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA1A S2_21_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA1A S2_21_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA1A S2_21_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA1A S2_21_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA1A S2_21_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA1A S2_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA1A S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA1A S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1A S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1A S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1A S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA1A S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1A S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1A S2_18_38 ( .A(\ab[18][38] ), .B(\CARRYB[17][38] ), .CI(\SUMB[17][39] ), 
        .CO(\CARRYB[18][38] ), .S(\SUMB[18][38] ) );
  FA1A S2_18_37 ( .A(\ab[18][37] ), .B(\CARRYB[17][37] ), .CI(\SUMB[17][38] ), 
        .CO(\CARRYB[18][37] ), .S(\SUMB[18][37] ) );
  FA1A S2_19_34 ( .A(\ab[19][34] ), .B(\CARRYB[18][34] ), .CI(\SUMB[18][35] ), 
        .CO(\CARRYB[19][34] ), .S(\SUMB[19][34] ) );
  FA1A S2_19_35 ( .A(\ab[19][35] ), .B(\CARRYB[18][35] ), .CI(\SUMB[18][36] ), 
        .CO(\CARRYB[19][35] ), .S(\SUMB[19][35] ) );
  FA1A S2_20_32 ( .A(\ab[20][32] ), .B(\CARRYB[19][32] ), .CI(\SUMB[19][33] ), 
        .CO(\CARRYB[20][32] ), .S(\SUMB[20][32] ) );
  FA1A S2_20_31 ( .A(\ab[20][31] ), .B(\CARRYB[19][31] ), .CI(\SUMB[19][32] ), 
        .CO(\CARRYB[20][31] ), .S(\SUMB[20][31] ) );
  FA1A S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA1A S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA1A S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA1A S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA1A S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA1A S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA1A S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA1A S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA1A S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA1A S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1A S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1A S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1A S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA1A S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1A S2_17_38 ( .A(\ab[17][38] ), .B(\CARRYB[16][38] ), .CI(\SUMB[16][39] ), 
        .CO(\CARRYB[17][38] ), .S(\SUMB[17][38] ) );
  FA1A S2_18_35 ( .A(\ab[18][35] ), .B(\CARRYB[17][35] ), .CI(\SUMB[17][36] ), 
        .CO(\CARRYB[18][35] ), .S(\SUMB[18][35] ) );
  FA1A S2_18_36 ( .A(\ab[18][36] ), .B(\CARRYB[17][36] ), .CI(\SUMB[17][37] ), 
        .CO(\CARRYB[18][36] ), .S(\SUMB[18][36] ) );
  FA1A S2_19_33 ( .A(\ab[19][33] ), .B(\CARRYB[18][33] ), .CI(\SUMB[18][34] ), 
        .CO(\CARRYB[19][33] ), .S(\SUMB[19][33] ) );
  FA1A S2_19_32 ( .A(\ab[19][32] ), .B(\CARRYB[18][32] ), .CI(\SUMB[18][33] ), 
        .CO(\CARRYB[19][32] ), .S(\SUMB[19][32] ) );
  FA1A S2_19_31 ( .A(\ab[19][31] ), .B(\CARRYB[18][31] ), .CI(\SUMB[18][32] ), 
        .CO(\CARRYB[19][31] ), .S(\SUMB[19][31] ) );
  FA1A S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA1A S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA1A S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA1A S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA1A S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA1A S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA1A S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA1A S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA1A S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1A S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1A S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1A S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA1A S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1A S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA1A S2_17_36 ( .A(\ab[17][36] ), .B(\CARRYB[16][36] ), .CI(\SUMB[16][37] ), 
        .CO(\CARRYB[17][36] ), .S(\SUMB[17][36] ) );
  FA1A S2_17_37 ( .A(\ab[17][37] ), .B(\CARRYB[16][37] ), .CI(\SUMB[16][38] ), 
        .CO(\CARRYB[17][37] ), .S(\SUMB[17][37] ) );
  FA1A S2_18_34 ( .A(\ab[18][34] ), .B(\CARRYB[17][34] ), .CI(\SUMB[17][35] ), 
        .CO(\CARRYB[18][34] ), .S(\SUMB[18][34] ) );
  FA1A S2_18_33 ( .A(\ab[18][33] ), .B(\CARRYB[17][33] ), .CI(\SUMB[17][34] ), 
        .CO(\CARRYB[18][33] ), .S(\SUMB[18][33] ) );
  FA1A S2_18_32 ( .A(\ab[18][32] ), .B(\CARRYB[17][32] ), .CI(\SUMB[17][33] ), 
        .CO(\CARRYB[18][32] ), .S(\SUMB[18][32] ) );
  FA1A S2_18_31 ( .A(\ab[18][31] ), .B(\CARRYB[17][31] ), .CI(\SUMB[17][32] ), 
        .CO(\CARRYB[18][31] ), .S(\SUMB[18][31] ) );
  FA1A S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA1A S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA1A S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA1A S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA1A S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA1A S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA1A S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA1A S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA1A S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1A S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1A S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1A S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1A S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1A S2_16_37 ( .A(\ab[16][37] ), .B(\CARRYB[15][37] ), .CI(\SUMB[15][38] ), 
        .CO(\CARRYB[16][37] ), .S(\SUMB[16][37] ) );
  FA1A S2_16_38 ( .A(\ab[16][38] ), .B(\CARRYB[15][38] ), .CI(\SUMB[15][39] ), 
        .CO(\CARRYB[16][38] ), .S(\SUMB[16][38] ) );
  FA1A S2_17_35 ( .A(\ab[17][35] ), .B(\CARRYB[16][35] ), .CI(\SUMB[16][36] ), 
        .CO(\CARRYB[17][35] ), .S(\SUMB[17][35] ) );
  FA1A S2_17_34 ( .A(\ab[17][34] ), .B(\CARRYB[16][34] ), .CI(\SUMB[16][35] ), 
        .CO(\CARRYB[17][34] ), .S(\SUMB[17][34] ) );
  FA1A S2_17_33 ( .A(\ab[17][33] ), .B(\CARRYB[16][33] ), .CI(\SUMB[16][34] ), 
        .CO(\CARRYB[17][33] ), .S(\SUMB[17][33] ) );
  FA1A S2_17_32 ( .A(\ab[17][32] ), .B(\CARRYB[16][32] ), .CI(\SUMB[16][33] ), 
        .CO(\CARRYB[17][32] ), .S(\SUMB[17][32] ) );
  FA1A S2_17_31 ( .A(\ab[17][31] ), .B(\CARRYB[16][31] ), .CI(\SUMB[16][32] ), 
        .CO(\CARRYB[17][31] ), .S(\SUMB[17][31] ) );
  FA1A S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA1A S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA1A S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA1A S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA1A S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA1A S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA1A S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA1A S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA1A S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1A S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1A S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1A S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1A S2_14_63 ( .A(\ab[14][63] ), .B(\CARRYB[13][63] ), .CI(\SUMB[13][64] ), 
        .CO(\CARRYB[14][63] ), .S(\SUMB[14][63] ) );
  FA1A S2_14_62 ( .A(\ab[14][62] ), .B(\CARRYB[13][62] ), .CI(\SUMB[13][63] ), 
        .CO(\CARRYB[14][62] ), .S(\SUMB[14][62] ) );
  FA1A S2_14_61 ( .A(\ab[14][61] ), .B(\CARRYB[13][61] ), .CI(\SUMB[13][62] ), 
        .CO(\CARRYB[14][61] ), .S(\SUMB[14][61] ) );
  FA1A S2_16_36 ( .A(\ab[16][36] ), .B(\CARRYB[15][36] ), .CI(\SUMB[15][37] ), 
        .CO(\CARRYB[16][36] ), .S(\SUMB[16][36] ) );
  FA1A S2_16_35 ( .A(\ab[16][35] ), .B(\CARRYB[15][35] ), .CI(\SUMB[15][36] ), 
        .CO(\CARRYB[16][35] ), .S(\SUMB[16][35] ) );
  FA1A S2_16_34 ( .A(\ab[16][34] ), .B(\CARRYB[15][34] ), .CI(\SUMB[15][35] ), 
        .CO(\CARRYB[16][34] ), .S(\SUMB[16][34] ) );
  FA1A S2_16_33 ( .A(\ab[16][33] ), .B(\CARRYB[15][33] ), .CI(\SUMB[15][34] ), 
        .CO(\CARRYB[16][33] ), .S(\SUMB[16][33] ) );
  FA1A S2_16_32 ( .A(\ab[16][32] ), .B(\CARRYB[15][32] ), .CI(\SUMB[15][33] ), 
        .CO(\CARRYB[16][32] ), .S(\SUMB[16][32] ) );
  FA1A S2_16_31 ( .A(\ab[16][31] ), .B(\CARRYB[15][31] ), .CI(\SUMB[15][32] ), 
        .CO(\CARRYB[16][31] ), .S(\SUMB[16][31] ) );
  FA1A S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA1A S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA1A S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA1A S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA1A S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA1A S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA1A S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA1A S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA1A S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1A S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1A S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA1A S2_13_63 ( .A(\ab[13][63] ), .B(\CARRYB[12][63] ), .CI(\SUMB[12][64] ), 
        .CO(\CARRYB[13][63] ), .S(\SUMB[13][63] ) );
  FA1A S2_13_62 ( .A(\ab[13][62] ), .B(\CARRYB[12][62] ), .CI(\SUMB[12][63] ), 
        .CO(\CARRYB[13][62] ), .S(\SUMB[13][62] ) );
  FA1A S2_13_61 ( .A(\ab[13][61] ), .B(\CARRYB[12][61] ), .CI(\SUMB[12][62] ), 
        .CO(\CARRYB[13][61] ), .S(\SUMB[13][61] ) );
  FA1A S2_15_37 ( .A(\ab[15][37] ), .B(\CARRYB[14][37] ), .CI(\SUMB[14][38] ), 
        .CO(\CARRYB[15][37] ), .S(\SUMB[15][37] ) );
  FA1A S2_15_36 ( .A(\ab[15][36] ), .B(\CARRYB[14][36] ), .CI(\SUMB[14][37] ), 
        .CO(\CARRYB[15][36] ), .S(\SUMB[15][36] ) );
  FA1A S2_15_35 ( .A(\ab[15][35] ), .B(\CARRYB[14][35] ), .CI(\SUMB[14][36] ), 
        .CO(\CARRYB[15][35] ), .S(\SUMB[15][35] ) );
  FA1A S2_15_34 ( .A(\ab[15][34] ), .B(\CARRYB[14][34] ), .CI(\SUMB[14][35] ), 
        .CO(\CARRYB[15][34] ), .S(\SUMB[15][34] ) );
  FA1A S2_15_33 ( .A(\ab[15][33] ), .B(\CARRYB[14][33] ), .CI(\SUMB[14][34] ), 
        .CO(\CARRYB[15][33] ), .S(\SUMB[15][33] ) );
  FA1A S2_15_32 ( .A(\ab[15][32] ), .B(\CARRYB[14][32] ), .CI(\SUMB[14][33] ), 
        .CO(\CARRYB[15][32] ), .S(\SUMB[15][32] ) );
  FA1A S2_15_31 ( .A(\ab[15][31] ), .B(\CARRYB[14][31] ), .CI(\SUMB[14][32] ), 
        .CO(\CARRYB[15][31] ), .S(\SUMB[15][31] ) );
  FA1A S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA1A S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA1A S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA1A S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA1A S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA1A S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA1A S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA1A S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S2_12_63 ( .A(\ab[12][63] ), .B(\CARRYB[11][63] ), .CI(\SUMB[11][64] ), 
        .CO(\CARRYB[12][63] ), .S(\SUMB[12][63] ) );
  FA1A S2_12_62 ( .A(\ab[12][62] ), .B(\CARRYB[11][62] ), .CI(\SUMB[11][63] ), 
        .CO(\CARRYB[12][62] ), .S(\SUMB[12][62] ) );
  FA1A S2_12_61 ( .A(\ab[12][61] ), .B(\CARRYB[11][61] ), .CI(\SUMB[11][62] ), 
        .CO(\CARRYB[12][61] ), .S(\SUMB[12][61] ) );
  FA1A S2_14_37 ( .A(\ab[14][37] ), .B(\CARRYB[13][37] ), .CI(\SUMB[13][38] ), 
        .CO(\CARRYB[14][37] ), .S(\SUMB[14][37] ) );
  FA1A S2_14_36 ( .A(\ab[14][36] ), .B(\CARRYB[13][36] ), .CI(\SUMB[13][37] ), 
        .CO(\CARRYB[14][36] ), .S(\SUMB[14][36] ) );
  FA1A S2_14_35 ( .A(\ab[14][35] ), .B(\CARRYB[13][35] ), .CI(\SUMB[13][36] ), 
        .CO(\CARRYB[14][35] ), .S(\SUMB[14][35] ) );
  FA1A S2_14_34 ( .A(\ab[14][34] ), .B(\CARRYB[13][34] ), .CI(\SUMB[13][35] ), 
        .CO(\CARRYB[14][34] ), .S(\SUMB[14][34] ) );
  FA1A S2_14_33 ( .A(\ab[14][33] ), .B(\CARRYB[13][33] ), .CI(\SUMB[13][34] ), 
        .CO(\CARRYB[14][33] ), .S(\SUMB[14][33] ) );
  FA1A S2_14_32 ( .A(\ab[14][32] ), .B(\CARRYB[13][32] ), .CI(\SUMB[13][33] ), 
        .CO(\CARRYB[14][32] ), .S(\SUMB[14][32] ) );
  FA1A S2_14_31 ( .A(\ab[14][31] ), .B(\CARRYB[13][31] ), .CI(\SUMB[13][32] ), 
        .CO(\CARRYB[14][31] ), .S(\SUMB[14][31] ) );
  FA1A S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA1A S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA1A S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA1A S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA1A S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA1A S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA1A S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA1A S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_11_63 ( .A(\ab[11][63] ), .B(\CARRYB[10][63] ), .CI(\SUMB[10][64] ), 
        .CO(\CARRYB[11][63] ), .S(\SUMB[11][63] ) );
  FA1A S2_11_62 ( .A(\ab[11][62] ), .B(\CARRYB[10][62] ), .CI(\SUMB[10][63] ), 
        .CO(\CARRYB[11][62] ), .S(\SUMB[11][62] ) );
  FA1A S2_11_61 ( .A(\ab[11][61] ), .B(\CARRYB[10][61] ), .CI(\SUMB[10][62] ), 
        .CO(\CARRYB[11][61] ), .S(\SUMB[11][61] ) );
  FA1A S2_13_37 ( .A(\ab[13][37] ), .B(\CARRYB[12][37] ), .CI(\SUMB[12][38] ), 
        .CO(\CARRYB[13][37] ), .S(\SUMB[13][37] ) );
  FA1A S2_13_36 ( .A(\ab[13][36] ), .B(\CARRYB[12][36] ), .CI(\SUMB[12][37] ), 
        .CO(\CARRYB[13][36] ), .S(\SUMB[13][36] ) );
  FA1A S2_13_35 ( .A(\ab[13][35] ), .B(\CARRYB[12][35] ), .CI(\SUMB[12][36] ), 
        .CO(\CARRYB[13][35] ), .S(\SUMB[13][35] ) );
  FA1A S2_13_34 ( .A(\ab[13][34] ), .B(\CARRYB[12][34] ), .CI(\SUMB[12][35] ), 
        .CO(\CARRYB[13][34] ), .S(\SUMB[13][34] ) );
  FA1A S2_13_33 ( .A(\ab[13][33] ), .B(\CARRYB[12][33] ), .CI(\SUMB[12][34] ), 
        .CO(\CARRYB[13][33] ), .S(\SUMB[13][33] ) );
  FA1A S2_13_32 ( .A(\ab[13][32] ), .B(\CARRYB[12][32] ), .CI(\SUMB[12][33] ), 
        .CO(\CARRYB[13][32] ), .S(\SUMB[13][32] ) );
  FA1A S2_13_31 ( .A(\ab[13][31] ), .B(\CARRYB[12][31] ), .CI(\SUMB[12][32] ), 
        .CO(\CARRYB[13][31] ), .S(\SUMB[13][31] ) );
  FA1A S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA1A S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA1A S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA1A S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA1A S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA1A S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA1A S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA1A S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_10_63 ( .A(\ab[10][63] ), .B(\CARRYB[9][63] ), .CI(\SUMB[9][64] ), 
        .CO(\CARRYB[10][63] ), .S(\SUMB[10][63] ) );
  FA1A S2_10_62 ( .A(\ab[10][62] ), .B(\CARRYB[9][62] ), .CI(\SUMB[9][63] ), 
        .CO(\CARRYB[10][62] ), .S(\SUMB[10][62] ) );
  FA1A S2_10_61 ( .A(\ab[10][61] ), .B(\CARRYB[9][61] ), .CI(\SUMB[9][62] ), 
        .CO(\CARRYB[10][61] ), .S(\SUMB[10][61] ) );
  FA1A S2_12_37 ( .A(\ab[12][37] ), .B(\CARRYB[11][37] ), .CI(\SUMB[11][38] ), 
        .CO(\CARRYB[12][37] ), .S(\SUMB[12][37] ) );
  FA1A S2_12_36 ( .A(\ab[12][36] ), .B(\CARRYB[11][36] ), .CI(\SUMB[11][37] ), 
        .CO(\CARRYB[12][36] ), .S(\SUMB[12][36] ) );
  FA1A S2_12_35 ( .A(\ab[12][35] ), .B(\CARRYB[11][35] ), .CI(\SUMB[11][36] ), 
        .CO(\CARRYB[12][35] ), .S(\SUMB[12][35] ) );
  FA1A S2_12_34 ( .A(\ab[12][34] ), .B(\CARRYB[11][34] ), .CI(\SUMB[11][35] ), 
        .CO(\CARRYB[12][34] ), .S(\SUMB[12][34] ) );
  FA1A S2_12_33 ( .A(\ab[12][33] ), .B(\CARRYB[11][33] ), .CI(\SUMB[11][34] ), 
        .CO(\CARRYB[12][33] ), .S(\SUMB[12][33] ) );
  FA1A S2_12_32 ( .A(\ab[12][32] ), .B(\CARRYB[11][32] ), .CI(\SUMB[11][33] ), 
        .CO(\CARRYB[12][32] ), .S(\SUMB[12][32] ) );
  FA1A S2_12_31 ( .A(\ab[12][31] ), .B(\CARRYB[11][31] ), .CI(\SUMB[11][32] ), 
        .CO(\CARRYB[12][31] ), .S(\SUMB[12][31] ) );
  FA1A S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA1A S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA1A S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA1A S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA1A S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA1A S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA1A S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA1A S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_9_63 ( .A(\ab[9][63] ), .B(\CARRYB[8][63] ), .CI(\SUMB[8][64] ), 
        .CO(\CARRYB[9][63] ), .S(\SUMB[9][63] ) );
  FA1A S2_9_62 ( .A(\ab[9][62] ), .B(\CARRYB[8][62] ), .CI(\SUMB[8][63] ), 
        .CO(\CARRYB[9][62] ), .S(\SUMB[9][62] ) );
  FA1A S2_9_61 ( .A(\ab[9][61] ), .B(\CARRYB[8][61] ), .CI(\SUMB[8][62] ), 
        .CO(\CARRYB[9][61] ), .S(\SUMB[9][61] ) );
  FA1A S2_11_37 ( .A(\ab[11][37] ), .B(\CARRYB[10][37] ), .CI(\SUMB[10][38] ), 
        .CO(\CARRYB[11][37] ), .S(\SUMB[11][37] ) );
  FA1A S2_11_36 ( .A(\ab[11][36] ), .B(\CARRYB[10][36] ), .CI(\SUMB[10][37] ), 
        .CO(\CARRYB[11][36] ), .S(\SUMB[11][36] ) );
  FA1A S2_11_35 ( .A(\ab[11][35] ), .B(\CARRYB[10][35] ), .CI(\SUMB[10][36] ), 
        .CO(\CARRYB[11][35] ), .S(\SUMB[11][35] ) );
  FA1A S2_11_34 ( .A(\ab[11][34] ), .B(\CARRYB[10][34] ), .CI(\SUMB[10][35] ), 
        .CO(\CARRYB[11][34] ), .S(\SUMB[11][34] ) );
  FA1A S2_11_33 ( .A(\ab[11][33] ), .B(\CARRYB[10][33] ), .CI(\SUMB[10][34] ), 
        .CO(\CARRYB[11][33] ), .S(\SUMB[11][33] ) );
  FA1A S2_11_32 ( .A(\ab[11][32] ), .B(\CARRYB[10][32] ), .CI(\SUMB[10][33] ), 
        .CO(\CARRYB[11][32] ), .S(\SUMB[11][32] ) );
  FA1A S2_11_31 ( .A(\ab[11][31] ), .B(\CARRYB[10][31] ), .CI(\SUMB[10][32] ), 
        .CO(\CARRYB[11][31] ), .S(\SUMB[11][31] ) );
  FA1A S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1A S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA1A S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1A S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1A S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1A S2_11_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1A S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1A S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_8_63 ( .A(\ab[8][63] ), .B(\CARRYB[7][63] ), .CI(\SUMB[7][64] ), 
        .CO(\CARRYB[8][63] ), .S(\SUMB[8][63] ) );
  FA1A S2_8_62 ( .A(\ab[8][62] ), .B(\CARRYB[7][62] ), .CI(\SUMB[7][63] ), 
        .CO(\CARRYB[8][62] ), .S(\SUMB[8][62] ) );
  FA1A S2_8_61 ( .A(\ab[8][61] ), .B(\CARRYB[7][61] ), .CI(\SUMB[7][62] ), 
        .CO(\CARRYB[8][61] ), .S(\SUMB[8][61] ) );
  FA1A S2_10_37 ( .A(\ab[10][37] ), .B(\CARRYB[9][37] ), .CI(\SUMB[9][38] ), 
        .CO(\CARRYB[10][37] ), .S(\SUMB[10][37] ) );
  FA1A S2_10_36 ( .A(\ab[10][36] ), .B(\CARRYB[9][36] ), .CI(\SUMB[9][37] ), 
        .CO(\CARRYB[10][36] ), .S(\SUMB[10][36] ) );
  FA1A S2_10_35 ( .A(\ab[10][35] ), .B(\CARRYB[9][35] ), .CI(\SUMB[9][36] ), 
        .CO(\CARRYB[10][35] ), .S(\SUMB[10][35] ) );
  FA1A S2_10_34 ( .A(\ab[10][34] ), .B(\CARRYB[9][34] ), .CI(\SUMB[9][35] ), 
        .CO(\CARRYB[10][34] ), .S(\SUMB[10][34] ) );
  FA1A S2_10_33 ( .A(\ab[10][33] ), .B(\CARRYB[9][33] ), .CI(\SUMB[9][34] ), 
        .CO(\CARRYB[10][33] ), .S(\SUMB[10][33] ) );
  FA1A S2_10_32 ( .A(\ab[10][32] ), .B(\CARRYB[9][32] ), .CI(\SUMB[9][33] ), 
        .CO(\CARRYB[10][32] ), .S(\SUMB[10][32] ) );
  FA1A S2_10_31 ( .A(\ab[10][31] ), .B(\CARRYB[9][31] ), .CI(\SUMB[9][32] ), 
        .CO(\CARRYB[10][31] ), .S(\SUMB[10][31] ) );
  FA1A S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1A S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA1A S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA1A S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1A S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1A S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA1A S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA1A S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_7_63 ( .A(\ab[7][63] ), .B(\CARRYB[6][63] ), .CI(\SUMB[6][64] ), 
        .CO(\CARRYB[7][63] ), .S(\SUMB[7][63] ) );
  FA1A S2_7_62 ( .A(\ab[7][62] ), .B(\CARRYB[6][62] ), .CI(\SUMB[6][63] ), 
        .CO(\CARRYB[7][62] ), .S(\SUMB[7][62] ) );
  FA1A S2_7_61 ( .A(\ab[7][61] ), .B(\CARRYB[6][61] ), .CI(\SUMB[6][62] ), 
        .CO(\CARRYB[7][61] ), .S(\SUMB[7][61] ) );
  FA1A S2_9_37 ( .A(\ab[9][37] ), .B(\CARRYB[8][37] ), .CI(\SUMB[8][38] ), 
        .CO(\CARRYB[9][37] ), .S(\SUMB[9][37] ) );
  FA1A S2_9_36 ( .A(\ab[9][36] ), .B(\CARRYB[8][36] ), .CI(\SUMB[8][37] ), 
        .CO(\CARRYB[9][36] ), .S(\SUMB[9][36] ) );
  FA1A S2_9_35 ( .A(\ab[9][35] ), .B(\CARRYB[8][35] ), .CI(\SUMB[8][36] ), 
        .CO(\CARRYB[9][35] ), .S(\SUMB[9][35] ) );
  FA1A S2_9_34 ( .A(\ab[9][34] ), .B(\CARRYB[8][34] ), .CI(\SUMB[8][35] ), 
        .CO(\CARRYB[9][34] ), .S(\SUMB[9][34] ) );
  FA1A S2_9_33 ( .A(\ab[9][33] ), .B(\CARRYB[8][33] ), .CI(\SUMB[8][34] ), 
        .CO(\CARRYB[9][33] ), .S(\SUMB[9][33] ) );
  FA1A S2_9_32 ( .A(\ab[9][32] ), .B(\CARRYB[8][32] ), .CI(\SUMB[8][33] ), 
        .CO(\CARRYB[9][32] ), .S(\SUMB[9][32] ) );
  FA1A S2_9_31 ( .A(\ab[9][31] ), .B(\CARRYB[8][31] ), .CI(\SUMB[8][32] ), 
        .CO(\CARRYB[9][31] ), .S(\SUMB[9][31] ) );
  FA1A S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1A S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1A S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1A S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1A S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1A S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA1A S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_6_63 ( .A(\ab[6][63] ), .B(\CARRYB[5][63] ), .CI(\SUMB[5][64] ), 
        .CO(\CARRYB[6][63] ), .S(\SUMB[6][63] ) );
  FA1A S2_6_62 ( .A(\ab[6][62] ), .B(\CARRYB[5][62] ), .CI(\SUMB[5][63] ), 
        .CO(\CARRYB[6][62] ), .S(\SUMB[6][62] ) );
  FA1A S2_6_61 ( .A(\ab[6][61] ), .B(\CARRYB[5][61] ), .CI(\SUMB[5][62] ), 
        .CO(\CARRYB[6][61] ), .S(\SUMB[6][61] ) );
  FA1A S2_8_37 ( .A(\ab[8][37] ), .B(\CARRYB[7][37] ), .CI(\SUMB[7][38] ), 
        .CO(\CARRYB[8][37] ), .S(\SUMB[8][37] ) );
  FA1A S2_8_36 ( .A(\ab[8][36] ), .B(\CARRYB[7][36] ), .CI(\SUMB[7][37] ), 
        .CO(\CARRYB[8][36] ), .S(\SUMB[8][36] ) );
  FA1A S2_8_35 ( .A(\ab[8][35] ), .B(\CARRYB[7][35] ), .CI(\SUMB[7][36] ), 
        .CO(\CARRYB[8][35] ), .S(\SUMB[8][35] ) );
  FA1A S2_8_34 ( .A(\ab[8][34] ), .B(\CARRYB[7][34] ), .CI(\SUMB[7][35] ), 
        .CO(\CARRYB[8][34] ), .S(\SUMB[8][34] ) );
  FA1A S2_8_33 ( .A(\ab[8][33] ), .B(\CARRYB[7][33] ), .CI(\SUMB[7][34] ), 
        .CO(\CARRYB[8][33] ), .S(\SUMB[8][33] ) );
  FA1A S2_8_32 ( .A(\ab[8][32] ), .B(\CARRYB[7][32] ), .CI(\SUMB[7][33] ), 
        .CO(\CARRYB[8][32] ), .S(\SUMB[8][32] ) );
  FA1A S2_8_31 ( .A(\ab[8][31] ), .B(\CARRYB[7][31] ), .CI(\SUMB[7][32] ), 
        .CO(\CARRYB[8][31] ), .S(\SUMB[8][31] ) );
  FA1A S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA1A S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1A S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1A S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1A S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1A S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1A S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1A S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_5_63 ( .A(\ab[5][63] ), .B(\CARRYB[4][63] ), .CI(\SUMB[4][64] ), 
        .CO(\CARRYB[5][63] ), .S(\SUMB[5][63] ) );
  FA1A S2_5_62 ( .A(\ab[5][62] ), .B(\CARRYB[4][62] ), .CI(\SUMB[4][63] ), 
        .CO(\CARRYB[5][62] ), .S(\SUMB[5][62] ) );
  FA1A S2_5_61 ( .A(\ab[5][61] ), .B(\CARRYB[4][61] ), .CI(\SUMB[4][62] ), 
        .CO(\CARRYB[5][61] ), .S(\SUMB[5][61] ) );
  FA1A S2_7_37 ( .A(\ab[7][37] ), .B(\CARRYB[6][37] ), .CI(\SUMB[6][38] ), 
        .CO(\CARRYB[7][37] ), .S(\SUMB[7][37] ) );
  FA1A S2_7_36 ( .A(\ab[7][36] ), .B(\CARRYB[6][36] ), .CI(\SUMB[6][37] ), 
        .CO(\CARRYB[7][36] ), .S(\SUMB[7][36] ) );
  FA1A S2_7_35 ( .A(\ab[7][35] ), .B(\CARRYB[6][35] ), .CI(\SUMB[6][36] ), 
        .CO(\CARRYB[7][35] ), .S(\SUMB[7][35] ) );
  FA1A S2_7_34 ( .A(\ab[7][34] ), .B(\CARRYB[6][34] ), .CI(\SUMB[6][35] ), 
        .CO(\CARRYB[7][34] ), .S(\SUMB[7][34] ) );
  FA1A S2_7_33 ( .A(\ab[7][33] ), .B(\CARRYB[6][33] ), .CI(\SUMB[6][34] ), 
        .CO(\CARRYB[7][33] ), .S(\SUMB[7][33] ) );
  FA1A S2_7_32 ( .A(\ab[7][32] ), .B(\CARRYB[6][32] ), .CI(\SUMB[6][33] ), 
        .CO(\CARRYB[7][32] ), .S(\SUMB[7][32] ) );
  FA1A S2_7_31 ( .A(\ab[7][31] ), .B(\CARRYB[6][31] ), .CI(\SUMB[6][32] ), 
        .CO(\CARRYB[7][31] ), .S(\SUMB[7][31] ) );
  FA1A S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA1A S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1A S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA1A S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA1A S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA1A S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA1A S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA1A S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_4_63 ( .A(\ab[4][63] ), .B(\CARRYB[3][63] ), .CI(\SUMB[3][64] ), 
        .CO(\CARRYB[4][63] ), .S(\SUMB[4][63] ) );
  FA1A S2_4_62 ( .A(\ab[4][62] ), .B(\CARRYB[3][62] ), .CI(\SUMB[3][63] ), 
        .CO(\CARRYB[4][62] ), .S(\SUMB[4][62] ) );
  FA1A S2_4_61 ( .A(\ab[4][61] ), .B(\CARRYB[3][61] ), .CI(\SUMB[3][62] ), 
        .CO(\CARRYB[4][61] ), .S(\SUMB[4][61] ) );
  FA1A S2_6_37 ( .A(\ab[6][37] ), .B(\CARRYB[5][37] ), .CI(\SUMB[5][38] ), 
        .CO(\CARRYB[6][37] ), .S(\SUMB[6][37] ) );
  FA1A S2_6_36 ( .A(\ab[6][36] ), .B(\CARRYB[5][36] ), .CI(\SUMB[5][37] ), 
        .CO(\CARRYB[6][36] ), .S(\SUMB[6][36] ) );
  FA1A S2_6_35 ( .A(\ab[6][35] ), .B(\CARRYB[5][35] ), .CI(\SUMB[5][36] ), 
        .CO(\CARRYB[6][35] ), .S(\SUMB[6][35] ) );
  FA1A S2_6_34 ( .A(\ab[6][34] ), .B(\CARRYB[5][34] ), .CI(\SUMB[5][35] ), 
        .CO(\CARRYB[6][34] ), .S(\SUMB[6][34] ) );
  FA1A S2_6_33 ( .A(\ab[6][33] ), .B(\CARRYB[5][33] ), .CI(\SUMB[5][34] ), 
        .CO(\CARRYB[6][33] ), .S(\SUMB[6][33] ) );
  FA1A S2_6_32 ( .A(\ab[6][32] ), .B(\CARRYB[5][32] ), .CI(\SUMB[5][33] ), 
        .CO(\CARRYB[6][32] ), .S(\SUMB[6][32] ) );
  FA1A S2_6_31 ( .A(\ab[6][31] ), .B(\CARRYB[5][31] ), .CI(\SUMB[5][32] ), 
        .CO(\CARRYB[6][31] ), .S(\SUMB[6][31] ) );
  FA1A S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1A S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA1A S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA1A S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA1A S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1A S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1A S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA1A S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_3_63 ( .A(\ab[3][63] ), .B(\CARRYB[2][63] ), .CI(\SUMB[2][64] ), 
        .CO(\CARRYB[3][63] ), .S(\SUMB[3][63] ) );
  FA1A S2_3_62 ( .A(\ab[3][62] ), .B(\CARRYB[2][62] ), .CI(\SUMB[2][63] ), 
        .CO(\CARRYB[3][62] ), .S(\SUMB[3][62] ) );
  FA1A S2_3_61 ( .A(\ab[3][61] ), .B(\CARRYB[2][61] ), .CI(\SUMB[2][62] ), 
        .CO(\CARRYB[3][61] ), .S(\SUMB[3][61] ) );
  FA1A S2_5_37 ( .A(\ab[5][37] ), .B(\CARRYB[4][37] ), .CI(\SUMB[4][38] ), 
        .CO(\CARRYB[5][37] ), .S(\SUMB[5][37] ) );
  FA1A S2_5_36 ( .A(\ab[5][36] ), .B(\CARRYB[4][36] ), .CI(\SUMB[4][37] ), 
        .CO(\CARRYB[5][36] ), .S(\SUMB[5][36] ) );
  FA1A S2_5_35 ( .A(\ab[5][35] ), .B(\CARRYB[4][35] ), .CI(\SUMB[4][36] ), 
        .CO(\CARRYB[5][35] ), .S(\SUMB[5][35] ) );
  FA1A S2_5_34 ( .A(\ab[5][34] ), .B(\CARRYB[4][34] ), .CI(\SUMB[4][35] ), 
        .CO(\CARRYB[5][34] ), .S(\SUMB[5][34] ) );
  FA1A S2_5_33 ( .A(\ab[5][33] ), .B(\CARRYB[4][33] ), .CI(\SUMB[4][34] ), 
        .CO(\CARRYB[5][33] ), .S(\SUMB[5][33] ) );
  FA1A S2_5_32 ( .A(\ab[5][32] ), .B(\CARRYB[4][32] ), .CI(\SUMB[4][33] ), 
        .CO(\CARRYB[5][32] ), .S(\SUMB[5][32] ) );
  FA1A S2_5_31 ( .A(\ab[5][31] ), .B(\CARRYB[4][31] ), .CI(\SUMB[4][32] ), 
        .CO(\CARRYB[5][31] ), .S(\SUMB[5][31] ) );
  FA1A S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA1A S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA1A S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1A S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1A S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1A S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1A S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_2_63 ( .A(\ab[2][63] ), .B(\CARRYB[1][63] ), .CI(\SUMB[1][64] ), 
        .CO(\CARRYB[2][63] ), .S(\SUMB[2][63] ) );
  FA1A S2_2_62 ( .A(\ab[2][62] ), .B(\CARRYB[1][62] ), .CI(\SUMB[1][63] ), 
        .CO(\CARRYB[2][62] ), .S(\SUMB[2][62] ) );
  FA1A S2_2_61 ( .A(\ab[2][61] ), .B(\CARRYB[1][61] ), .CI(\SUMB[1][62] ), 
        .CO(\CARRYB[2][61] ), .S(\SUMB[2][61] ) );
  FA1A S2_4_37 ( .A(\ab[4][37] ), .B(\CARRYB[3][37] ), .CI(\SUMB[3][38] ), 
        .CO(\CARRYB[4][37] ), .S(\SUMB[4][37] ) );
  FA1A S2_4_36 ( .A(\ab[4][36] ), .B(\CARRYB[3][36] ), .CI(\SUMB[3][37] ), 
        .CO(\CARRYB[4][36] ), .S(\SUMB[4][36] ) );
  FA1A S2_4_35 ( .A(\ab[4][35] ), .B(\CARRYB[3][35] ), .CI(\SUMB[3][36] ), 
        .CO(\CARRYB[4][35] ), .S(\SUMB[4][35] ) );
  FA1A S2_4_34 ( .A(\ab[4][34] ), .B(\CARRYB[3][34] ), .CI(\SUMB[3][35] ), 
        .CO(\CARRYB[4][34] ), .S(\SUMB[4][34] ) );
  FA1A S2_4_33 ( .A(\ab[4][33] ), .B(\CARRYB[3][33] ), .CI(\SUMB[3][34] ), 
        .CO(\CARRYB[4][33] ), .S(\SUMB[4][33] ) );
  FA1A S2_4_32 ( .A(\ab[4][32] ), .B(\CARRYB[3][32] ), .CI(\SUMB[3][33] ), 
        .CO(\CARRYB[4][32] ), .S(\SUMB[4][32] ) );
  FA1A S2_4_31 ( .A(\ab[4][31] ), .B(\CARRYB[3][31] ), .CI(\SUMB[3][32] ), 
        .CO(\CARRYB[4][31] ), .S(\SUMB[4][31] ) );
  FA1A S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1A S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1A S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1A S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1A S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1A S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA1A S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA1A S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_3_37 ( .A(\ab[3][37] ), .B(\CARRYB[2][37] ), .CI(\SUMB[2][38] ), 
        .CO(\CARRYB[3][37] ), .S(\SUMB[3][37] ) );
  FA1A S2_3_36 ( .A(\ab[3][36] ), .B(\CARRYB[2][36] ), .CI(\SUMB[2][37] ), 
        .CO(\CARRYB[3][36] ), .S(\SUMB[3][36] ) );
  FA1A S2_3_35 ( .A(\ab[3][35] ), .B(\CARRYB[2][35] ), .CI(\SUMB[2][36] ), 
        .CO(\CARRYB[3][35] ), .S(\SUMB[3][35] ) );
  FA1A S2_3_34 ( .A(\ab[3][34] ), .B(\CARRYB[2][34] ), .CI(\SUMB[2][35] ), 
        .CO(\CARRYB[3][34] ), .S(\SUMB[3][34] ) );
  FA1A S2_3_33 ( .A(\ab[3][33] ), .B(\CARRYB[2][33] ), .CI(\SUMB[2][34] ), 
        .CO(\CARRYB[3][33] ), .S(\SUMB[3][33] ) );
  FA1A S2_3_32 ( .A(\ab[3][32] ), .B(\CARRYB[2][32] ), .CI(\SUMB[2][33] ), 
        .CO(\CARRYB[3][32] ), .S(\SUMB[3][32] ) );
  FA1A S2_3_31 ( .A(\ab[3][31] ), .B(\CARRYB[2][31] ), .CI(\SUMB[2][32] ), 
        .CO(\CARRYB[3][31] ), .S(\SUMB[3][31] ) );
  FA1A S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA1A S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1A S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1A S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA1A S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA1A S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA1A S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA1A S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_2_36 ( .A(\ab[2][36] ), .B(\CARRYB[1][36] ), .CI(\SUMB[1][37] ), 
        .CO(\CARRYB[2][36] ), .S(\SUMB[2][36] ) );
  FA1A S2_2_35 ( .A(\ab[2][35] ), .B(\CARRYB[1][35] ), .CI(\SUMB[1][36] ), 
        .CO(\CARRYB[2][35] ), .S(\SUMB[2][35] ) );
  FA1A S2_2_34 ( .A(\ab[2][34] ), .B(\CARRYB[1][34] ), .CI(\SUMB[1][35] ), 
        .CO(\CARRYB[2][34] ), .S(\SUMB[2][34] ) );
  FA1A S2_2_33 ( .A(\ab[2][33] ), .B(\CARRYB[1][33] ), .CI(\SUMB[1][34] ), 
        .CO(\CARRYB[2][33] ), .S(\SUMB[2][33] ) );
  FA1A S2_2_32 ( .A(\ab[2][32] ), .B(\CARRYB[1][32] ), .CI(\SUMB[1][33] ), 
        .CO(\CARRYB[2][32] ), .S(\SUMB[2][32] ) );
  FA1A S2_2_31 ( .A(\ab[2][31] ), .B(\CARRYB[1][31] ), .CI(\SUMB[1][32] ), 
        .CO(\CARRYB[2][31] ), .S(\SUMB[2][31] ) );
  FA1A S2_2_28 ( .A(\ab[2][28] ), .B(\CARRYB[1][28] ), .CI(\SUMB[1][29] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FA1A S2_2_27 ( .A(\ab[2][27] ), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1A S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1A S2_2_25 ( .A(\ab[2][25] ), .B(\CARRYB[1][25] ), .CI(\SUMB[1][26] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1A S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), 
        .CO(\CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA1A S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1A S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA1A S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), 
        .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA1A S4_32 ( .A(\ab[29][32] ), .B(\CARRYB[28][32] ), .CI(\SUMB[28][33] ), 
        .CO(\CARRYB[29][32] ), .S(\SUMB[29][32] ) );
  FA1A S4_36 ( .A(\ab[29][36] ), .B(\CARRYB[28][36] ), .CI(\SUMB[28][37] ), 
        .CO(\CARRYB[29][36] ), .S(\SUMB[29][36] ) );
  FA1A S4_35 ( .A(\ab[29][35] ), .B(\CARRYB[28][35] ), .CI(\SUMB[28][36] ), 
        .CO(\CARRYB[29][35] ), .S(\SUMB[29][35] ) );
  FA1A S4_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA1A S4_3 ( .A(\ab[29][3] ), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), .CO(
        \CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA1A S4_38 ( .A(\ab[29][38] ), .B(\CARRYB[28][38] ), .CI(\SUMB[28][39] ), 
        .CO(\CARRYB[29][38] ), .S(\SUMB[29][38] ) );
  FA1A S4_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA1A S4_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), .CO(
        \CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA1A S4_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), 
        .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FA1A S4_6 ( .A(\ab[29][6] ), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), .CO(
        \CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA1A S4_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), 
        .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA1A S4_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA1A S4_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA1A S4_5 ( .A(\ab[29][5] ), .B(\CARRYB[28][5] ), .CI(\SUMB[28][6] ), .CO(
        \CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA1A S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA1A S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), 
        .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA1A S2_28_12 ( .A(\ab[28][12] ), .B(\CARRYB[27][12] ), .CI(\SUMB[27][13] ), 
        .CO(\CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA1A S2_28_5 ( .A(\ab[28][5] ), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA1A S4_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA1A S4_14 ( .A(\ab[29][14] ), .B(\CARRYB[28][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA1A S4_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), 
        .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA1A S4_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA1A S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), 
        .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA1A S2_27_5 ( .A(\ab[27][5] ), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA1A S4_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), .CO(
        \CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA1A S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA1A S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA1A S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA1A S2_28_14 ( .A(\ab[28][14] ), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA1A S2_28_13 ( .A(\ab[28][13] ), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), 
        .CO(\CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA1A S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA1A S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA1A S2_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA1A S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA1A S2_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\SUMB[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA1A S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA1A S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA1A S2_27_15 ( .A(\ab[27][15] ), .B(\CARRYB[26][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA1A S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA1A S2_27_13 ( .A(\ab[27][13] ), .B(\CARRYB[26][13] ), .CI(\SUMB[26][14] ), 
        .CO(\CARRYB[27][13] ), .S(\SUMB[27][13] ) );
  FA1A S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA1A S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA1A S2_27_11 ( .A(\ab[27][11] ), .B(\CARRYB[26][11] ), .CI(\SUMB[26][12] ), 
        .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FA1A S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA1A S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA1A S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA1A S2_26_18 ( .A(\ab[26][18] ), .B(\CARRYB[25][18] ), .CI(\SUMB[25][19] ), 
        .CO(\CARRYB[26][18] ), .S(\SUMB[26][18] ) );
  FA1A S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA1A S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA1A S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA1A S2_26_14 ( .A(\ab[26][14] ), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), 
        .CO(\CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA1A S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), 
        .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA1A S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA1A S2_26_12 ( .A(\ab[26][12] ), .B(\CARRYB[25][12] ), .CI(\SUMB[25][13] ), 
        .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FA1A S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), 
        .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA1A S2_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA1A S2_26_9 ( .A(\ab[26][9] ), .B(\CARRYB[25][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA1A S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA1A S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA1A S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA1A S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA1A S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA1A S2_25_14 ( .A(\ab[25][14] ), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), 
        .CO(\CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA1A S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA1A S2_25_13 ( .A(\ab[25][13] ), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), 
        .CO(\CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA1A S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), 
        .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA1A S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), 
        .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA1A S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA1A S2_25_9 ( .A(\ab[25][9] ), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA1A S2_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\SUMB[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA1A S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA1A S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA1A S2_24_16 ( .A(\ab[24][16] ), .B(\CARRYB[23][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA1A S2_24_15 ( .A(\ab[24][15] ), .B(\CARRYB[23][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA1A S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA1A S2_24_14 ( .A(\ab[24][14] ), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), 
        .CO(\CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA1A S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), 
        .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA1A S2_24_12 ( .A(\ab[24][12] ), .B(\CARRYB[23][12] ), .CI(\SUMB[23][13] ), 
        .CO(\CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA1A S2_24_11 ( .A(\ab[24][11] ), .B(\CARRYB[23][11] ), .CI(\SUMB[23][12] ), 
        .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA1A S2_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA1A S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA1A S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA1A S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA1A S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA1A S2_23_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA1A S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1A S2_23_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA1A S2_23_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA1A S2_23_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA1A S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA1A S2_23_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA1A S2_23_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA1A S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA1A S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA1A S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA1A S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA1A S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA1A S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA1A S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA1A S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA1A S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA1A S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA1A S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA1A S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA1A S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA1A S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA1A S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA1A S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1A S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA1A S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA1A S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA1A S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA1A S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA1A S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA1A S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA1A S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1A S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1A S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA1A S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1A S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA1A S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA1A S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA1A S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA1A S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA1A S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA1A S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA1A S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA1A S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA1A S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1A S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA1A S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1A S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA1A S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA1A S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA1A S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA1A S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA1A S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA1A S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA1A S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA1A S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA1A S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA1A S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1A S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA1A S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA1A S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA1A S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA1A S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA1A S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA1A S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA1A S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA1A S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA1A S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA1A S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA1A S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1A S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA1A S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA1A S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA1A S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA1A S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA1A S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA1A S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA1A S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA1A S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA1A S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA1A S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1A S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA1A S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA1A S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA1A S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA1A S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA1A S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA1A S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA1A S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA1A S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA1A S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1A S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA1A S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA1A S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA1A S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA1A S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA1A S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA1A S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA1A S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA1A S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA1A S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1A S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA1A S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA1A S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA1A S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA1A S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA1A S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA1A S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA1A S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA1A S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA1A S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA1A S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA1A S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA1A S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1A S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1A S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1A S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1A S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1A S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1A S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1A S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1A S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1A S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1A S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1A S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1A S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA1A S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1A S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1A S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1A S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA1A S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1A S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1A S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1A S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1A S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1A S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1A S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1A S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1A S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1A S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1A S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA1A S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1A S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1A S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1A S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1A S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1A S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1A S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1A S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1A S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1A S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1A S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S4_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA1A S4_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA1A S4_12 ( .A(\ab[29][12] ), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), 
        .CO(\CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA1A S4_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA1A S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA1A S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA1A S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA1A S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA1A S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA1A S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA1A S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA1A S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA1A S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA1A S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA1A S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA1A S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA1A S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA1A S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA1A S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA1A S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA1A S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA1A S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1A S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1A S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1A S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA1A S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1A S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1A S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA1A S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1A S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  AN2P U2 ( .A(n173), .B(n305), .Z(n3) );
  IVDA U3 ( .A(n557), .Z(n4) );
  IVP U4 ( .A(A[22]), .Z(n557) );
  IVP U5 ( .A(n10), .Z(n8) );
  IVP U6 ( .A(n10), .Z(n9) );
  IVP U7 ( .A(n10), .Z(n7) );
  IVP U8 ( .A(n10), .Z(n6) );
  IVP U9 ( .A(n10), .Z(n5) );
  IVP U10 ( .A(n181), .Z(n174) );
  IVP U11 ( .A(n172), .Z(n165) );
  IVP U12 ( .A(n181), .Z(n176) );
  IVP U13 ( .A(n181), .Z(n177) );
  IVP U14 ( .A(n181), .Z(n173) );
  IVP U15 ( .A(n172), .Z(n164) );
  IVP U16 ( .A(n181), .Z(n175) );
  IVP U17 ( .A(n172), .Z(n167) );
  IVP U18 ( .A(n190), .Z(n183) );
  IVP U19 ( .A(n190), .Z(n185) );
  IVP U20 ( .A(n172), .Z(n168) );
  IVP U21 ( .A(n181), .Z(n178) );
  IVP U22 ( .A(n190), .Z(n186) );
  IVP U23 ( .A(n190), .Z(n182) );
  IVP U24 ( .A(n172), .Z(n166) );
  IVP U25 ( .A(n190), .Z(n184) );
  IVP U26 ( .A(n172), .Z(n169) );
  IVP U27 ( .A(n199), .Z(n192) );
  IVP U28 ( .A(n181), .Z(n179) );
  IVP U29 ( .A(n190), .Z(n187) );
  IVP U30 ( .A(n199), .Z(n193) );
  IVP U31 ( .A(n199), .Z(n194) );
  IVP U32 ( .A(n172), .Z(n170) );
  IVP U33 ( .A(n199), .Z(n191) );
  IVP U34 ( .A(n190), .Z(n188) );
  IVP U35 ( .A(n199), .Z(n195) );
  IVP U36 ( .A(n181), .Z(n180) );
  IVP U37 ( .A(n208), .Z(n201) );
  IVP U38 ( .A(n199), .Z(n196) );
  IVP U39 ( .A(n172), .Z(n171) );
  IVP U40 ( .A(n208), .Z(n203) );
  IVP U41 ( .A(n208), .Z(n204) );
  IVP U42 ( .A(n190), .Z(n189) );
  IVP U43 ( .A(n208), .Z(n200) );
  IVP U44 ( .A(n208), .Z(n202) );
  IVP U45 ( .A(n199), .Z(n197) );
  IVP U46 ( .A(n208), .Z(n205) );
  IVP U47 ( .A(n217), .Z(n210) );
  IVP U48 ( .A(n199), .Z(n198) );
  IVP U49 ( .A(n217), .Z(n211) );
  IVP U50 ( .A(n217), .Z(n212) );
  IVP U51 ( .A(n217), .Z(n209) );
  IVP U52 ( .A(n208), .Z(n206) );
  IVP U53 ( .A(n217), .Z(n213) );
  IVP U54 ( .A(n226), .Z(n219) );
  IVP U55 ( .A(n217), .Z(n214) );
  IVP U56 ( .A(n208), .Z(n207) );
  IVP U57 ( .A(n226), .Z(n221) );
  IVP U58 ( .A(n226), .Z(n222) );
  IVP U59 ( .A(n226), .Z(n218) );
  IVP U60 ( .A(n226), .Z(n220) );
  IVP U61 ( .A(n235), .Z(n228) );
  IVP U62 ( .A(n235), .Z(n230) );
  IVP U63 ( .A(n217), .Z(n215) );
  IVP U64 ( .A(n235), .Z(n227) );
  IVP U65 ( .A(n226), .Z(n223) );
  IVP U66 ( .A(n235), .Z(n231) );
  IVP U67 ( .A(n235), .Z(n229) );
  IVP U68 ( .A(n217), .Z(n216) );
  IVP U69 ( .A(n244), .Z(n237) );
  IVP U70 ( .A(n226), .Z(n224) );
  IVP U71 ( .A(n235), .Z(n232) );
  IVP U72 ( .A(n244), .Z(n239) );
  IVP U73 ( .A(n235), .Z(n233) );
  IVP U74 ( .A(n244), .Z(n240) );
  IVP U75 ( .A(n226), .Z(n225) );
  IVP U76 ( .A(n244), .Z(n236) );
  IVP U77 ( .A(n244), .Z(n238) );
  IVP U78 ( .A(n244), .Z(n241) );
  IVP U79 ( .A(n253), .Z(n246) );
  IVP U80 ( .A(n235), .Z(n234) );
  IVP U81 ( .A(n253), .Z(n245) );
  IVP U82 ( .A(n253), .Z(n248) );
  IVP U83 ( .A(n244), .Z(n242) );
  IVP U84 ( .A(n253), .Z(n249) );
  IVP U85 ( .A(n253), .Z(n247) );
  IVP U86 ( .A(n262), .Z(n255) );
  IVP U87 ( .A(n253), .Z(n250) );
  IVP U88 ( .A(n244), .Z(n243) );
  IVP U89 ( .A(n262), .Z(n254) );
  IVP U90 ( .A(n262), .Z(n256) );
  IVP U91 ( .A(n262), .Z(n257) );
  IVP U92 ( .A(n262), .Z(n258) );
  IVP U93 ( .A(n271), .Z(n264) );
  IVP U94 ( .A(n253), .Z(n251) );
  IVP U95 ( .A(n262), .Z(n259) );
  IVP U96 ( .A(n271), .Z(n263) );
  IVP U97 ( .A(n262), .Z(n260) );
  IVP U98 ( .A(n271), .Z(n266) );
  IVP U99 ( .A(n271), .Z(n267) );
  IVP U100 ( .A(n253), .Z(n252) );
  IVP U101 ( .A(n271), .Z(n265) );
  IVP U102 ( .A(n271), .Z(n268) );
  IVP U103 ( .A(n280), .Z(n273) );
  IVP U104 ( .A(n262), .Z(n261) );
  IVP U105 ( .A(n280), .Z(n274) );
  IVP U106 ( .A(n280), .Z(n275) );
  IVP U107 ( .A(n280), .Z(n276) );
  IVP U108 ( .A(n271), .Z(n269) );
  IVP U109 ( .A(n280), .Z(n272) );
  IVP U110 ( .A(n289), .Z(n282) );
  IVP U111 ( .A(n289), .Z(n281) );
  IVP U112 ( .A(n280), .Z(n277) );
  IVP U113 ( .A(n289), .Z(n285) );
  IVP U114 ( .A(n271), .Z(n270) );
  IVP U115 ( .A(n289), .Z(n283) );
  IVP U116 ( .A(n289), .Z(n284) );
  IVP U117 ( .A(n289), .Z(n286) );
  IVP U118 ( .A(n280), .Z(n278) );
  IVP U119 ( .A(n298), .Z(n291) );
  IVP U120 ( .A(n298), .Z(n293) );
  IVP U121 ( .A(n298), .Z(n294) );
  IVP U122 ( .A(n289), .Z(n287) );
  IVP U123 ( .A(n280), .Z(n279) );
  IVP U124 ( .A(n298), .Z(n290) );
  IVP U125 ( .A(n298), .Z(n292) );
  IVP U126 ( .A(n549), .Z(n10) );
  IVP U127 ( .A(n298), .Z(n295) );
  IVP U128 ( .A(n289), .Z(n288) );
  IVP U129 ( .A(n549), .Z(n13) );
  IVP U130 ( .A(n298), .Z(n296) );
  IVP U131 ( .A(n549), .Z(n12) );
  IVP U132 ( .A(n549), .Z(n14) );
  IVP U133 ( .A(n549), .Z(n15) );
  IVP U134 ( .A(n158), .Z(n156) );
  IVP U135 ( .A(n549), .Z(n11) );
  IVP U136 ( .A(n298), .Z(n297) );
  IVP U137 ( .A(n158), .Z(n157) );
  IVP U138 ( .A(n158), .Z(n155) );
  IVP U139 ( .A(n158), .Z(n154) );
  IVP U140 ( .A(n147), .Z(n145) );
  IVP U141 ( .A(n147), .Z(n146) );
  IVP U142 ( .A(n147), .Z(n144) );
  IVP U143 ( .A(n136), .Z(n134) );
  IVP U144 ( .A(n158), .Z(n153) );
  IVP U145 ( .A(n136), .Z(n135) );
  IVP U146 ( .A(n147), .Z(n143) );
  IVP U147 ( .A(n136), .Z(n133) );
  IVP U148 ( .A(n125), .Z(n123) );
  IVP U149 ( .A(n136), .Z(n132) );
  IVP U150 ( .A(n147), .Z(n142) );
  IVP U151 ( .A(n125), .Z(n124) );
  IVP U152 ( .A(n125), .Z(n122) );
  IVP U153 ( .A(n125), .Z(n121) );
  IVP U154 ( .A(n114), .Z(n112) );
  IVP U155 ( .A(n136), .Z(n131) );
  IVP U156 ( .A(n114), .Z(n113) );
  IVP U157 ( .A(n114), .Z(n111) );
  IVP U158 ( .A(n125), .Z(n120) );
  IVP U159 ( .A(n103), .Z(n101) );
  IVP U160 ( .A(n114), .Z(n110) );
  IVP U161 ( .A(n103), .Z(n102) );
  IVP U162 ( .A(n103), .Z(n100) );
  IVP U163 ( .A(n114), .Z(n109) );
  IVP U164 ( .A(n103), .Z(n99) );
  IVP U165 ( .A(n103), .Z(n98) );
  IVP U166 ( .A(n87), .Z(n85) );
  IVP U167 ( .A(n87), .Z(n86) );
  IVP U168 ( .A(n87), .Z(n84) );
  IVP U169 ( .A(n76), .Z(n74) );
  IVP U170 ( .A(n76), .Z(n75) );
  IVP U171 ( .A(n87), .Z(n83) );
  IVP U172 ( .A(n76), .Z(n73) );
  IVP U173 ( .A(n65), .Z(n63) );
  IVP U174 ( .A(n87), .Z(n82) );
  IVP U175 ( .A(n76), .Z(n72) );
  IVP U176 ( .A(n65), .Z(n64) );
  IVP U177 ( .A(n65), .Z(n62) );
  IVP U178 ( .A(n54), .Z(n52) );
  IVP U179 ( .A(n65), .Z(n61) );
  IVP U180 ( .A(n76), .Z(n71) );
  IVP U181 ( .A(n54), .Z(n53) );
  IVP U182 ( .A(n54), .Z(n51) );
  IVP U183 ( .A(n65), .Z(n60) );
  IVP U184 ( .A(n43), .Z(n41) );
  IVP U185 ( .A(n54), .Z(n50) );
  IVP U186 ( .A(n43), .Z(n42) );
  IVP U187 ( .A(n43), .Z(n40) );
  IVP U188 ( .A(n32), .Z(n30) );
  IVP U189 ( .A(n54), .Z(n49) );
  IVP U190 ( .A(n32), .Z(n31) );
  IVP U191 ( .A(n32), .Z(n29) );
  IVP U192 ( .A(n43), .Z(n39) );
  IVP U193 ( .A(n21), .Z(n19) );
  IVP U194 ( .A(n43), .Z(n38) );
  IVP U195 ( .A(n32), .Z(n28) );
  IVP U196 ( .A(n21), .Z(n20) );
  IVP U197 ( .A(n21), .Z(n18) );
  IVP U198 ( .A(n32), .Z(n27) );
  IVP U199 ( .A(n21), .Z(n17) );
  IVP U200 ( .A(n21), .Z(n16) );
  IVP U201 ( .A(A[1]), .Z(n181) );
  IVP U202 ( .A(A[0]), .Z(n172) );
  IVP U203 ( .A(A[2]), .Z(n190) );
  IVP U204 ( .A(A[3]), .Z(n199) );
  IVP U205 ( .A(A[4]), .Z(n208) );
  IVP U206 ( .A(A[5]), .Z(n217) );
  IVP U207 ( .A(A[6]), .Z(n226) );
  IVP U208 ( .A(A[7]), .Z(n235) );
  IVP U209 ( .A(A[8]), .Z(n244) );
  IVP U210 ( .A(A[9]), .Z(n253) );
  IVP U211 ( .A(A[10]), .Z(n262) );
  IVP U212 ( .A(A[11]), .Z(n271) );
  IVP U213 ( .A(A[12]), .Z(n280) );
  IVP U214 ( .A(A[13]), .Z(n289) );
  IVP U215 ( .A(A[14]), .Z(n298) );
  IVP U216 ( .A(A[15]), .Z(n549) );
  IVP U217 ( .A(n563), .Z(n158) );
  IVP U218 ( .A(n563), .Z(n161) );
  IVP U219 ( .A(n563), .Z(n162) );
  IVP U220 ( .A(n563), .Z(n160) );
  IVP U221 ( .A(n563), .Z(n159) );
  IVP U222 ( .A(n563), .Z(n163) );
  IVP U223 ( .A(n562), .Z(n147) );
  IVP U224 ( .A(n562), .Z(n150) );
  IVP U225 ( .A(n562), .Z(n151) );
  IVP U226 ( .A(n562), .Z(n149) );
  IVP U227 ( .A(n562), .Z(n148) );
  IVP U228 ( .A(n562), .Z(n152) );
  IVP U229 ( .A(n561), .Z(n136) );
  IVP U230 ( .A(n561), .Z(n139) );
  IVP U231 ( .A(n561), .Z(n140) );
  IVP U232 ( .A(n561), .Z(n138) );
  IVP U233 ( .A(n561), .Z(n137) );
  IVP U234 ( .A(n561), .Z(n141) );
  IVP U235 ( .A(n560), .Z(n125) );
  IVP U236 ( .A(n560), .Z(n129) );
  IVP U237 ( .A(n560), .Z(n128) );
  IVP U238 ( .A(n560), .Z(n127) );
  IVP U239 ( .A(n560), .Z(n126) );
  IVP U240 ( .A(n560), .Z(n130) );
  IVP U241 ( .A(n559), .Z(n114) );
  IVP U242 ( .A(n559), .Z(n118) );
  IVP U243 ( .A(n559), .Z(n117) );
  IVP U244 ( .A(n559), .Z(n116) );
  IVP U245 ( .A(n559), .Z(n115) );
  IVP U246 ( .A(n559), .Z(n119) );
  IVP U247 ( .A(n558), .Z(n103) );
  IVP U248 ( .A(n558), .Z(n107) );
  IVP U249 ( .A(n558), .Z(n106) );
  IVP U250 ( .A(n558), .Z(n105) );
  IVP U251 ( .A(n558), .Z(n104) );
  IVP U252 ( .A(n557), .Z(n96) );
  IVP U253 ( .A(n557), .Z(n95) );
  IVP U254 ( .A(n558), .Z(n108) );
  IVP U255 ( .A(n557), .Z(n94) );
  IVP U256 ( .A(n557), .Z(n93) );
  IVP U257 ( .A(n557), .Z(n97) );
  IVP U258 ( .A(n556), .Z(n87) );
  IVP U259 ( .A(n556), .Z(n91) );
  IVP U260 ( .A(n556), .Z(n90) );
  IVP U261 ( .A(n556), .Z(n89) );
  IVP U262 ( .A(n556), .Z(n88) );
  IVP U263 ( .A(n556), .Z(n92) );
  IVP U264 ( .A(n555), .Z(n76) );
  IVP U265 ( .A(n555), .Z(n80) );
  IVP U266 ( .A(n555), .Z(n79) );
  IVP U267 ( .A(n555), .Z(n78) );
  IVP U268 ( .A(n555), .Z(n77) );
  IVP U269 ( .A(n555), .Z(n81) );
  IVP U270 ( .A(n554), .Z(n65) );
  IVP U271 ( .A(n554), .Z(n68) );
  IVP U272 ( .A(n554), .Z(n69) );
  IVP U273 ( .A(n554), .Z(n70) );
  IVP U274 ( .A(n554), .Z(n67) );
  IVP U275 ( .A(n554), .Z(n66) );
  IVP U276 ( .A(n553), .Z(n54) );
  IVP U277 ( .A(n553), .Z(n57) );
  IVP U278 ( .A(n553), .Z(n56) );
  IVP U279 ( .A(n553), .Z(n58) );
  IVP U280 ( .A(n553), .Z(n59) );
  IVP U281 ( .A(n553), .Z(n55) );
  IVP U282 ( .A(n552), .Z(n43) );
  IVP U283 ( .A(n552), .Z(n47) );
  IVP U284 ( .A(n552), .Z(n46) );
  IVP U285 ( .A(n552), .Z(n45) );
  IVP U286 ( .A(n552), .Z(n44) );
  IVP U287 ( .A(n552), .Z(n48) );
  IVP U288 ( .A(n551), .Z(n32) );
  IVP U289 ( .A(n551), .Z(n36) );
  IVP U290 ( .A(n551), .Z(n35) );
  IVP U291 ( .A(n551), .Z(n34) );
  IVP U292 ( .A(n551), .Z(n33) );
  IVP U293 ( .A(n551), .Z(n37) );
  IVP U294 ( .A(n550), .Z(n21) );
  IVP U295 ( .A(n550), .Z(n24) );
  IVP U296 ( .A(n550), .Z(n25) );
  IVP U297 ( .A(n550), .Z(n23) );
  IVP U298 ( .A(n550), .Z(n22) );
  IVP U299 ( .A(n550), .Z(n26) );
  EO U300 ( .A(\CARRYB[29][19] ), .B(\SUMB[29][20] ), .Z(\A1[47] ) );
  EO U301 ( .A(\CARRYB[29][10] ), .B(\SUMB[29][11] ), .Z(\A1[38] ) );
  EO U302 ( .A(\CARRYB[29][15] ), .B(\SUMB[29][16] ), .Z(\A1[43] ) );
  EO U303 ( .A(\CARRYB[29][14] ), .B(\SUMB[29][15] ), .Z(\A1[42] ) );
  EO U304 ( .A(\CARRYB[29][5] ), .B(\SUMB[29][6] ), .Z(\A1[33] ) );
  EO U305 ( .A(\CARRYB[29][13] ), .B(\SUMB[29][14] ), .Z(\A1[41] ) );
  EO U306 ( .A(\CARRYB[29][9] ), .B(\SUMB[29][10] ), .Z(\A1[37] ) );
  EO U307 ( .A(\CARRYB[29][17] ), .B(\SUMB[29][18] ), .Z(\A1[45] ) );
  EO U308 ( .A(\CARRYB[29][18] ), .B(\SUMB[29][19] ), .Z(\A1[46] ) );
  EO U309 ( .A(\CARRYB[29][11] ), .B(\SUMB[29][12] ), .Z(\A1[39] ) );
  EO U310 ( .A(\CARRYB[29][16] ), .B(\SUMB[29][17] ), .Z(\A1[44] ) );
  EO U311 ( .A(\CARRYB[29][22] ), .B(\SUMB[29][23] ), .Z(\A1[50] ) );
  EO U312 ( .A(\CARRYB[29][23] ), .B(\SUMB[29][24] ), .Z(\A1[51] ) );
  EO U313 ( .A(\CARRYB[29][7] ), .B(\SUMB[29][8] ), .Z(\A1[35] ) );
  EO U314 ( .A(\CARRYB[29][25] ), .B(\SUMB[29][26] ), .Z(\A1[53] ) );
  EO U315 ( .A(\CARRYB[29][6] ), .B(\SUMB[29][7] ), .Z(\A1[34] ) );
  EO U316 ( .A(\CARRYB[29][21] ), .B(\SUMB[29][22] ), .Z(\A1[49] ) );
  EO U317 ( .A(\CARRYB[29][27] ), .B(\SUMB[29][28] ), .Z(\A1[55] ) );
  EO U318 ( .A(\CARRYB[29][26] ), .B(\SUMB[29][27] ), .Z(\A1[54] ) );
  EO U319 ( .A(\CARRYB[29][2] ), .B(\SUMB[29][3] ), .Z(\A1[30] ) );
  EO U320 ( .A(\CARRYB[29][37] ), .B(\SUMB[29][38] ), .Z(\A1[65] ) );
  EO U321 ( .A(\CARRYB[29][31] ), .B(\SUMB[29][32] ), .Z(\A1[59] ) );
  EO U322 ( .A(\CARRYB[29][34] ), .B(\SUMB[29][35] ), .Z(\A1[62] ) );
  EO U323 ( .A(\CARRYB[29][33] ), .B(\SUMB[29][34] ), .Z(\A1[61] ) );
  EO U324 ( .A(\CARRYB[29][35] ), .B(\SUMB[29][36] ), .Z(\A1[63] ) );
  EO U325 ( .A(\CARRYB[29][8] ), .B(\SUMB[29][9] ), .Z(\A1[36] ) );
  EO U326 ( .A(\CARRYB[29][4] ), .B(\SUMB[29][5] ), .Z(\A1[32] ) );
  EO U327 ( .A(\CARRYB[29][24] ), .B(\SUMB[29][25] ), .Z(\A1[52] ) );
  EO U328 ( .A(\CARRYB[29][12] ), .B(\SUMB[29][13] ), .Z(\A1[40] ) );
  EO U329 ( .A(\CARRYB[29][29] ), .B(\SUMB[29][30] ), .Z(\A1[57] ) );
  EO U330 ( .A(\CARRYB[29][30] ), .B(\SUMB[29][31] ), .Z(\A1[58] ) );
  EO U331 ( .A(\CARRYB[29][20] ), .B(\SUMB[29][21] ), .Z(\A1[48] ) );
  EO U332 ( .A(\CARRYB[29][3] ), .B(\SUMB[29][4] ), .Z(\A1[31] ) );
  EO U333 ( .A(\CARRYB[29][28] ), .B(\SUMB[29][29] ), .Z(\A1[56] ) );
  EO U334 ( .A(\CARRYB[29][36] ), .B(\SUMB[29][37] ), .Z(\A1[64] ) );
  EO U335 ( .A(\CARRYB[29][32] ), .B(\SUMB[29][33] ), .Z(\A1[60] ) );
  EO U336 ( .A(\CARRYB[29][1] ), .B(\SUMB[29][2] ), .Z(\A1[29] ) );
  EO U337 ( .A(\ab[0][2] ), .B(n3), .Z(\SUMB[1][1] ) );
  IVP U338 ( .A(A[16]), .Z(n563) );
  IVP U339 ( .A(A[17]), .Z(n562) );
  IVP U340 ( .A(A[18]), .Z(n561) );
  IVP U341 ( .A(A[19]), .Z(n560) );
  IVP U342 ( .A(A[20]), .Z(n559) );
  IVP U343 ( .A(A[21]), .Z(n558) );
  IVP U344 ( .A(A[23]), .Z(n556) );
  IVP U345 ( .A(A[24]), .Z(n555) );
  IVP U346 ( .A(A[25]), .Z(n554) );
  IVP U347 ( .A(A[26]), .Z(n553) );
  IVP U348 ( .A(A[27]), .Z(n552) );
  IVP U349 ( .A(A[28]), .Z(n551) );
  IVP U350 ( .A(A[29]), .Z(n550) );
  EO U351 ( .A(\CARRYB[29][0] ), .B(\SUMB[29][1] ), .Z(\A1[28] ) );
  EO U352 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Z(\SUMB[1][20] ) );
  EO U353 ( .A(\CARRYB[29][46] ), .B(\SUMB[29][47] ), .Z(\A1[74] ) );
  EO U354 ( .A(\CARRYB[29][50] ), .B(\SUMB[29][51] ), .Z(\A1[78] ) );
  EO U355 ( .A(\CARRYB[29][49] ), .B(\SUMB[29][50] ), .Z(\A1[77] ) );
  EO U356 ( .A(\CARRYB[29][45] ), .B(\SUMB[29][46] ), .Z(\A1[73] ) );
  EO U357 ( .A(\CARRYB[29][47] ), .B(\SUMB[29][48] ), .Z(\A1[75] ) );
  EO U358 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U359 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U360 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U361 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U362 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U363 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U364 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Z(\SUMB[1][16] ) );
  EO U365 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Z(\SUMB[1][17] ) );
  EO U366 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Z(\SUMB[1][18] ) );
  EO U367 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Z(\SUMB[1][19] ) );
  EO U368 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Z(\SUMB[1][21] ) );
  EO U369 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U370 ( .A(\CARRYB[29][39] ), .B(\SUMB[29][40] ), .Z(\A1[67] ) );
  EO U371 ( .A(\CARRYB[29][41] ), .B(\SUMB[29][42] ), .Z(\A1[69] ) );
  EO U372 ( .A(\CARRYB[29][42] ), .B(\SUMB[29][43] ), .Z(\A1[70] ) );
  EO U373 ( .A(\CARRYB[29][62] ), .B(\SUMB[29][63] ), .Z(\A1[90] ) );
  EO U374 ( .A(\CARRYB[29][61] ), .B(\SUMB[29][62] ), .Z(\A1[89] ) );
  EO U375 ( .A(\CARRYB[29][40] ), .B(\SUMB[29][41] ), .Z(\A1[68] ) );
  EO U376 ( .A(\CARRYB[29][51] ), .B(\SUMB[29][52] ), .Z(\A1[79] ) );
  EO U377 ( .A(\CARRYB[29][38] ), .B(\SUMB[29][39] ), .Z(\A1[66] ) );
  EO U378 ( .A(\CARRYB[29][43] ), .B(\SUMB[29][44] ), .Z(\A1[71] ) );
  EO U379 ( .A(\CARRYB[29][44] ), .B(\SUMB[29][45] ), .Z(\A1[72] ) );
  EO U380 ( .A(\CARRYB[29][48] ), .B(\SUMB[29][49] ), .Z(\A1[76] ) );
  EO U381 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Z(\SUMB[1][22] ) );
  EO U382 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Z(\SUMB[1][23] ) );
  EO U383 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Z(\SUMB[1][24] ) );
  EO U384 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Z(\SUMB[1][25] ) );
  EO U385 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Z(\SUMB[1][26] ) );
  EO U386 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Z(\SUMB[1][27] ) );
  EO U387 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Z(\SUMB[1][28] ) );
  EO U388 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Z(\SUMB[1][29] ) );
  EO U389 ( .A(\ab[0][33] ), .B(\ab[1][32] ), .Z(\SUMB[1][32] ) );
  EO U390 ( .A(\ab[0][34] ), .B(\ab[1][33] ), .Z(\SUMB[1][33] ) );
  EO U391 ( .A(\ab[0][35] ), .B(\ab[1][34] ), .Z(\SUMB[1][34] ) );
  EO U392 ( .A(\ab[0][36] ), .B(\ab[1][35] ), .Z(\SUMB[1][35] ) );
  EO U393 ( .A(\ab[0][37] ), .B(\ab[1][36] ), .Z(\SUMB[1][36] ) );
  EO U394 ( .A(\ab[0][38] ), .B(\ab[1][37] ), .Z(\SUMB[1][37] ) );
  EO U395 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U396 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U397 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U398 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U399 ( .A(\ab[0][63] ), .B(\ab[1][62] ), .Z(\SUMB[1][62] ) );
  EO U400 ( .A(\ab[0][64] ), .B(\ab[1][63] ), .Z(\SUMB[1][63] ) );
  EO U401 ( .A(\ab[0][65] ), .B(\ab[1][64] ), .Z(\SUMB[1][64] ) );
  EO U402 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U403 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U404 ( .A(\CARRYB[29][59] ), .B(\SUMB[29][60] ), .Z(\A1[87] ) );
  EO U405 ( .A(\CARRYB[29][66] ), .B(\SUMB[29][67] ), .Z(\A1[94] ) );
  EO U406 ( .A(\CARRYB[29][67] ), .B(\SUMB[29][68] ), .Z(\A1[95] ) );
  EO U407 ( .A(\CARRYB[29][65] ), .B(\SUMB[29][66] ), .Z(\A1[93] ) );
  EO U408 ( .A(\CARRYB[29][64] ), .B(\SUMB[29][65] ), .Z(\A1[92] ) );
  EO U409 ( .A(\CARRYB[29][63] ), .B(\SUMB[29][64] ), .Z(\A1[91] ) );
  EO U410 ( .A(\CARRYB[29][60] ), .B(\SUMB[29][61] ), .Z(\A1[88] ) );
  EO U411 ( .A(\CARRYB[29][53] ), .B(\SUMB[29][54] ), .Z(\A1[81] ) );
  EO U412 ( .A(\CARRYB[29][55] ), .B(\SUMB[29][56] ), .Z(\A1[83] ) );
  EO U413 ( .A(\CARRYB[29][58] ), .B(\SUMB[29][59] ), .Z(\A1[86] ) );
  EO U414 ( .A(\CARRYB[29][54] ), .B(\SUMB[29][55] ), .Z(\A1[82] ) );
  EO U415 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Z(\SUMB[1][30] ) );
  EO U416 ( .A(\ab[0][32] ), .B(\ab[1][31] ), .Z(\SUMB[1][31] ) );
  EO U417 ( .A(\ab[0][62] ), .B(\ab[1][61] ), .Z(\SUMB[1][61] ) );
  EO U418 ( .A(\ab[0][66] ), .B(\ab[1][65] ), .Z(\SUMB[1][65] ) );
  EO U419 ( .A(\ab[0][67] ), .B(\ab[1][66] ), .Z(\SUMB[1][66] ) );
  EO U420 ( .A(\ab[0][68] ), .B(\ab[1][67] ), .Z(\SUMB[1][67] ) );
  EO U421 ( .A(\ab[0][69] ), .B(\ab[1][68] ), .Z(\SUMB[1][68] ) );
  EO U422 ( .A(\ab[0][70] ), .B(\ab[1][69] ), .Z(\SUMB[1][69] ) );
  EO U423 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U424 ( .A(\CARRYB[29][71] ), .B(\SUMB[29][72] ), .Z(\A1[99] ) );
  EO U425 ( .A(\CARRYB[29][56] ), .B(\SUMB[29][57] ), .Z(\A1[84] ) );
  EO U426 ( .A(\CARRYB[29][69] ), .B(\SUMB[29][70] ), .Z(\A1[97] ) );
  EO U427 ( .A(\CARRYB[29][70] ), .B(\SUMB[29][71] ), .Z(\A1[98] ) );
  EO U428 ( .A(\CARRYB[29][75] ), .B(\SUMB[29][76] ), .Z(\A1[103] ) );
  EO U429 ( .A(\CARRYB[29][77] ), .B(\SUMB[29][78] ), .Z(\A1[105] ) );
  EO U430 ( .A(\CARRYB[29][78] ), .B(\SUMB[29][79] ), .Z(\A1[106] ) );
  EO U431 ( .A(\CARRYB[29][73] ), .B(\SUMB[29][74] ), .Z(\A1[101] ) );
  EO U432 ( .A(\CARRYB[29][74] ), .B(\SUMB[29][75] ), .Z(\A1[102] ) );
  EO U433 ( .A(\CARRYB[29][52] ), .B(\SUMB[29][53] ), .Z(\A1[80] ) );
  EO U434 ( .A(\CARRYB[29][68] ), .B(\SUMB[29][69] ), .Z(\A1[96] ) );
  EO U435 ( .A(\CARRYB[29][72] ), .B(\SUMB[29][73] ), .Z(\A1[100] ) );
  EO U436 ( .A(\CARRYB[29][57] ), .B(\SUMB[29][58] ), .Z(\A1[85] ) );
  EO U437 ( .A(\ab[0][71] ), .B(\ab[1][70] ), .Z(\SUMB[1][70] ) );
  EO U438 ( .A(\ab[0][72] ), .B(\ab[1][71] ), .Z(\SUMB[1][71] ) );
  EO U439 ( .A(\ab[0][73] ), .B(\ab[1][72] ), .Z(\SUMB[1][72] ) );
  EO U440 ( .A(\ab[0][74] ), .B(\ab[1][73] ), .Z(\SUMB[1][73] ) );
  EO U441 ( .A(\ab[0][75] ), .B(\ab[1][74] ), .Z(\SUMB[1][74] ) );
  EO U442 ( .A(\ab[0][76] ), .B(\ab[1][75] ), .Z(\SUMB[1][75] ) );
  EO U443 ( .A(\ab[0][77] ), .B(\ab[1][76] ), .Z(\SUMB[1][76] ) );
  EO U444 ( .A(\ab[0][78] ), .B(\ab[1][77] ), .Z(\SUMB[1][77] ) );
  EO U445 ( .A(\ab[0][79] ), .B(\ab[1][78] ), .Z(\SUMB[1][78] ) );
  EO U446 ( .A(\ab[0][80] ), .B(\ab[1][79] ), .Z(\SUMB[1][79] ) );
  EO U447 ( .A(\ab[0][81] ), .B(\ab[1][80] ), .Z(\SUMB[1][80] ) );
  EO U448 ( .A(\CARRYB[29][83] ), .B(\SUMB[29][84] ), .Z(\A1[111] ) );
  EO U449 ( .A(\CARRYB[29][76] ), .B(\SUMB[29][77] ), .Z(\A1[104] ) );
  EO U450 ( .A(\CARRYB[29][82] ), .B(\SUMB[29][83] ), .Z(\A1[110] ) );
  EO U451 ( .A(\ab[0][82] ), .B(\ab[1][81] ), .Z(\SUMB[1][81] ) );
  EO U452 ( .A(\ab[0][84] ), .B(\ab[1][83] ), .Z(\SUMB[1][83] ) );
  EO U453 ( .A(\ab[0][85] ), .B(\ab[1][84] ), .Z(\SUMB[1][84] ) );
  EO U454 ( .A(\ab[0][86] ), .B(\ab[1][85] ), .Z(\SUMB[1][85] ) );
  EO U455 ( .A(\CARRYB[29][81] ), .B(\SUMB[29][82] ), .Z(\A1[109] ) );
  EO U456 ( .A(\CARRYB[29][79] ), .B(\SUMB[29][80] ), .Z(\A1[107] ) );
  EO U457 ( .A(\CARRYB[29][80] ), .B(\SUMB[29][81] ), .Z(\A1[108] ) );
  EO U458 ( .A(\ab[0][83] ), .B(\ab[1][82] ), .Z(\SUMB[1][82] ) );
  EO U459 ( .A(\ab[0][87] ), .B(\ab[1][86] ), .Z(\SUMB[1][86] ) );
  EO U460 ( .A(\ab[0][88] ), .B(\ab[1][87] ), .Z(\SUMB[1][87] ) );
  EO U461 ( .A(\CARRYB[29][84] ), .B(\SUMB[29][85] ), .Z(\A1[112] ) );
  EO U462 ( .A(\ab[0][89] ), .B(\ab[1][88] ), .Z(\SUMB[1][88] ) );
  EO U463 ( .A(\CARRYB[29][85] ), .B(\SUMB[29][86] ), .Z(\A1[113] ) );
  EO U464 ( .A(\ab[0][90] ), .B(\ab[1][89] ), .Z(\SUMB[1][89] ) );
  EO U465 ( .A(\CARRYB[29][86] ), .B(\SUMB[29][87] ), .Z(\A1[114] ) );
  EO U466 ( .A(\CARRYB[29][87] ), .B(\SUMB[29][88] ), .Z(\A1[115] ) );
  EO U467 ( .A(\ab[0][91] ), .B(\ab[1][90] ), .Z(\SUMB[1][90] ) );
  EO U468 ( .A(\ab[0][92] ), .B(\ab[1][91] ), .Z(\SUMB[1][91] ) );
  EO U469 ( .A(\CARRYB[29][88] ), .B(\SUMB[29][89] ), .Z(\A1[116] ) );
  EO U470 ( .A(\ab[0][93] ), .B(\ab[1][92] ), .Z(\SUMB[1][92] ) );
  EO U471 ( .A(\ab[0][94] ), .B(\ab[1][93] ), .Z(\SUMB[1][93] ) );
  EO U472 ( .A(\ab[0][95] ), .B(\ab[1][94] ), .Z(\SUMB[1][94] ) );
  EO U473 ( .A(\CARRYB[29][89] ), .B(\SUMB[29][90] ), .Z(\A1[117] ) );
  EO U474 ( .A(\CARRYB[29][90] ), .B(\SUMB[29][91] ), .Z(\A1[118] ) );
  EO U475 ( .A(\CARRYB[29][91] ), .B(\SUMB[29][92] ), .Z(\A1[119] ) );
  EO U476 ( .A(\CARRYB[29][92] ), .B(\SUMB[29][93] ), .Z(\A1[120] ) );
  EO U477 ( .A(\CARRYB[29][93] ), .B(\SUMB[29][94] ), .Z(\A1[121] ) );
  EO U478 ( .A(\CARRYB[29][94] ), .B(\ab[29][95] ), .Z(\A1[122] ) );
  EO U479 ( .A(\ab[0][39] ), .B(\ab[1][38] ), .Z(\SUMB[1][38] ) );
  EO U480 ( .A(\ab[0][40] ), .B(\ab[1][39] ), .Z(\SUMB[1][39] ) );
  EO U481 ( .A(\ab[0][57] ), .B(\ab[1][56] ), .Z(\SUMB[1][56] ) );
  IVP U482 ( .A(n526), .Z(n488) );
  IVP U483 ( .A(n532), .Z(n490) );
  IVP U484 ( .A(n527), .Z(n489) );
  IVP U485 ( .A(n525), .Z(n487) );
  IVP U486 ( .A(n524), .Z(n486) );
  IVP U487 ( .A(n523), .Z(n485) );
  IVP U488 ( .A(n522), .Z(n484) );
  IVP U489 ( .A(n521), .Z(n483) );
  IVP U490 ( .A(n520), .Z(n482) );
  IVP U491 ( .A(n519), .Z(n481) );
  IVP U492 ( .A(n518), .Z(n480) );
  IVP U493 ( .A(n517), .Z(n479) );
  IVP U494 ( .A(n516), .Z(n478) );
  IVP U495 ( .A(n515), .Z(n477) );
  IVP U496 ( .A(n514), .Z(n476) );
  IVP U497 ( .A(n513), .Z(n475) );
  IVP U498 ( .A(n512), .Z(n474) );
  IVP U499 ( .A(n510), .Z(n472) );
  IVP U500 ( .A(n509), .Z(n471) );
  IVP U501 ( .A(n508), .Z(n470) );
  IVP U502 ( .A(n511), .Z(n473) );
  IVP U503 ( .A(n507), .Z(n469) );
  IVP U504 ( .A(n506), .Z(n468) );
  IVP U505 ( .A(n504), .Z(n466) );
  IVP U506 ( .A(n503), .Z(n465) );
  IVP U507 ( .A(n502), .Z(n464) );
  IVP U508 ( .A(n505), .Z(n467) );
  IVP U509 ( .A(n501), .Z(n463) );
  IVP U510 ( .A(n500), .Z(n462) );
  IVP U511 ( .A(n499), .Z(n461) );
  IVP U512 ( .A(n498), .Z(n460) );
  IVP U513 ( .A(n338), .Z(n336) );
  IVP U514 ( .A(n342), .Z(n340) );
  IVP U515 ( .A(n346), .Z(n344) );
  IVP U516 ( .A(n350), .Z(n348) );
  IVP U517 ( .A(n354), .Z(n352) );
  IVP U518 ( .A(n358), .Z(n356) );
  IVP U519 ( .A(n362), .Z(n360) );
  IVP U520 ( .A(n366), .Z(n364) );
  IVP U521 ( .A(n370), .Z(n368) );
  IVP U522 ( .A(n374), .Z(n372) );
  IVP U523 ( .A(n378), .Z(n376) );
  IVP U524 ( .A(n382), .Z(n380) );
  IVP U525 ( .A(n497), .Z(n459) );
  IVP U526 ( .A(n386), .Z(n384) );
  IVP U527 ( .A(n390), .Z(n388) );
  IVP U528 ( .A(n394), .Z(n392) );
  IVP U529 ( .A(n398), .Z(n396) );
  IVP U530 ( .A(n402), .Z(n400) );
  IVP U531 ( .A(n406), .Z(n404) );
  IVP U532 ( .A(n438), .Z(n436) );
  IVP U533 ( .A(n450), .Z(n448) );
  IVP U534 ( .A(n454), .Z(n452) );
  IVP U535 ( .A(n326), .Z(n324) );
  IVP U536 ( .A(n330), .Z(n328) );
  IVP U537 ( .A(n334), .Z(n332) );
  IVP U538 ( .A(n322), .Z(n320) );
  IVP U539 ( .A(n310), .Z(n308) );
  IVP U540 ( .A(n314), .Z(n312) );
  IVP U541 ( .A(n496), .Z(n458) );
  IVP U542 ( .A(n410), .Z(n408) );
  IVP U543 ( .A(n414), .Z(n412) );
  IVP U544 ( .A(n418), .Z(n416) );
  IVP U545 ( .A(n422), .Z(n420) );
  IVP U546 ( .A(n426), .Z(n424) );
  IVP U547 ( .A(n430), .Z(n428) );
  IVP U548 ( .A(n434), .Z(n432) );
  IVP U549 ( .A(n442), .Z(n440) );
  IVP U550 ( .A(n446), .Z(n444) );
  IVP U551 ( .A(n318), .Z(n316) );
  IVP U552 ( .A(n306), .Z(n304) );
  IVP U553 ( .A(n495), .Z(n457) );
  IVP U554 ( .A(n302), .Z(n300) );
  IVP U555 ( .A(n494), .Z(n456) );
  IVP U556 ( .A(n493), .Z(n455) );
  IVP U557 ( .A(n492), .Z(n491) );
  IVP U558 ( .A(n338), .Z(n335) );
  IVP U559 ( .A(n342), .Z(n339) );
  IVP U560 ( .A(n346), .Z(n343) );
  IVP U561 ( .A(n350), .Z(n347) );
  IVP U562 ( .A(n354), .Z(n351) );
  IVP U563 ( .A(n358), .Z(n355) );
  IVP U564 ( .A(n362), .Z(n359) );
  IVP U565 ( .A(n366), .Z(n363) );
  IVP U566 ( .A(n370), .Z(n367) );
  IVP U567 ( .A(n374), .Z(n371) );
  IVP U568 ( .A(n378), .Z(n375) );
  IVP U569 ( .A(n382), .Z(n379) );
  IVP U570 ( .A(n386), .Z(n383) );
  IVP U571 ( .A(n390), .Z(n387) );
  IVP U572 ( .A(n394), .Z(n391) );
  IVP U573 ( .A(n398), .Z(n395) );
  IVP U574 ( .A(n402), .Z(n399) );
  IVP U575 ( .A(n406), .Z(n403) );
  IVP U576 ( .A(n438), .Z(n435) );
  IVP U577 ( .A(n326), .Z(n323) );
  IVP U578 ( .A(n330), .Z(n327) );
  IVP U579 ( .A(n334), .Z(n331) );
  IVP U580 ( .A(n322), .Z(n319) );
  IVP U581 ( .A(n454), .Z(n451) );
  IVP U582 ( .A(n310), .Z(n307) );
  IVP U583 ( .A(n314), .Z(n311) );
  IVP U584 ( .A(n450), .Z(n447) );
  IVP U585 ( .A(n410), .Z(n407) );
  IVP U586 ( .A(n414), .Z(n411) );
  IVP U587 ( .A(n418), .Z(n415) );
  IVP U588 ( .A(n422), .Z(n419) );
  IVP U589 ( .A(n426), .Z(n423) );
  IVP U590 ( .A(n430), .Z(n427) );
  IVP U591 ( .A(n434), .Z(n431) );
  IVP U592 ( .A(n446), .Z(n443) );
  IVP U593 ( .A(n318), .Z(n315) );
  IVP U594 ( .A(n442), .Z(n439) );
  IVP U595 ( .A(n306), .Z(n303) );
  IVP U596 ( .A(n302), .Z(n299) );
  EO U597 ( .A(\ab[0][47] ), .B(\ab[1][46] ), .Z(\SUMB[1][46] ) );
  EO U598 ( .A(\ab[0][48] ), .B(\ab[1][47] ), .Z(\SUMB[1][47] ) );
  EO U599 ( .A(\ab[0][49] ), .B(\ab[1][48] ), .Z(\SUMB[1][48] ) );
  EO U600 ( .A(\ab[0][50] ), .B(\ab[1][49] ), .Z(\SUMB[1][49] ) );
  EO U601 ( .A(\ab[0][51] ), .B(\ab[1][50] ), .Z(\SUMB[1][50] ) );
  EO U602 ( .A(\ab[0][52] ), .B(\ab[1][51] ), .Z(\SUMB[1][51] ) );
  EO U603 ( .A(\ab[0][53] ), .B(\ab[1][52] ), .Z(\SUMB[1][52] ) );
  EO U604 ( .A(\ab[0][41] ), .B(\ab[1][40] ), .Z(\SUMB[1][40] ) );
  EO U605 ( .A(\ab[0][42] ), .B(\ab[1][41] ), .Z(\SUMB[1][41] ) );
  EO U606 ( .A(\ab[0][43] ), .B(\ab[1][42] ), .Z(\SUMB[1][42] ) );
  EO U607 ( .A(\ab[0][44] ), .B(\ab[1][43] ), .Z(\SUMB[1][43] ) );
  EO U608 ( .A(\ab[0][45] ), .B(\ab[1][44] ), .Z(\SUMB[1][44] ) );
  EO U609 ( .A(\ab[0][46] ), .B(\ab[1][45] ), .Z(\SUMB[1][45] ) );
  EO U610 ( .A(\ab[0][54] ), .B(\ab[1][53] ), .Z(\SUMB[1][53] ) );
  EO U611 ( .A(\ab[0][55] ), .B(\ab[1][54] ), .Z(\SUMB[1][54] ) );
  EO U612 ( .A(\ab[0][56] ), .B(\ab[1][55] ), .Z(\SUMB[1][55] ) );
  EO U613 ( .A(\ab[0][58] ), .B(\ab[1][57] ), .Z(\SUMB[1][57] ) );
  EO U614 ( .A(\ab[0][60] ), .B(\ab[1][59] ), .Z(\SUMB[1][59] ) );
  EO U615 ( .A(\ab[0][61] ), .B(\ab[1][60] ), .Z(\SUMB[1][60] ) );
  EO U616 ( .A(\ab[0][59] ), .B(\ab[1][58] ), .Z(\SUMB[1][58] ) );
  IVP U617 ( .A(B[61]), .Z(n526) );
  IVP U618 ( .A(B[55]), .Z(n532) );
  IVP U619 ( .A(B[60]), .Z(n527) );
  IVP U620 ( .A(B[62]), .Z(n525) );
  IVP U621 ( .A(B[63]), .Z(n524) );
  IVP U622 ( .A(B[64]), .Z(n523) );
  IVP U623 ( .A(B[65]), .Z(n522) );
  IVP U624 ( .A(B[66]), .Z(n521) );
  IVP U625 ( .A(B[67]), .Z(n520) );
  IVP U626 ( .A(B[68]), .Z(n519) );
  IVP U627 ( .A(B[69]), .Z(n518) );
  IVP U628 ( .A(B[70]), .Z(n517) );
  IVP U629 ( .A(B[71]), .Z(n516) );
  IVP U630 ( .A(B[72]), .Z(n515) );
  IVP U631 ( .A(B[73]), .Z(n514) );
  IVP U632 ( .A(B[74]), .Z(n513) );
  IVP U633 ( .A(B[75]), .Z(n512) );
  IVP U634 ( .A(B[77]), .Z(n510) );
  IVP U635 ( .A(B[78]), .Z(n509) );
  IVP U636 ( .A(B[79]), .Z(n508) );
  IVP U637 ( .A(B[76]), .Z(n511) );
  IVP U638 ( .A(B[80]), .Z(n507) );
  IVP U639 ( .A(B[81]), .Z(n506) );
  IVP U640 ( .A(B[83]), .Z(n504) );
  IVP U641 ( .A(B[84]), .Z(n503) );
  IVP U642 ( .A(B[85]), .Z(n502) );
  IVP U643 ( .A(B[82]), .Z(n505) );
  IVP U644 ( .A(B[86]), .Z(n501) );
  IVP U645 ( .A(B[87]), .Z(n500) );
  IVP U646 ( .A(B[88]), .Z(n499) );
  IVP U647 ( .A(B[89]), .Z(n498) );
  IVP U648 ( .A(B[90]), .Z(n497) );
  IVP U649 ( .A(B[91]), .Z(n496) );
  IVP U650 ( .A(B[92]), .Z(n495) );
  IVP U651 ( .A(B[93]), .Z(n494) );
  IVP U652 ( .A(B[94]), .Z(n493) );
  IVP U653 ( .A(B[45]), .Z(n542) );
  IVP U654 ( .A(B[46]), .Z(n541) );
  IVP U655 ( .A(B[47]), .Z(n540) );
  IVP U656 ( .A(B[48]), .Z(n539) );
  IVP U657 ( .A(B[49]), .Z(n538) );
  IVP U658 ( .A(B[50]), .Z(n537) );
  IVP U659 ( .A(B[51]), .Z(n536) );
  IVP U660 ( .A(B[39]), .Z(n548) );
  IVP U661 ( .A(B[58]), .Z(n529) );
  IVP U662 ( .A(B[40]), .Z(n547) );
  IVP U663 ( .A(B[41]), .Z(n546) );
  IVP U664 ( .A(B[42]), .Z(n545) );
  IVP U665 ( .A(B[43]), .Z(n544) );
  IVP U666 ( .A(B[44]), .Z(n543) );
  IVP U667 ( .A(B[52]), .Z(n535) );
  IVP U668 ( .A(B[53]), .Z(n534) );
  IVP U669 ( .A(B[57]), .Z(n530) );
  IVP U670 ( .A(B[59]), .Z(n528) );
  IVP U671 ( .A(B[54]), .Z(n533) );
  IVP U672 ( .A(B[56]), .Z(n531) );
  IVP U673 ( .A(B[95]), .Z(n492) );
  AN2P U674 ( .A(\CARRYB[29][0] ), .B(\SUMB[29][1] ), .Z(\A2[29] ) );
  AN2P U675 ( .A(\CARRYB[29][1] ), .B(\SUMB[29][2] ), .Z(\A2[30] ) );
  AN2P U676 ( .A(\CARRYB[29][2] ), .B(\SUMB[29][3] ), .Z(\A2[31] ) );
  AN2P U677 ( .A(\CARRYB[29][3] ), .B(\SUMB[29][4] ), .Z(\A2[32] ) );
  AN2P U678 ( .A(\CARRYB[29][4] ), .B(\SUMB[29][5] ), .Z(\A2[33] ) );
  AN2P U679 ( .A(\CARRYB[29][5] ), .B(\SUMB[29][6] ), .Z(\A2[34] ) );
  AN2P U680 ( .A(\CARRYB[29][6] ), .B(\SUMB[29][7] ), .Z(\A2[35] ) );
  AN2P U681 ( .A(\CARRYB[29][7] ), .B(\SUMB[29][8] ), .Z(\A2[36] ) );
  AN2P U682 ( .A(\CARRYB[29][8] ), .B(\SUMB[29][9] ), .Z(\A2[37] ) );
  AN2P U683 ( .A(\CARRYB[29][9] ), .B(\SUMB[29][10] ), .Z(\A2[38] ) );
  AN2P U684 ( .A(\CARRYB[29][10] ), .B(\SUMB[29][11] ), .Z(\A2[39] ) );
  AN2P U685 ( .A(\CARRYB[29][11] ), .B(\SUMB[29][12] ), .Z(\A2[40] ) );
  AN2P U686 ( .A(\CARRYB[29][12] ), .B(\SUMB[29][13] ), .Z(\A2[41] ) );
  AN2P U687 ( .A(\CARRYB[29][13] ), .B(\SUMB[29][14] ), .Z(\A2[42] ) );
  AN2P U688 ( .A(\CARRYB[29][14] ), .B(\SUMB[29][15] ), .Z(\A2[43] ) );
  AN2P U689 ( .A(\CARRYB[29][15] ), .B(\SUMB[29][16] ), .Z(\A2[44] ) );
  AN2P U690 ( .A(\CARRYB[29][16] ), .B(\SUMB[29][17] ), .Z(\A2[45] ) );
  AN2P U691 ( .A(\CARRYB[29][17] ), .B(\SUMB[29][18] ), .Z(\A2[46] ) );
  AN2P U692 ( .A(\CARRYB[29][18] ), .B(\SUMB[29][19] ), .Z(\A2[47] ) );
  AN2P U693 ( .A(\CARRYB[29][19] ), .B(\SUMB[29][20] ), .Z(\A2[48] ) );
  AN2P U694 ( .A(\CARRYB[29][20] ), .B(\SUMB[29][21] ), .Z(\A2[49] ) );
  AN2P U695 ( .A(\CARRYB[29][21] ), .B(\SUMB[29][22] ), .Z(\A2[50] ) );
  AN2P U696 ( .A(\CARRYB[29][22] ), .B(\SUMB[29][23] ), .Z(\A2[51] ) );
  AN2P U697 ( .A(\CARRYB[29][23] ), .B(\SUMB[29][24] ), .Z(\A2[52] ) );
  AN2P U698 ( .A(\CARRYB[29][24] ), .B(\SUMB[29][25] ), .Z(\A2[53] ) );
  AN2P U699 ( .A(\CARRYB[29][25] ), .B(\SUMB[29][26] ), .Z(\A2[54] ) );
  AN2P U700 ( .A(\CARRYB[29][26] ), .B(\SUMB[29][27] ), .Z(\A2[55] ) );
  AN2P U701 ( .A(\CARRYB[29][27] ), .B(\SUMB[29][28] ), .Z(\A2[56] ) );
  AN2P U702 ( .A(\CARRYB[29][28] ), .B(\SUMB[29][29] ), .Z(\A2[57] ) );
  AN2P U703 ( .A(\CARRYB[29][29] ), .B(\SUMB[29][30] ), .Z(\A2[58] ) );
  AN2P U704 ( .A(\CARRYB[29][30] ), .B(\SUMB[29][31] ), .Z(\A2[59] ) );
  AN2P U705 ( .A(\CARRYB[29][31] ), .B(\SUMB[29][32] ), .Z(\A2[60] ) );
  AN2P U706 ( .A(\CARRYB[29][32] ), .B(\SUMB[29][33] ), .Z(\A2[61] ) );
  AN2P U707 ( .A(\CARRYB[29][33] ), .B(\SUMB[29][34] ), .Z(\A2[62] ) );
  AN2P U708 ( .A(\CARRYB[29][34] ), .B(\SUMB[29][35] ), .Z(\A2[63] ) );
  AN2P U709 ( .A(\CARRYB[29][35] ), .B(\SUMB[29][36] ), .Z(\A2[64] ) );
  AN2P U710 ( .A(\CARRYB[29][36] ), .B(\SUMB[29][37] ), .Z(\A2[65] ) );
  AN2P U711 ( .A(\CARRYB[29][37] ), .B(\SUMB[29][38] ), .Z(\A2[66] ) );
  AN2P U712 ( .A(\CARRYB[29][38] ), .B(\SUMB[29][39] ), .Z(\A2[67] ) );
  AN2P U713 ( .A(\CARRYB[29][39] ), .B(\SUMB[29][40] ), .Z(\A2[68] ) );
  AN2P U714 ( .A(\CARRYB[29][40] ), .B(\SUMB[29][41] ), .Z(\A2[69] ) );
  AN2P U715 ( .A(\CARRYB[29][41] ), .B(\SUMB[29][42] ), .Z(\A2[70] ) );
  AN2P U716 ( .A(\CARRYB[29][42] ), .B(\SUMB[29][43] ), .Z(\A2[71] ) );
  AN2P U717 ( .A(\CARRYB[29][43] ), .B(\SUMB[29][44] ), .Z(\A2[72] ) );
  AN2P U718 ( .A(\CARRYB[29][44] ), .B(\SUMB[29][45] ), .Z(\A2[73] ) );
  AN2P U719 ( .A(\CARRYB[29][45] ), .B(\SUMB[29][46] ), .Z(\A2[74] ) );
  AN2P U720 ( .A(\CARRYB[29][46] ), .B(\SUMB[29][47] ), .Z(\A2[75] ) );
  AN2P U721 ( .A(\CARRYB[29][47] ), .B(\SUMB[29][48] ), .Z(\A2[76] ) );
  AN2P U722 ( .A(\CARRYB[29][48] ), .B(\SUMB[29][49] ), .Z(\A2[77] ) );
  AN2P U723 ( .A(\CARRYB[29][49] ), .B(\SUMB[29][50] ), .Z(\A2[78] ) );
  AN2P U724 ( .A(\CARRYB[29][50] ), .B(\SUMB[29][51] ), .Z(\A2[79] ) );
  AN2P U725 ( .A(\CARRYB[29][51] ), .B(\SUMB[29][52] ), .Z(\A2[80] ) );
  AN2P U726 ( .A(\CARRYB[29][52] ), .B(\SUMB[29][53] ), .Z(\A2[81] ) );
  AN2P U727 ( .A(\CARRYB[29][53] ), .B(\SUMB[29][54] ), .Z(\A2[82] ) );
  AN2P U728 ( .A(\CARRYB[29][54] ), .B(\SUMB[29][55] ), .Z(\A2[83] ) );
  AN2P U729 ( .A(\CARRYB[29][55] ), .B(\SUMB[29][56] ), .Z(\A2[84] ) );
  AN2P U730 ( .A(\CARRYB[29][56] ), .B(\SUMB[29][57] ), .Z(\A2[85] ) );
  AN2P U731 ( .A(\CARRYB[29][57] ), .B(\SUMB[29][58] ), .Z(\A2[86] ) );
  AN2P U732 ( .A(\CARRYB[29][58] ), .B(\SUMB[29][59] ), .Z(\A2[87] ) );
  AN2P U733 ( .A(\CARRYB[29][59] ), .B(\SUMB[29][60] ), .Z(\A2[88] ) );
  AN2P U734 ( .A(\CARRYB[29][60] ), .B(\SUMB[29][61] ), .Z(\A2[89] ) );
  AN2P U735 ( .A(\CARRYB[29][61] ), .B(\SUMB[29][62] ), .Z(\A2[90] ) );
  AN2P U736 ( .A(\CARRYB[29][62] ), .B(\SUMB[29][63] ), .Z(\A2[91] ) );
  AN2P U737 ( .A(\CARRYB[29][63] ), .B(\SUMB[29][64] ), .Z(\A2[92] ) );
  AN2P U738 ( .A(\CARRYB[29][64] ), .B(\SUMB[29][65] ), .Z(\A2[93] ) );
  AN2P U739 ( .A(\CARRYB[29][66] ), .B(\SUMB[29][67] ), .Z(\A2[95] ) );
  AN2P U740 ( .A(\CARRYB[29][67] ), .B(\SUMB[29][68] ), .Z(\A2[96] ) );
  AN2P U741 ( .A(\CARRYB[29][68] ), .B(\SUMB[29][69] ), .Z(\A2[97] ) );
  AN2P U742 ( .A(\CARRYB[29][69] ), .B(\SUMB[29][70] ), .Z(\A2[98] ) );
  AN2P U743 ( .A(\CARRYB[29][70] ), .B(\SUMB[29][71] ), .Z(\A2[99] ) );
  AN2P U744 ( .A(\CARRYB[29][71] ), .B(\SUMB[29][72] ), .Z(\A2[100] ) );
  AN2P U745 ( .A(\CARRYB[29][72] ), .B(\SUMB[29][73] ), .Z(\A2[101] ) );
  AN2P U746 ( .A(\CARRYB[29][73] ), .B(\SUMB[29][74] ), .Z(\A2[102] ) );
  AN2P U747 ( .A(\CARRYB[29][74] ), .B(\SUMB[29][75] ), .Z(\A2[103] ) );
  AN2P U748 ( .A(\CARRYB[29][75] ), .B(\SUMB[29][76] ), .Z(\A2[104] ) );
  AN2P U749 ( .A(\CARRYB[29][76] ), .B(\SUMB[29][77] ), .Z(\A2[105] ) );
  AN2P U750 ( .A(\CARRYB[29][77] ), .B(\SUMB[29][78] ), .Z(\A2[106] ) );
  AN2P U751 ( .A(\CARRYB[29][78] ), .B(\SUMB[29][79] ), .Z(\A2[107] ) );
  AN2P U752 ( .A(\CARRYB[29][79] ), .B(\SUMB[29][80] ), .Z(\A2[108] ) );
  AN2P U753 ( .A(\CARRYB[29][80] ), .B(\SUMB[29][81] ), .Z(\A2[109] ) );
  AN2P U754 ( .A(\CARRYB[29][81] ), .B(\SUMB[29][82] ), .Z(\A2[110] ) );
  AN2P U755 ( .A(\CARRYB[29][82] ), .B(\SUMB[29][83] ), .Z(\A2[111] ) );
  AN2P U756 ( .A(\CARRYB[29][83] ), .B(\SUMB[29][84] ), .Z(\A2[112] ) );
  AN2P U757 ( .A(\CARRYB[29][84] ), .B(\SUMB[29][85] ), .Z(\A2[113] ) );
  AN2P U758 ( .A(\CARRYB[29][85] ), .B(\SUMB[29][86] ), .Z(\A2[114] ) );
  AN2P U759 ( .A(\CARRYB[29][86] ), .B(\SUMB[29][87] ), .Z(\A2[115] ) );
  AN2P U760 ( .A(\CARRYB[29][87] ), .B(\SUMB[29][88] ), .Z(\A2[116] ) );
  AN2P U761 ( .A(\CARRYB[29][88] ), .B(\SUMB[29][89] ), .Z(\A2[117] ) );
  AN2P U762 ( .A(\CARRYB[29][89] ), .B(\SUMB[29][90] ), .Z(\A2[118] ) );
  AN2P U763 ( .A(\CARRYB[29][90] ), .B(\SUMB[29][91] ), .Z(\A2[119] ) );
  AN2P U764 ( .A(\CARRYB[29][91] ), .B(\SUMB[29][92] ), .Z(\A2[120] ) );
  AN2P U765 ( .A(\CARRYB[29][92] ), .B(\SUMB[29][93] ), .Z(\A2[121] ) );
  AN2P U766 ( .A(\CARRYB[29][93] ), .B(\SUMB[29][94] ), .Z(\A2[122] ) );
  AN2P U767 ( .A(\CARRYB[29][94] ), .B(\ab[29][95] ), .Z(\A2[123] ) );
  AN2P U768 ( .A(n3), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U769 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U770 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U771 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U772 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U773 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U774 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U775 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U776 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U777 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U778 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U779 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U780 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U781 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U782 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U783 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\CARRYB[1][16] ) );
  AN2P U784 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\CARRYB[1][17] ) );
  AN2P U785 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\CARRYB[1][18] ) );
  AN2P U786 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\CARRYB[1][19] ) );
  AN2P U787 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\CARRYB[1][20] ) );
  AN2P U788 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\CARRYB[1][21] ) );
  AN2P U789 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(\CARRYB[1][22] ) );
  AN2P U790 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(\CARRYB[1][23] ) );
  AN2P U791 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(\CARRYB[1][24] ) );
  AN2P U792 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(\CARRYB[1][25] ) );
  AN2P U793 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\CARRYB[1][26] ) );
  AN2P U794 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(\CARRYB[1][27] ) );
  AN2P U795 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(\CARRYB[1][28] ) );
  AN2P U796 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(\CARRYB[1][29] ) );
  AN2P U797 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(\CARRYB[1][30] ) );
  AN2P U798 ( .A(\ab[1][31] ), .B(\ab[0][32] ), .Z(\CARRYB[1][31] ) );
  AN2P U799 ( .A(\ab[1][32] ), .B(\ab[0][33] ), .Z(\CARRYB[1][32] ) );
  AN2P U800 ( .A(\ab[1][33] ), .B(\ab[0][34] ), .Z(\CARRYB[1][33] ) );
  AN2P U801 ( .A(\ab[1][34] ), .B(\ab[0][35] ), .Z(\CARRYB[1][34] ) );
  AN2P U802 ( .A(\ab[1][35] ), .B(\ab[0][36] ), .Z(\CARRYB[1][35] ) );
  AN2P U803 ( .A(\ab[1][36] ), .B(\ab[0][37] ), .Z(\CARRYB[1][36] ) );
  AN2P U804 ( .A(\ab[1][37] ), .B(\ab[0][38] ), .Z(\CARRYB[1][37] ) );
  AN2P U805 ( .A(\ab[1][38] ), .B(\ab[0][39] ), .Z(\CARRYB[1][38] ) );
  AN2P U806 ( .A(\ab[1][39] ), .B(\ab[0][40] ), .Z(\CARRYB[1][39] ) );
  AN2P U807 ( .A(\ab[1][40] ), .B(\ab[0][41] ), .Z(\CARRYB[1][40] ) );
  AN2P U808 ( .A(\ab[1][41] ), .B(\ab[0][42] ), .Z(\CARRYB[1][41] ) );
  AN2P U809 ( .A(\ab[1][42] ), .B(\ab[0][43] ), .Z(\CARRYB[1][42] ) );
  AN2P U810 ( .A(\ab[1][43] ), .B(\ab[0][44] ), .Z(\CARRYB[1][43] ) );
  AN2P U811 ( .A(\ab[1][44] ), .B(\ab[0][45] ), .Z(\CARRYB[1][44] ) );
  AN2P U812 ( .A(\ab[1][45] ), .B(\ab[0][46] ), .Z(\CARRYB[1][45] ) );
  AN2P U813 ( .A(\ab[1][46] ), .B(\ab[0][47] ), .Z(\CARRYB[1][46] ) );
  AN2P U814 ( .A(\ab[1][47] ), .B(\ab[0][48] ), .Z(\CARRYB[1][47] ) );
  AN2P U815 ( .A(\ab[1][48] ), .B(\ab[0][49] ), .Z(\CARRYB[1][48] ) );
  AN2P U816 ( .A(\ab[1][49] ), .B(\ab[0][50] ), .Z(\CARRYB[1][49] ) );
  AN2P U817 ( .A(\ab[1][50] ), .B(\ab[0][51] ), .Z(\CARRYB[1][50] ) );
  AN2P U818 ( .A(\ab[1][51] ), .B(\ab[0][52] ), .Z(\CARRYB[1][51] ) );
  AN2P U819 ( .A(\ab[1][52] ), .B(\ab[0][53] ), .Z(\CARRYB[1][52] ) );
  AN2P U820 ( .A(\ab[1][53] ), .B(\ab[0][54] ), .Z(\CARRYB[1][53] ) );
  AN2P U821 ( .A(\ab[1][54] ), .B(\ab[0][55] ), .Z(\CARRYB[1][54] ) );
  AN2P U822 ( .A(\ab[1][55] ), .B(\ab[0][56] ), .Z(\CARRYB[1][55] ) );
  AN2P U823 ( .A(\ab[1][56] ), .B(\ab[0][57] ), .Z(\CARRYB[1][56] ) );
  AN2P U824 ( .A(\ab[1][57] ), .B(\ab[0][58] ), .Z(\CARRYB[1][57] ) );
  AN2P U825 ( .A(\ab[1][58] ), .B(\ab[0][59] ), .Z(\CARRYB[1][58] ) );
  AN2P U826 ( .A(\ab[1][59] ), .B(\ab[0][60] ), .Z(\CARRYB[1][59] ) );
  AN2P U827 ( .A(\ab[1][60] ), .B(\ab[0][61] ), .Z(\CARRYB[1][60] ) );
  AN2P U828 ( .A(\ab[1][61] ), .B(\ab[0][62] ), .Z(\CARRYB[1][61] ) );
  AN2P U829 ( .A(\ab[1][62] ), .B(\ab[0][63] ), .Z(\CARRYB[1][62] ) );
  AN2P U830 ( .A(\ab[1][63] ), .B(\ab[0][64] ), .Z(\CARRYB[1][63] ) );
  AN2P U831 ( .A(\ab[1][64] ), .B(\ab[0][65] ), .Z(\CARRYB[1][64] ) );
  AN2P U832 ( .A(\ab[1][65] ), .B(\ab[0][66] ), .Z(\CARRYB[1][65] ) );
  AN2P U833 ( .A(\ab[1][66] ), .B(\ab[0][67] ), .Z(\CARRYB[1][66] ) );
  AN2P U834 ( .A(\ab[1][67] ), .B(\ab[0][68] ), .Z(\CARRYB[1][67] ) );
  AN2P U835 ( .A(\ab[1][68] ), .B(\ab[0][69] ), .Z(\CARRYB[1][68] ) );
  AN2P U836 ( .A(\ab[1][69] ), .B(\ab[0][70] ), .Z(\CARRYB[1][69] ) );
  AN2P U837 ( .A(\ab[1][70] ), .B(\ab[0][71] ), .Z(\CARRYB[1][70] ) );
  AN2P U838 ( .A(\ab[1][71] ), .B(\ab[0][72] ), .Z(\CARRYB[1][71] ) );
  AN2P U839 ( .A(\ab[1][72] ), .B(\ab[0][73] ), .Z(\CARRYB[1][72] ) );
  AN2P U840 ( .A(\ab[1][73] ), .B(\ab[0][74] ), .Z(\CARRYB[1][73] ) );
  AN2P U841 ( .A(\ab[1][74] ), .B(\ab[0][75] ), .Z(\CARRYB[1][74] ) );
  AN2P U842 ( .A(\ab[1][75] ), .B(\ab[0][76] ), .Z(\CARRYB[1][75] ) );
  AN2P U843 ( .A(\ab[1][76] ), .B(\ab[0][77] ), .Z(\CARRYB[1][76] ) );
  AN2P U844 ( .A(\ab[1][77] ), .B(\ab[0][78] ), .Z(\CARRYB[1][77] ) );
  AN2P U845 ( .A(\ab[1][78] ), .B(\ab[0][79] ), .Z(\CARRYB[1][78] ) );
  AN2P U846 ( .A(\ab[1][79] ), .B(\ab[0][80] ), .Z(\CARRYB[1][79] ) );
  AN2P U847 ( .A(\ab[1][80] ), .B(\ab[0][81] ), .Z(\CARRYB[1][80] ) );
  AN2P U848 ( .A(\ab[1][81] ), .B(\ab[0][82] ), .Z(\CARRYB[1][81] ) );
  AN2P U849 ( .A(\ab[1][82] ), .B(\ab[0][83] ), .Z(\CARRYB[1][82] ) );
  AN2P U850 ( .A(\ab[1][83] ), .B(\ab[0][84] ), .Z(\CARRYB[1][83] ) );
  AN2P U851 ( .A(\ab[1][84] ), .B(\ab[0][85] ), .Z(\CARRYB[1][84] ) );
  AN2P U852 ( .A(\ab[1][85] ), .B(\ab[0][86] ), .Z(\CARRYB[1][85] ) );
  AN2P U853 ( .A(\ab[1][86] ), .B(\ab[0][87] ), .Z(\CARRYB[1][86] ) );
  AN2P U854 ( .A(\ab[1][87] ), .B(\ab[0][88] ), .Z(\CARRYB[1][87] ) );
  AN2P U855 ( .A(\ab[1][88] ), .B(\ab[0][89] ), .Z(\CARRYB[1][88] ) );
  AN2P U856 ( .A(\ab[1][89] ), .B(\ab[0][90] ), .Z(\CARRYB[1][89] ) );
  AN2P U857 ( .A(\ab[1][90] ), .B(\ab[0][91] ), .Z(\CARRYB[1][90] ) );
  AN2P U858 ( .A(\ab[1][91] ), .B(\ab[0][92] ), .Z(\CARRYB[1][91] ) );
  AN2P U859 ( .A(\ab[1][92] ), .B(\ab[0][93] ), .Z(\CARRYB[1][92] ) );
  AN2P U860 ( .A(\ab[1][93] ), .B(\ab[0][94] ), .Z(\CARRYB[1][93] ) );
  AN2P U861 ( .A(\ab[1][94] ), .B(\ab[0][95] ), .Z(\CARRYB[1][94] ) );
  AN2P U862 ( .A(\CARRYB[29][65] ), .B(\SUMB[29][66] ), .Z(\A2[94] ) );
  IVA U863 ( .A(n302), .Z(n301) );
  IVA U864 ( .A(B[0]), .Z(n302) );
  IVA U865 ( .A(n306), .Z(n305) );
  IVA U866 ( .A(B[1]), .Z(n306) );
  IVA U867 ( .A(n310), .Z(n309) );
  IVA U868 ( .A(B[2]), .Z(n310) );
  IVA U869 ( .A(n314), .Z(n313) );
  IVA U870 ( .A(B[3]), .Z(n314) );
  IVA U871 ( .A(n318), .Z(n317) );
  IVA U872 ( .A(B[4]), .Z(n318) );
  IVA U873 ( .A(n322), .Z(n321) );
  IVA U874 ( .A(B[5]), .Z(n322) );
  IVA U875 ( .A(n326), .Z(n325) );
  IVA U876 ( .A(B[6]), .Z(n326) );
  IVA U877 ( .A(n330), .Z(n329) );
  IVA U878 ( .A(B[7]), .Z(n330) );
  IVA U879 ( .A(n334), .Z(n333) );
  IVA U880 ( .A(B[8]), .Z(n334) );
  IVA U881 ( .A(n338), .Z(n337) );
  IVA U882 ( .A(B[9]), .Z(n338) );
  IVA U883 ( .A(n342), .Z(n341) );
  IVA U884 ( .A(B[10]), .Z(n342) );
  IVA U885 ( .A(n346), .Z(n345) );
  IVA U886 ( .A(B[11]), .Z(n346) );
  IVA U887 ( .A(n350), .Z(n349) );
  IVA U888 ( .A(B[12]), .Z(n350) );
  IVA U889 ( .A(n354), .Z(n353) );
  IVA U890 ( .A(B[13]), .Z(n354) );
  IVA U891 ( .A(n358), .Z(n357) );
  IVA U892 ( .A(B[14]), .Z(n358) );
  IVA U893 ( .A(n362), .Z(n361) );
  IVA U894 ( .A(B[15]), .Z(n362) );
  IVA U895 ( .A(n366), .Z(n365) );
  IVA U896 ( .A(B[16]), .Z(n366) );
  IVA U897 ( .A(n370), .Z(n369) );
  IVA U898 ( .A(B[17]), .Z(n370) );
  IVA U899 ( .A(n374), .Z(n373) );
  IVA U900 ( .A(B[18]), .Z(n374) );
  IVA U901 ( .A(n378), .Z(n377) );
  IVA U902 ( .A(B[19]), .Z(n378) );
  IVA U903 ( .A(n382), .Z(n381) );
  IVA U904 ( .A(B[20]), .Z(n382) );
  IVA U905 ( .A(n386), .Z(n385) );
  IVA U906 ( .A(B[21]), .Z(n386) );
  IVA U907 ( .A(n390), .Z(n389) );
  IVA U908 ( .A(B[22]), .Z(n390) );
  IVA U909 ( .A(n394), .Z(n393) );
  IVA U910 ( .A(B[23]), .Z(n394) );
  IVA U911 ( .A(n398), .Z(n397) );
  IVA U912 ( .A(B[24]), .Z(n398) );
  IVA U913 ( .A(n402), .Z(n401) );
  IVA U914 ( .A(B[25]), .Z(n402) );
  IVA U915 ( .A(n406), .Z(n405) );
  IVA U916 ( .A(B[26]), .Z(n406) );
  IVA U917 ( .A(n410), .Z(n409) );
  IVA U918 ( .A(B[27]), .Z(n410) );
  IVA U919 ( .A(n414), .Z(n413) );
  IVA U920 ( .A(B[28]), .Z(n414) );
  IVA U921 ( .A(n418), .Z(n417) );
  IVA U922 ( .A(B[29]), .Z(n418) );
  IVA U923 ( .A(n422), .Z(n421) );
  IVA U924 ( .A(B[30]), .Z(n422) );
  IVA U925 ( .A(n426), .Z(n425) );
  IVA U926 ( .A(B[31]), .Z(n426) );
  IVA U927 ( .A(n430), .Z(n429) );
  IVA U928 ( .A(B[32]), .Z(n430) );
  IVA U929 ( .A(n434), .Z(n433) );
  IVA U930 ( .A(B[33]), .Z(n434) );
  IVA U931 ( .A(n438), .Z(n437) );
  IVA U932 ( .A(B[34]), .Z(n438) );
  IVA U933 ( .A(n442), .Z(n441) );
  IVA U934 ( .A(B[35]), .Z(n442) );
  IVA U935 ( .A(n446), .Z(n445) );
  IVA U936 ( .A(B[36]), .Z(n446) );
  IVA U937 ( .A(n450), .Z(n449) );
  IVA U938 ( .A(B[37]), .Z(n450) );
  IVA U939 ( .A(n454), .Z(n453) );
  IVA U940 ( .A(B[38]), .Z(n454) );
  AN2P U941 ( .A(n171), .B(n491), .Z(\ab[0][95] ) );
  AN2P U942 ( .A(n180), .B(n455), .Z(\ab[1][94] ) );
  AN2P U943 ( .A(n171), .B(n455), .Z(\ab[0][94] ) );
  AN2P U944 ( .A(n180), .B(n456), .Z(\ab[1][93] ) );
  AN2P U945 ( .A(n171), .B(n456), .Z(\ab[0][93] ) );
  AN2P U946 ( .A(n180), .B(n457), .Z(\ab[1][92] ) );
  AN2P U947 ( .A(n171), .B(n457), .Z(\ab[0][92] ) );
  AN2P U948 ( .A(n180), .B(n458), .Z(\ab[1][91] ) );
  AN2P U949 ( .A(n171), .B(n458), .Z(\ab[0][91] ) );
  AN2P U950 ( .A(n180), .B(n459), .Z(\ab[1][90] ) );
  AN2P U951 ( .A(n171), .B(n459), .Z(\ab[0][90] ) );
  AN2P U952 ( .A(n180), .B(n460), .Z(\ab[1][89] ) );
  AN2P U953 ( .A(n171), .B(n460), .Z(\ab[0][89] ) );
  AN2P U954 ( .A(n180), .B(n461), .Z(\ab[1][88] ) );
  AN2P U955 ( .A(n171), .B(n461), .Z(\ab[0][88] ) );
  AN2P U956 ( .A(n180), .B(n462), .Z(\ab[1][87] ) );
  AN2P U957 ( .A(n171), .B(n462), .Z(\ab[0][87] ) );
  AN2P U958 ( .A(n180), .B(n463), .Z(\ab[1][86] ) );
  AN2P U959 ( .A(n171), .B(n463), .Z(\ab[0][86] ) );
  AN2P U960 ( .A(n180), .B(n464), .Z(\ab[1][85] ) );
  AN2P U961 ( .A(n171), .B(n464), .Z(\ab[0][85] ) );
  AN2P U962 ( .A(n180), .B(n465), .Z(\ab[1][84] ) );
  AN2P U963 ( .A(n170), .B(n465), .Z(\ab[0][84] ) );
  AN2P U964 ( .A(n179), .B(n466), .Z(\ab[1][83] ) );
  AN2P U965 ( .A(n170), .B(n466), .Z(\ab[0][83] ) );
  AN2P U966 ( .A(n179), .B(n467), .Z(\ab[1][82] ) );
  AN2P U967 ( .A(n170), .B(n467), .Z(\ab[0][82] ) );
  AN2P U968 ( .A(n179), .B(n468), .Z(\ab[1][81] ) );
  AN2P U969 ( .A(n170), .B(n468), .Z(\ab[0][81] ) );
  AN2P U970 ( .A(n179), .B(n469), .Z(\ab[1][80] ) );
  AN2P U971 ( .A(n170), .B(n469), .Z(\ab[0][80] ) );
  AN2P U972 ( .A(n179), .B(n470), .Z(\ab[1][79] ) );
  AN2P U973 ( .A(n170), .B(n470), .Z(\ab[0][79] ) );
  AN2P U974 ( .A(n179), .B(n471), .Z(\ab[1][78] ) );
  AN2P U975 ( .A(n170), .B(n471), .Z(\ab[0][78] ) );
  AN2P U976 ( .A(n179), .B(n472), .Z(\ab[1][77] ) );
  AN2P U977 ( .A(n170), .B(n472), .Z(\ab[0][77] ) );
  AN2P U978 ( .A(n179), .B(n473), .Z(\ab[1][76] ) );
  AN2P U979 ( .A(n170), .B(n473), .Z(\ab[0][76] ) );
  AN2P U980 ( .A(n179), .B(n474), .Z(\ab[1][75] ) );
  AN2P U981 ( .A(n170), .B(n474), .Z(\ab[0][75] ) );
  AN2P U982 ( .A(n179), .B(n475), .Z(\ab[1][74] ) );
  AN2P U983 ( .A(n170), .B(n475), .Z(\ab[0][74] ) );
  AN2P U984 ( .A(n179), .B(n476), .Z(\ab[1][73] ) );
  AN2P U985 ( .A(n170), .B(n476), .Z(\ab[0][73] ) );
  AN2P U986 ( .A(n179), .B(n477), .Z(\ab[1][72] ) );
  AN2P U987 ( .A(n169), .B(n477), .Z(\ab[0][72] ) );
  AN2P U988 ( .A(n178), .B(n478), .Z(\ab[1][71] ) );
  AN2P U989 ( .A(n169), .B(n478), .Z(\ab[0][71] ) );
  AN2P U990 ( .A(n178), .B(n479), .Z(\ab[1][70] ) );
  AN2P U991 ( .A(n169), .B(n479), .Z(\ab[0][70] ) );
  AN2P U992 ( .A(n178), .B(n480), .Z(\ab[1][69] ) );
  AN2P U993 ( .A(n169), .B(n480), .Z(\ab[0][69] ) );
  AN2P U994 ( .A(n178), .B(n481), .Z(\ab[1][68] ) );
  AN2P U995 ( .A(n169), .B(n481), .Z(\ab[0][68] ) );
  AN2P U996 ( .A(n178), .B(n482), .Z(\ab[1][67] ) );
  AN2P U997 ( .A(n169), .B(n482), .Z(\ab[0][67] ) );
  AN2P U998 ( .A(n178), .B(n483), .Z(\ab[1][66] ) );
  AN2P U999 ( .A(n169), .B(n483), .Z(\ab[0][66] ) );
  AN2P U1000 ( .A(n178), .B(n484), .Z(\ab[1][65] ) );
  AN2P U1001 ( .A(n169), .B(n484), .Z(\ab[0][65] ) );
  AN2P U1002 ( .A(n178), .B(n485), .Z(\ab[1][64] ) );
  AN2P U1003 ( .A(n169), .B(n485), .Z(\ab[0][64] ) );
  AN2P U1004 ( .A(n178), .B(n486), .Z(\ab[1][63] ) );
  AN2P U1005 ( .A(n169), .B(n486), .Z(\ab[0][63] ) );
  AN2P U1006 ( .A(n178), .B(n487), .Z(\ab[1][62] ) );
  AN2P U1007 ( .A(n169), .B(n487), .Z(\ab[0][62] ) );
  AN2P U1008 ( .A(n178), .B(n488), .Z(\ab[1][61] ) );
  AN2P U1009 ( .A(n169), .B(n488), .Z(\ab[0][61] ) );
  AN2P U1010 ( .A(n178), .B(n489), .Z(\ab[1][60] ) );
  AN2P U1011 ( .A(n168), .B(n489), .Z(\ab[0][60] ) );
  AN2P U1012 ( .A(n177), .B(B[59]), .Z(\ab[1][59] ) );
  AN2P U1013 ( .A(n168), .B(B[59]), .Z(\ab[0][59] ) );
  AN2P U1014 ( .A(n177), .B(B[58]), .Z(\ab[1][58] ) );
  AN2P U1015 ( .A(n168), .B(B[58]), .Z(\ab[0][58] ) );
  AN2P U1016 ( .A(n177), .B(B[57]), .Z(\ab[1][57] ) );
  AN2P U1017 ( .A(n168), .B(B[57]), .Z(\ab[0][57] ) );
  AN2P U1018 ( .A(n177), .B(B[56]), .Z(\ab[1][56] ) );
  AN2P U1019 ( .A(n168), .B(B[56]), .Z(\ab[0][56] ) );
  AN2P U1020 ( .A(n177), .B(n490), .Z(\ab[1][55] ) );
  AN2P U1021 ( .A(n168), .B(n490), .Z(\ab[0][55] ) );
  AN2P U1022 ( .A(n177), .B(B[54]), .Z(\ab[1][54] ) );
  AN2P U1023 ( .A(n168), .B(B[54]), .Z(\ab[0][54] ) );
  AN2P U1024 ( .A(n177), .B(B[53]), .Z(\ab[1][53] ) );
  AN2P U1025 ( .A(n168), .B(B[53]), .Z(\ab[0][53] ) );
  AN2P U1026 ( .A(n177), .B(B[52]), .Z(\ab[1][52] ) );
  AN2P U1027 ( .A(n168), .B(B[52]), .Z(\ab[0][52] ) );
  AN2P U1028 ( .A(n177), .B(B[51]), .Z(\ab[1][51] ) );
  AN2P U1029 ( .A(n168), .B(B[51]), .Z(\ab[0][51] ) );
  AN2P U1030 ( .A(n177), .B(B[50]), .Z(\ab[1][50] ) );
  AN2P U1031 ( .A(n168), .B(B[50]), .Z(\ab[0][50] ) );
  AN2P U1032 ( .A(n177), .B(B[49]), .Z(\ab[1][49] ) );
  AN2P U1033 ( .A(n168), .B(B[49]), .Z(\ab[0][49] ) );
  AN2P U1034 ( .A(n177), .B(B[48]), .Z(\ab[1][48] ) );
  AN2P U1035 ( .A(n167), .B(B[48]), .Z(\ab[0][48] ) );
  AN2P U1036 ( .A(n176), .B(B[47]), .Z(\ab[1][47] ) );
  AN2P U1037 ( .A(n167), .B(B[47]), .Z(\ab[0][47] ) );
  AN2P U1038 ( .A(n176), .B(B[46]), .Z(\ab[1][46] ) );
  AN2P U1039 ( .A(n167), .B(B[46]), .Z(\ab[0][46] ) );
  AN2P U1040 ( .A(n176), .B(B[45]), .Z(\ab[1][45] ) );
  AN2P U1041 ( .A(n167), .B(B[45]), .Z(\ab[0][45] ) );
  AN2P U1042 ( .A(n176), .B(B[44]), .Z(\ab[1][44] ) );
  AN2P U1043 ( .A(n167), .B(B[44]), .Z(\ab[0][44] ) );
  AN2P U1044 ( .A(n176), .B(B[43]), .Z(\ab[1][43] ) );
  AN2P U1045 ( .A(n167), .B(B[43]), .Z(\ab[0][43] ) );
  AN2P U1046 ( .A(n176), .B(B[42]), .Z(\ab[1][42] ) );
  AN2P U1047 ( .A(n167), .B(B[42]), .Z(\ab[0][42] ) );
  AN2P U1048 ( .A(n176), .B(B[41]), .Z(\ab[1][41] ) );
  AN2P U1049 ( .A(n167), .B(B[41]), .Z(\ab[0][41] ) );
  AN2P U1050 ( .A(n176), .B(B[40]), .Z(\ab[1][40] ) );
  AN2P U1051 ( .A(n167), .B(B[40]), .Z(\ab[0][40] ) );
  AN2P U1052 ( .A(n176), .B(B[39]), .Z(\ab[1][39] ) );
  AN2P U1053 ( .A(n167), .B(B[39]), .Z(\ab[0][39] ) );
  AN2P U1054 ( .A(n176), .B(n453), .Z(\ab[1][38] ) );
  AN2P U1055 ( .A(n167), .B(n453), .Z(\ab[0][38] ) );
  AN2P U1056 ( .A(n176), .B(n449), .Z(\ab[1][37] ) );
  AN2P U1057 ( .A(n167), .B(n449), .Z(\ab[0][37] ) );
  AN2P U1058 ( .A(n176), .B(n445), .Z(\ab[1][36] ) );
  AN2P U1059 ( .A(n166), .B(n445), .Z(\ab[0][36] ) );
  AN2P U1060 ( .A(n175), .B(n441), .Z(\ab[1][35] ) );
  AN2P U1061 ( .A(n166), .B(n441), .Z(\ab[0][35] ) );
  AN2P U1062 ( .A(n175), .B(n437), .Z(\ab[1][34] ) );
  AN2P U1063 ( .A(n166), .B(n437), .Z(\ab[0][34] ) );
  AN2P U1064 ( .A(n175), .B(n433), .Z(\ab[1][33] ) );
  AN2P U1065 ( .A(n166), .B(n433), .Z(\ab[0][33] ) );
  AN2P U1066 ( .A(n175), .B(n429), .Z(\ab[1][32] ) );
  AN2P U1067 ( .A(n166), .B(n429), .Z(\ab[0][32] ) );
  AN2P U1068 ( .A(n175), .B(n425), .Z(\ab[1][31] ) );
  AN2P U1069 ( .A(n166), .B(n425), .Z(\ab[0][31] ) );
  AN2P U1070 ( .A(n175), .B(n421), .Z(\ab[1][30] ) );
  AN2P U1071 ( .A(n166), .B(n421), .Z(\ab[0][30] ) );
  AN2P U1072 ( .A(n175), .B(n417), .Z(\ab[1][29] ) );
  AN2P U1073 ( .A(n166), .B(n417), .Z(\ab[0][29] ) );
  AN2P U1074 ( .A(n175), .B(n413), .Z(\ab[1][28] ) );
  AN2P U1075 ( .A(n166), .B(n413), .Z(\ab[0][28] ) );
  AN2P U1076 ( .A(n175), .B(n409), .Z(\ab[1][27] ) );
  AN2P U1077 ( .A(n166), .B(n409), .Z(\ab[0][27] ) );
  AN2P U1078 ( .A(n175), .B(n405), .Z(\ab[1][26] ) );
  AN2P U1079 ( .A(n166), .B(n405), .Z(\ab[0][26] ) );
  AN2P U1080 ( .A(n175), .B(n401), .Z(\ab[1][25] ) );
  AN2P U1081 ( .A(n166), .B(n401), .Z(\ab[0][25] ) );
  AN2P U1082 ( .A(n175), .B(n397), .Z(\ab[1][24] ) );
  AN2P U1083 ( .A(n165), .B(n397), .Z(\ab[0][24] ) );
  AN2P U1084 ( .A(n174), .B(n393), .Z(\ab[1][23] ) );
  AN2P U1085 ( .A(n165), .B(n393), .Z(\ab[0][23] ) );
  AN2P U1086 ( .A(n174), .B(n389), .Z(\ab[1][22] ) );
  AN2P U1087 ( .A(n165), .B(n389), .Z(\ab[0][22] ) );
  AN2P U1088 ( .A(n174), .B(n385), .Z(\ab[1][21] ) );
  AN2P U1089 ( .A(n165), .B(n385), .Z(\ab[0][21] ) );
  AN2P U1090 ( .A(n174), .B(n381), .Z(\ab[1][20] ) );
  AN2P U1091 ( .A(n165), .B(n381), .Z(\ab[0][20] ) );
  AN2P U1092 ( .A(n174), .B(n377), .Z(\ab[1][19] ) );
  AN2P U1093 ( .A(n165), .B(n377), .Z(\ab[0][19] ) );
  AN2P U1094 ( .A(n174), .B(n373), .Z(\ab[1][18] ) );
  AN2P U1095 ( .A(n165), .B(n373), .Z(\ab[0][18] ) );
  AN2P U1096 ( .A(n174), .B(n369), .Z(\ab[1][17] ) );
  AN2P U1097 ( .A(n165), .B(n369), .Z(\ab[0][17] ) );
  AN2P U1098 ( .A(n174), .B(n365), .Z(\ab[1][16] ) );
  AN2P U1099 ( .A(n165), .B(n365), .Z(\ab[0][16] ) );
  AN2P U1100 ( .A(n174), .B(n361), .Z(\ab[1][15] ) );
  AN2P U1101 ( .A(n165), .B(n361), .Z(\ab[0][15] ) );
  AN2P U1102 ( .A(n174), .B(n357), .Z(\ab[1][14] ) );
  AN2P U1103 ( .A(n165), .B(n357), .Z(\ab[0][14] ) );
  AN2P U1104 ( .A(n174), .B(n353), .Z(\ab[1][13] ) );
  AN2P U1105 ( .A(n165), .B(n353), .Z(\ab[0][13] ) );
  AN2P U1106 ( .A(n174), .B(n349), .Z(\ab[1][12] ) );
  AN2P U1107 ( .A(n164), .B(n349), .Z(\ab[0][12] ) );
  AN2P U1108 ( .A(n173), .B(n345), .Z(\ab[1][11] ) );
  AN2P U1109 ( .A(n164), .B(n345), .Z(\ab[0][11] ) );
  AN2P U1110 ( .A(n173), .B(n341), .Z(\ab[1][10] ) );
  AN2P U1111 ( .A(n164), .B(n341), .Z(\ab[0][10] ) );
  AN2P U1112 ( .A(n173), .B(n337), .Z(\ab[1][9] ) );
  AN2P U1113 ( .A(n164), .B(n337), .Z(\ab[0][9] ) );
  AN2P U1114 ( .A(n173), .B(n333), .Z(\ab[1][8] ) );
  AN2P U1115 ( .A(n164), .B(n333), .Z(\ab[0][8] ) );
  AN2P U1116 ( .A(n173), .B(n329), .Z(\ab[1][7] ) );
  AN2P U1117 ( .A(n164), .B(n329), .Z(\ab[0][7] ) );
  AN2P U1118 ( .A(n173), .B(n325), .Z(\ab[1][6] ) );
  AN2P U1119 ( .A(n164), .B(n325), .Z(\ab[0][6] ) );
  AN2P U1120 ( .A(n173), .B(n321), .Z(\ab[1][5] ) );
  AN2P U1121 ( .A(n164), .B(n321), .Z(\ab[0][5] ) );
  AN2P U1122 ( .A(n173), .B(n317), .Z(\ab[1][4] ) );
  AN2P U1123 ( .A(n164), .B(n317), .Z(\ab[0][4] ) );
  AN2P U1124 ( .A(n173), .B(n313), .Z(\ab[1][3] ) );
  AN2P U1125 ( .A(n164), .B(n313), .Z(\ab[0][3] ) );
  AN2P U1126 ( .A(n173), .B(n309), .Z(\ab[1][2] ) );
  AN2P U1127 ( .A(n164), .B(n309), .Z(\ab[0][2] ) );
  AN2P U1128 ( .A(n189), .B(n455), .Z(\ab[2][94] ) );
  AN2P U1129 ( .A(n173), .B(n491), .Z(\ab[1][95] ) );
  AN2P U1130 ( .A(n189), .B(n456), .Z(\ab[2][93] ) );
  AN2P U1131 ( .A(n189), .B(n457), .Z(\ab[2][92] ) );
  AN2P U1132 ( .A(n189), .B(n458), .Z(\ab[2][91] ) );
  AN2P U1133 ( .A(n189), .B(n459), .Z(\ab[2][90] ) );
  AN2P U1134 ( .A(n189), .B(n460), .Z(\ab[2][89] ) );
  AN2P U1135 ( .A(n189), .B(n461), .Z(\ab[2][88] ) );
  AN2P U1136 ( .A(n189), .B(n462), .Z(\ab[2][87] ) );
  AN2P U1137 ( .A(n189), .B(n463), .Z(\ab[2][86] ) );
  AN2P U1138 ( .A(n189), .B(n464), .Z(\ab[2][85] ) );
  AN2P U1139 ( .A(n189), .B(n465), .Z(\ab[2][84] ) );
  AN2P U1140 ( .A(n189), .B(n466), .Z(\ab[2][83] ) );
  AN2P U1141 ( .A(n188), .B(n467), .Z(\ab[2][82] ) );
  AN2P U1142 ( .A(n188), .B(n468), .Z(\ab[2][81] ) );
  AN2P U1143 ( .A(n188), .B(n469), .Z(\ab[2][80] ) );
  AN2P U1144 ( .A(n188), .B(n470), .Z(\ab[2][79] ) );
  AN2P U1145 ( .A(n188), .B(n471), .Z(\ab[2][78] ) );
  AN2P U1146 ( .A(n188), .B(n472), .Z(\ab[2][77] ) );
  AN2P U1147 ( .A(n188), .B(n473), .Z(\ab[2][76] ) );
  AN2P U1148 ( .A(n188), .B(n474), .Z(\ab[2][75] ) );
  AN2P U1149 ( .A(n188), .B(n475), .Z(\ab[2][74] ) );
  AN2P U1150 ( .A(n188), .B(n476), .Z(\ab[2][73] ) );
  AN2P U1151 ( .A(n188), .B(n477), .Z(\ab[2][72] ) );
  AN2P U1152 ( .A(n188), .B(n478), .Z(\ab[2][71] ) );
  AN2P U1153 ( .A(n187), .B(n479), .Z(\ab[2][70] ) );
  AN2P U1154 ( .A(n187), .B(n480), .Z(\ab[2][69] ) );
  AN2P U1155 ( .A(n187), .B(n481), .Z(\ab[2][68] ) );
  AN2P U1156 ( .A(n187), .B(n482), .Z(\ab[2][67] ) );
  AN2P U1157 ( .A(n187), .B(n483), .Z(\ab[2][66] ) );
  AN2P U1158 ( .A(n187), .B(n484), .Z(\ab[2][65] ) );
  AN2P U1159 ( .A(n187), .B(n485), .Z(\ab[2][64] ) );
  AN2P U1160 ( .A(n187), .B(n486), .Z(\ab[2][63] ) );
  AN2P U1161 ( .A(n187), .B(n487), .Z(\ab[2][62] ) );
  AN2P U1162 ( .A(n187), .B(n488), .Z(\ab[2][61] ) );
  AN2P U1163 ( .A(n187), .B(n489), .Z(\ab[2][60] ) );
  AN2P U1164 ( .A(n187), .B(B[59]), .Z(\ab[2][59] ) );
  AN2P U1165 ( .A(n186), .B(B[58]), .Z(\ab[2][58] ) );
  AN2P U1166 ( .A(n186), .B(B[57]), .Z(\ab[2][57] ) );
  AN2P U1167 ( .A(n186), .B(B[56]), .Z(\ab[2][56] ) );
  AN2P U1168 ( .A(n186), .B(n490), .Z(\ab[2][55] ) );
  AN2P U1169 ( .A(n186), .B(B[54]), .Z(\ab[2][54] ) );
  AN2P U1170 ( .A(n186), .B(B[53]), .Z(\ab[2][53] ) );
  AN2P U1171 ( .A(n186), .B(B[52]), .Z(\ab[2][52] ) );
  AN2P U1172 ( .A(n186), .B(B[51]), .Z(\ab[2][51] ) );
  AN2P U1173 ( .A(n186), .B(B[50]), .Z(\ab[2][50] ) );
  AN2P U1174 ( .A(n186), .B(B[49]), .Z(\ab[2][49] ) );
  AN2P U1175 ( .A(n186), .B(B[48]), .Z(\ab[2][48] ) );
  AN2P U1176 ( .A(n186), .B(B[47]), .Z(\ab[2][47] ) );
  AN2P U1177 ( .A(n185), .B(B[46]), .Z(\ab[2][46] ) );
  AN2P U1178 ( .A(n185), .B(B[45]), .Z(\ab[2][45] ) );
  AN2P U1179 ( .A(n185), .B(B[44]), .Z(\ab[2][44] ) );
  AN2P U1180 ( .A(n185), .B(B[43]), .Z(\ab[2][43] ) );
  AN2P U1181 ( .A(n185), .B(B[42]), .Z(\ab[2][42] ) );
  AN2P U1182 ( .A(n185), .B(B[41]), .Z(\ab[2][41] ) );
  AN2P U1183 ( .A(n185), .B(B[40]), .Z(\ab[2][40] ) );
  AN2P U1184 ( .A(n185), .B(B[39]), .Z(\ab[2][39] ) );
  AN2P U1185 ( .A(n185), .B(n453), .Z(\ab[2][38] ) );
  AN2P U1186 ( .A(n185), .B(n449), .Z(\ab[2][37] ) );
  AN2P U1187 ( .A(n185), .B(n445), .Z(\ab[2][36] ) );
  AN2P U1188 ( .A(n185), .B(n441), .Z(\ab[2][35] ) );
  AN2P U1189 ( .A(n184), .B(n437), .Z(\ab[2][34] ) );
  AN2P U1190 ( .A(n184), .B(n433), .Z(\ab[2][33] ) );
  AN2P U1191 ( .A(n184), .B(n429), .Z(\ab[2][32] ) );
  AN2P U1192 ( .A(n184), .B(n425), .Z(\ab[2][31] ) );
  AN2P U1193 ( .A(n184), .B(n421), .Z(\ab[2][30] ) );
  AN2P U1194 ( .A(n184), .B(n417), .Z(\ab[2][29] ) );
  AN2P U1195 ( .A(n184), .B(n413), .Z(\ab[2][28] ) );
  AN2P U1196 ( .A(n184), .B(n409), .Z(\ab[2][27] ) );
  AN2P U1197 ( .A(n184), .B(n405), .Z(\ab[2][26] ) );
  AN2P U1198 ( .A(n184), .B(n401), .Z(\ab[2][25] ) );
  AN2P U1199 ( .A(n184), .B(n397), .Z(\ab[2][24] ) );
  AN2P U1200 ( .A(n184), .B(n393), .Z(\ab[2][23] ) );
  AN2P U1201 ( .A(n183), .B(n389), .Z(\ab[2][22] ) );
  AN2P U1202 ( .A(n183), .B(n385), .Z(\ab[2][21] ) );
  AN2P U1203 ( .A(n183), .B(n381), .Z(\ab[2][20] ) );
  AN2P U1204 ( .A(n183), .B(n377), .Z(\ab[2][19] ) );
  AN2P U1205 ( .A(n183), .B(n373), .Z(\ab[2][18] ) );
  AN2P U1206 ( .A(n183), .B(n369), .Z(\ab[2][17] ) );
  AN2P U1207 ( .A(n183), .B(n365), .Z(\ab[2][16] ) );
  AN2P U1208 ( .A(n183), .B(n361), .Z(\ab[2][15] ) );
  AN2P U1209 ( .A(n183), .B(n357), .Z(\ab[2][14] ) );
  AN2P U1210 ( .A(n183), .B(n353), .Z(\ab[2][13] ) );
  AN2P U1211 ( .A(n183), .B(n349), .Z(\ab[2][12] ) );
  AN2P U1212 ( .A(n183), .B(n345), .Z(\ab[2][11] ) );
  AN2P U1213 ( .A(n182), .B(n341), .Z(\ab[2][10] ) );
  AN2P U1214 ( .A(n182), .B(n337), .Z(\ab[2][9] ) );
  AN2P U1215 ( .A(n182), .B(n333), .Z(\ab[2][8] ) );
  AN2P U1216 ( .A(n182), .B(n329), .Z(\ab[2][7] ) );
  AN2P U1217 ( .A(n182), .B(n325), .Z(\ab[2][6] ) );
  AN2P U1218 ( .A(n182), .B(n321), .Z(\ab[2][5] ) );
  AN2P U1219 ( .A(n182), .B(n317), .Z(\ab[2][4] ) );
  AN2P U1220 ( .A(n182), .B(n313), .Z(\ab[2][3] ) );
  AN2P U1221 ( .A(n182), .B(n309), .Z(\ab[2][2] ) );
  AN2P U1222 ( .A(n182), .B(n305), .Z(\ab[2][1] ) );
  AN2P U1223 ( .A(n182), .B(n301), .Z(\ab[2][0] ) );
  AN3 U1224 ( .A(n164), .B(n301), .C(n3), .Z(\CARRYB[1][0] ) );
  AN2P U1225 ( .A(n198), .B(n455), .Z(\ab[3][94] ) );
  AN2P U1226 ( .A(n182), .B(n491), .Z(\ab[2][95] ) );
  AN2P U1227 ( .A(n198), .B(n456), .Z(\ab[3][93] ) );
  AN2P U1228 ( .A(n198), .B(n457), .Z(\ab[3][92] ) );
  AN2P U1229 ( .A(n198), .B(n458), .Z(\ab[3][91] ) );
  AN2P U1230 ( .A(n198), .B(n459), .Z(\ab[3][90] ) );
  AN2P U1231 ( .A(n198), .B(n460), .Z(\ab[3][89] ) );
  AN2P U1232 ( .A(n198), .B(n461), .Z(\ab[3][88] ) );
  AN2P U1233 ( .A(n198), .B(n462), .Z(\ab[3][87] ) );
  AN2P U1234 ( .A(n198), .B(n463), .Z(\ab[3][86] ) );
  AN2P U1235 ( .A(n198), .B(n464), .Z(\ab[3][85] ) );
  AN2P U1236 ( .A(n198), .B(n465), .Z(\ab[3][84] ) );
  AN2P U1237 ( .A(n198), .B(n466), .Z(\ab[3][83] ) );
  AN2P U1238 ( .A(n197), .B(n467), .Z(\ab[3][82] ) );
  AN2P U1239 ( .A(n197), .B(n468), .Z(\ab[3][81] ) );
  AN2P U1240 ( .A(n197), .B(n469), .Z(\ab[3][80] ) );
  AN2P U1241 ( .A(n197), .B(n470), .Z(\ab[3][79] ) );
  AN2P U1242 ( .A(n197), .B(n471), .Z(\ab[3][78] ) );
  AN2P U1243 ( .A(n197), .B(n472), .Z(\ab[3][77] ) );
  AN2P U1244 ( .A(n197), .B(n473), .Z(\ab[3][76] ) );
  AN2P U1245 ( .A(n197), .B(n474), .Z(\ab[3][75] ) );
  AN2P U1246 ( .A(n197), .B(n475), .Z(\ab[3][74] ) );
  AN2P U1247 ( .A(n197), .B(n476), .Z(\ab[3][73] ) );
  AN2P U1248 ( .A(n197), .B(n477), .Z(\ab[3][72] ) );
  AN2P U1249 ( .A(n197), .B(n478), .Z(\ab[3][71] ) );
  AN2P U1250 ( .A(n196), .B(n479), .Z(\ab[3][70] ) );
  AN2P U1251 ( .A(n196), .B(n480), .Z(\ab[3][69] ) );
  AN2P U1252 ( .A(n196), .B(n481), .Z(\ab[3][68] ) );
  AN2P U1253 ( .A(n196), .B(n482), .Z(\ab[3][67] ) );
  AN2P U1254 ( .A(n196), .B(n483), .Z(\ab[3][66] ) );
  AN2P U1255 ( .A(n196), .B(n484), .Z(\ab[3][65] ) );
  AN2P U1256 ( .A(n196), .B(n485), .Z(\ab[3][64] ) );
  AN2P U1257 ( .A(n196), .B(n486), .Z(\ab[3][63] ) );
  AN2P U1258 ( .A(n196), .B(n487), .Z(\ab[3][62] ) );
  AN2P U1259 ( .A(n196), .B(n488), .Z(\ab[3][61] ) );
  AN2P U1260 ( .A(n196), .B(n489), .Z(\ab[3][60] ) );
  AN2P U1261 ( .A(n196), .B(B[59]), .Z(\ab[3][59] ) );
  AN2P U1262 ( .A(n195), .B(B[58]), .Z(\ab[3][58] ) );
  AN2P U1263 ( .A(n195), .B(B[57]), .Z(\ab[3][57] ) );
  AN2P U1264 ( .A(n195), .B(B[56]), .Z(\ab[3][56] ) );
  AN2P U1265 ( .A(n195), .B(n490), .Z(\ab[3][55] ) );
  AN2P U1266 ( .A(n195), .B(B[54]), .Z(\ab[3][54] ) );
  AN2P U1267 ( .A(n195), .B(B[53]), .Z(\ab[3][53] ) );
  AN2P U1268 ( .A(n195), .B(B[52]), .Z(\ab[3][52] ) );
  AN2P U1269 ( .A(n195), .B(B[51]), .Z(\ab[3][51] ) );
  AN2P U1270 ( .A(n195), .B(B[50]), .Z(\ab[3][50] ) );
  AN2P U1271 ( .A(n195), .B(B[49]), .Z(\ab[3][49] ) );
  AN2P U1272 ( .A(n195), .B(B[48]), .Z(\ab[3][48] ) );
  AN2P U1273 ( .A(n195), .B(B[47]), .Z(\ab[3][47] ) );
  AN2P U1274 ( .A(n194), .B(B[46]), .Z(\ab[3][46] ) );
  AN2P U1275 ( .A(n194), .B(B[45]), .Z(\ab[3][45] ) );
  AN2P U1276 ( .A(n194), .B(B[44]), .Z(\ab[3][44] ) );
  AN2P U1277 ( .A(n194), .B(B[43]), .Z(\ab[3][43] ) );
  AN2P U1278 ( .A(n194), .B(B[42]), .Z(\ab[3][42] ) );
  AN2P U1279 ( .A(n194), .B(B[41]), .Z(\ab[3][41] ) );
  AN2P U1280 ( .A(n194), .B(B[40]), .Z(\ab[3][40] ) );
  AN2P U1281 ( .A(n194), .B(B[39]), .Z(\ab[3][39] ) );
  AN2P U1282 ( .A(n194), .B(n453), .Z(\ab[3][38] ) );
  AN2P U1283 ( .A(n194), .B(n449), .Z(\ab[3][37] ) );
  AN2P U1284 ( .A(n194), .B(n445), .Z(\ab[3][36] ) );
  AN2P U1285 ( .A(n194), .B(n441), .Z(\ab[3][35] ) );
  AN2P U1286 ( .A(n193), .B(n437), .Z(\ab[3][34] ) );
  AN2P U1287 ( .A(n193), .B(n433), .Z(\ab[3][33] ) );
  AN2P U1288 ( .A(n193), .B(n429), .Z(\ab[3][32] ) );
  AN2P U1289 ( .A(n193), .B(n425), .Z(\ab[3][31] ) );
  AN2P U1290 ( .A(n193), .B(n421), .Z(\ab[3][30] ) );
  AN2P U1291 ( .A(n193), .B(n417), .Z(\ab[3][29] ) );
  AN2P U1292 ( .A(n193), .B(n413), .Z(\ab[3][28] ) );
  AN2P U1293 ( .A(n193), .B(n409), .Z(\ab[3][27] ) );
  AN2P U1294 ( .A(n193), .B(n405), .Z(\ab[3][26] ) );
  AN2P U1295 ( .A(n193), .B(n401), .Z(\ab[3][25] ) );
  AN2P U1296 ( .A(n193), .B(n397), .Z(\ab[3][24] ) );
  AN2P U1297 ( .A(n193), .B(n393), .Z(\ab[3][23] ) );
  AN2P U1298 ( .A(n192), .B(n389), .Z(\ab[3][22] ) );
  AN2P U1299 ( .A(n192), .B(n385), .Z(\ab[3][21] ) );
  AN2P U1300 ( .A(n192), .B(n381), .Z(\ab[3][20] ) );
  AN2P U1301 ( .A(n192), .B(n377), .Z(\ab[3][19] ) );
  AN2P U1302 ( .A(n192), .B(n373), .Z(\ab[3][18] ) );
  AN2P U1303 ( .A(n192), .B(n369), .Z(\ab[3][17] ) );
  AN2P U1304 ( .A(n192), .B(n365), .Z(\ab[3][16] ) );
  AN2P U1305 ( .A(n192), .B(n361), .Z(\ab[3][15] ) );
  AN2P U1306 ( .A(n192), .B(n357), .Z(\ab[3][14] ) );
  AN2P U1307 ( .A(n192), .B(n353), .Z(\ab[3][13] ) );
  AN2P U1308 ( .A(n192), .B(n349), .Z(\ab[3][12] ) );
  AN2P U1309 ( .A(n192), .B(n345), .Z(\ab[3][11] ) );
  AN2P U1310 ( .A(n191), .B(n341), .Z(\ab[3][10] ) );
  AN2P U1311 ( .A(n191), .B(n337), .Z(\ab[3][9] ) );
  AN2P U1312 ( .A(n191), .B(n333), .Z(\ab[3][8] ) );
  AN2P U1313 ( .A(n191), .B(n329), .Z(\ab[3][7] ) );
  AN2P U1314 ( .A(n191), .B(n325), .Z(\ab[3][6] ) );
  AN2P U1315 ( .A(n191), .B(n321), .Z(\ab[3][5] ) );
  AN2P U1316 ( .A(n191), .B(n317), .Z(\ab[3][4] ) );
  AN2P U1317 ( .A(n191), .B(n313), .Z(\ab[3][3] ) );
  AN2P U1318 ( .A(n191), .B(n309), .Z(\ab[3][2] ) );
  AN2P U1319 ( .A(n191), .B(n305), .Z(\ab[3][1] ) );
  AN2P U1320 ( .A(n191), .B(n301), .Z(\ab[3][0] ) );
  AN2P U1321 ( .A(n207), .B(n455), .Z(\ab[4][94] ) );
  AN2P U1322 ( .A(n191), .B(n491), .Z(\ab[3][95] ) );
  AN2P U1323 ( .A(n207), .B(n456), .Z(\ab[4][93] ) );
  AN2P U1324 ( .A(n207), .B(n457), .Z(\ab[4][92] ) );
  AN2P U1325 ( .A(n207), .B(n458), .Z(\ab[4][91] ) );
  AN2P U1326 ( .A(n207), .B(n459), .Z(\ab[4][90] ) );
  AN2P U1327 ( .A(n207), .B(n460), .Z(\ab[4][89] ) );
  AN2P U1328 ( .A(n207), .B(n461), .Z(\ab[4][88] ) );
  AN2P U1329 ( .A(n207), .B(n462), .Z(\ab[4][87] ) );
  AN2P U1330 ( .A(n207), .B(n463), .Z(\ab[4][86] ) );
  AN2P U1331 ( .A(n207), .B(n464), .Z(\ab[4][85] ) );
  AN2P U1332 ( .A(n207), .B(n465), .Z(\ab[4][84] ) );
  AN2P U1333 ( .A(n207), .B(n466), .Z(\ab[4][83] ) );
  AN2P U1334 ( .A(n206), .B(n467), .Z(\ab[4][82] ) );
  AN2P U1335 ( .A(n206), .B(n468), .Z(\ab[4][81] ) );
  AN2P U1336 ( .A(n206), .B(n469), .Z(\ab[4][80] ) );
  AN2P U1337 ( .A(n206), .B(n470), .Z(\ab[4][79] ) );
  AN2P U1338 ( .A(n206), .B(n471), .Z(\ab[4][78] ) );
  AN2P U1339 ( .A(n206), .B(n472), .Z(\ab[4][77] ) );
  AN2P U1340 ( .A(n206), .B(n473), .Z(\ab[4][76] ) );
  AN2P U1341 ( .A(n206), .B(n474), .Z(\ab[4][75] ) );
  AN2P U1342 ( .A(n206), .B(n475), .Z(\ab[4][74] ) );
  AN2P U1343 ( .A(n206), .B(n476), .Z(\ab[4][73] ) );
  AN2P U1344 ( .A(n206), .B(n477), .Z(\ab[4][72] ) );
  AN2P U1345 ( .A(n206), .B(n478), .Z(\ab[4][71] ) );
  AN2P U1346 ( .A(n205), .B(n479), .Z(\ab[4][70] ) );
  AN2P U1347 ( .A(n205), .B(n480), .Z(\ab[4][69] ) );
  AN2P U1348 ( .A(n205), .B(n481), .Z(\ab[4][68] ) );
  AN2P U1349 ( .A(n205), .B(n482), .Z(\ab[4][67] ) );
  AN2P U1350 ( .A(n205), .B(n483), .Z(\ab[4][66] ) );
  AN2P U1351 ( .A(n205), .B(n484), .Z(\ab[4][65] ) );
  AN2P U1352 ( .A(n205), .B(n485), .Z(\ab[4][64] ) );
  AN2P U1353 ( .A(n205), .B(n486), .Z(\ab[4][63] ) );
  AN2P U1354 ( .A(n205), .B(n487), .Z(\ab[4][62] ) );
  AN2P U1355 ( .A(n205), .B(n488), .Z(\ab[4][61] ) );
  AN2P U1356 ( .A(n205), .B(n489), .Z(\ab[4][60] ) );
  AN2P U1357 ( .A(n205), .B(B[59]), .Z(\ab[4][59] ) );
  AN2P U1358 ( .A(n204), .B(B[58]), .Z(\ab[4][58] ) );
  AN2P U1359 ( .A(n204), .B(B[57]), .Z(\ab[4][57] ) );
  AN2P U1360 ( .A(n204), .B(B[56]), .Z(\ab[4][56] ) );
  AN2P U1361 ( .A(n204), .B(n490), .Z(\ab[4][55] ) );
  AN2P U1362 ( .A(n204), .B(B[54]), .Z(\ab[4][54] ) );
  AN2P U1363 ( .A(n204), .B(B[53]), .Z(\ab[4][53] ) );
  AN2P U1364 ( .A(n204), .B(B[52]), .Z(\ab[4][52] ) );
  AN2P U1365 ( .A(n204), .B(B[51]), .Z(\ab[4][51] ) );
  AN2P U1366 ( .A(n204), .B(B[50]), .Z(\ab[4][50] ) );
  AN2P U1367 ( .A(n204), .B(B[49]), .Z(\ab[4][49] ) );
  AN2P U1368 ( .A(n204), .B(B[48]), .Z(\ab[4][48] ) );
  AN2P U1369 ( .A(n204), .B(B[47]), .Z(\ab[4][47] ) );
  AN2P U1370 ( .A(n203), .B(B[46]), .Z(\ab[4][46] ) );
  AN2P U1371 ( .A(n203), .B(B[45]), .Z(\ab[4][45] ) );
  AN2P U1372 ( .A(n203), .B(B[44]), .Z(\ab[4][44] ) );
  AN2P U1373 ( .A(n203), .B(B[43]), .Z(\ab[4][43] ) );
  AN2P U1374 ( .A(n203), .B(B[42]), .Z(\ab[4][42] ) );
  AN2P U1375 ( .A(n203), .B(B[41]), .Z(\ab[4][41] ) );
  AN2P U1376 ( .A(n203), .B(B[40]), .Z(\ab[4][40] ) );
  AN2P U1377 ( .A(n203), .B(B[39]), .Z(\ab[4][39] ) );
  AN2P U1378 ( .A(n203), .B(n453), .Z(\ab[4][38] ) );
  AN2P U1379 ( .A(n203), .B(n449), .Z(\ab[4][37] ) );
  AN2P U1380 ( .A(n203), .B(n445), .Z(\ab[4][36] ) );
  AN2P U1381 ( .A(n203), .B(n441), .Z(\ab[4][35] ) );
  AN2P U1382 ( .A(n202), .B(n437), .Z(\ab[4][34] ) );
  AN2P U1383 ( .A(n202), .B(n433), .Z(\ab[4][33] ) );
  AN2P U1384 ( .A(n202), .B(n429), .Z(\ab[4][32] ) );
  AN2P U1385 ( .A(n202), .B(n425), .Z(\ab[4][31] ) );
  AN2P U1386 ( .A(n202), .B(n421), .Z(\ab[4][30] ) );
  AN2P U1387 ( .A(n202), .B(n417), .Z(\ab[4][29] ) );
  AN2P U1388 ( .A(n202), .B(n413), .Z(\ab[4][28] ) );
  AN2P U1389 ( .A(n202), .B(n409), .Z(\ab[4][27] ) );
  AN2P U1390 ( .A(n202), .B(n405), .Z(\ab[4][26] ) );
  AN2P U1391 ( .A(n202), .B(n401), .Z(\ab[4][25] ) );
  AN2P U1392 ( .A(n202), .B(n397), .Z(\ab[4][24] ) );
  AN2P U1393 ( .A(n202), .B(n393), .Z(\ab[4][23] ) );
  AN2P U1394 ( .A(n201), .B(n389), .Z(\ab[4][22] ) );
  AN2P U1395 ( .A(n201), .B(n385), .Z(\ab[4][21] ) );
  AN2P U1396 ( .A(n201), .B(n381), .Z(\ab[4][20] ) );
  AN2P U1397 ( .A(n201), .B(n377), .Z(\ab[4][19] ) );
  AN2P U1398 ( .A(n201), .B(n373), .Z(\ab[4][18] ) );
  AN2P U1399 ( .A(n201), .B(n369), .Z(\ab[4][17] ) );
  AN2P U1400 ( .A(n201), .B(n365), .Z(\ab[4][16] ) );
  AN2P U1401 ( .A(n201), .B(n361), .Z(\ab[4][15] ) );
  AN2P U1402 ( .A(n201), .B(n357), .Z(\ab[4][14] ) );
  AN2P U1403 ( .A(n201), .B(n353), .Z(\ab[4][13] ) );
  AN2P U1404 ( .A(n201), .B(n349), .Z(\ab[4][12] ) );
  AN2P U1405 ( .A(n201), .B(n345), .Z(\ab[4][11] ) );
  AN2P U1406 ( .A(n200), .B(n341), .Z(\ab[4][10] ) );
  AN2P U1407 ( .A(n200), .B(n337), .Z(\ab[4][9] ) );
  AN2P U1408 ( .A(n200), .B(n333), .Z(\ab[4][8] ) );
  AN2P U1409 ( .A(n200), .B(n329), .Z(\ab[4][7] ) );
  AN2P U1410 ( .A(n200), .B(n325), .Z(\ab[4][6] ) );
  AN2P U1411 ( .A(n200), .B(n321), .Z(\ab[4][5] ) );
  AN2P U1412 ( .A(n200), .B(n317), .Z(\ab[4][4] ) );
  AN2P U1413 ( .A(n200), .B(n313), .Z(\ab[4][3] ) );
  AN2P U1414 ( .A(n200), .B(n309), .Z(\ab[4][2] ) );
  AN2P U1415 ( .A(n200), .B(n305), .Z(\ab[4][1] ) );
  AN2P U1416 ( .A(n200), .B(n301), .Z(\ab[4][0] ) );
  AN2P U1417 ( .A(n216), .B(n455), .Z(\ab[5][94] ) );
  AN2P U1418 ( .A(n200), .B(n491), .Z(\ab[4][95] ) );
  AN2P U1419 ( .A(n216), .B(n456), .Z(\ab[5][93] ) );
  AN2P U1420 ( .A(n216), .B(n457), .Z(\ab[5][92] ) );
  AN2P U1421 ( .A(n216), .B(n458), .Z(\ab[5][91] ) );
  AN2P U1422 ( .A(n216), .B(n459), .Z(\ab[5][90] ) );
  AN2P U1423 ( .A(n216), .B(n460), .Z(\ab[5][89] ) );
  AN2P U1424 ( .A(n216), .B(n461), .Z(\ab[5][88] ) );
  AN2P U1425 ( .A(n216), .B(n462), .Z(\ab[5][87] ) );
  AN2P U1426 ( .A(n216), .B(n463), .Z(\ab[5][86] ) );
  AN2P U1427 ( .A(n216), .B(n464), .Z(\ab[5][85] ) );
  AN2P U1428 ( .A(n216), .B(n465), .Z(\ab[5][84] ) );
  AN2P U1429 ( .A(n216), .B(n466), .Z(\ab[5][83] ) );
  AN2P U1430 ( .A(n215), .B(n467), .Z(\ab[5][82] ) );
  AN2P U1431 ( .A(n215), .B(n468), .Z(\ab[5][81] ) );
  AN2P U1432 ( .A(n215), .B(n469), .Z(\ab[5][80] ) );
  AN2P U1433 ( .A(n215), .B(n470), .Z(\ab[5][79] ) );
  AN2P U1434 ( .A(n215), .B(n471), .Z(\ab[5][78] ) );
  AN2P U1435 ( .A(n215), .B(n472), .Z(\ab[5][77] ) );
  AN2P U1436 ( .A(n215), .B(n473), .Z(\ab[5][76] ) );
  AN2P U1437 ( .A(n215), .B(n474), .Z(\ab[5][75] ) );
  AN2P U1438 ( .A(n215), .B(n475), .Z(\ab[5][74] ) );
  AN2P U1439 ( .A(n215), .B(n476), .Z(\ab[5][73] ) );
  AN2P U1440 ( .A(n215), .B(n477), .Z(\ab[5][72] ) );
  AN2P U1441 ( .A(n215), .B(n478), .Z(\ab[5][71] ) );
  AN2P U1442 ( .A(n214), .B(n479), .Z(\ab[5][70] ) );
  AN2P U1443 ( .A(n214), .B(n480), .Z(\ab[5][69] ) );
  AN2P U1444 ( .A(n214), .B(n481), .Z(\ab[5][68] ) );
  AN2P U1445 ( .A(n214), .B(n482), .Z(\ab[5][67] ) );
  AN2P U1446 ( .A(n214), .B(n483), .Z(\ab[5][66] ) );
  AN2P U1447 ( .A(n214), .B(n484), .Z(\ab[5][65] ) );
  AN2P U1448 ( .A(n214), .B(n485), .Z(\ab[5][64] ) );
  AN2P U1449 ( .A(n214), .B(n486), .Z(\ab[5][63] ) );
  AN2P U1450 ( .A(n214), .B(n487), .Z(\ab[5][62] ) );
  AN2P U1451 ( .A(n214), .B(n488), .Z(\ab[5][61] ) );
  AN2P U1452 ( .A(n214), .B(n489), .Z(\ab[5][60] ) );
  AN2P U1453 ( .A(n214), .B(B[59]), .Z(\ab[5][59] ) );
  AN2P U1454 ( .A(n213), .B(B[58]), .Z(\ab[5][58] ) );
  AN2P U1455 ( .A(n213), .B(B[57]), .Z(\ab[5][57] ) );
  AN2P U1456 ( .A(n213), .B(B[56]), .Z(\ab[5][56] ) );
  AN2P U1457 ( .A(n213), .B(n490), .Z(\ab[5][55] ) );
  AN2P U1458 ( .A(n213), .B(B[54]), .Z(\ab[5][54] ) );
  AN2P U1459 ( .A(n213), .B(B[53]), .Z(\ab[5][53] ) );
  AN2P U1460 ( .A(n213), .B(B[52]), .Z(\ab[5][52] ) );
  AN2P U1461 ( .A(n213), .B(B[51]), .Z(\ab[5][51] ) );
  AN2P U1462 ( .A(n213), .B(B[50]), .Z(\ab[5][50] ) );
  AN2P U1463 ( .A(n213), .B(B[49]), .Z(\ab[5][49] ) );
  AN2P U1464 ( .A(n213), .B(B[48]), .Z(\ab[5][48] ) );
  AN2P U1465 ( .A(n213), .B(B[47]), .Z(\ab[5][47] ) );
  AN2P U1466 ( .A(n212), .B(B[46]), .Z(\ab[5][46] ) );
  AN2P U1467 ( .A(n212), .B(B[45]), .Z(\ab[5][45] ) );
  AN2P U1468 ( .A(n212), .B(B[44]), .Z(\ab[5][44] ) );
  AN2P U1469 ( .A(n212), .B(B[43]), .Z(\ab[5][43] ) );
  AN2P U1470 ( .A(n212), .B(B[42]), .Z(\ab[5][42] ) );
  AN2P U1471 ( .A(n212), .B(B[41]), .Z(\ab[5][41] ) );
  AN2P U1472 ( .A(n212), .B(B[40]), .Z(\ab[5][40] ) );
  AN2P U1473 ( .A(n212), .B(B[39]), .Z(\ab[5][39] ) );
  AN2P U1474 ( .A(n212), .B(n453), .Z(\ab[5][38] ) );
  AN2P U1475 ( .A(n212), .B(n449), .Z(\ab[5][37] ) );
  AN2P U1476 ( .A(n212), .B(n445), .Z(\ab[5][36] ) );
  AN2P U1477 ( .A(n212), .B(n441), .Z(\ab[5][35] ) );
  AN2P U1478 ( .A(n211), .B(n437), .Z(\ab[5][34] ) );
  AN2P U1479 ( .A(n211), .B(n433), .Z(\ab[5][33] ) );
  AN2P U1480 ( .A(n211), .B(n429), .Z(\ab[5][32] ) );
  AN2P U1481 ( .A(n211), .B(n425), .Z(\ab[5][31] ) );
  AN2P U1482 ( .A(n211), .B(n421), .Z(\ab[5][30] ) );
  AN2P U1483 ( .A(n211), .B(n417), .Z(\ab[5][29] ) );
  AN2P U1484 ( .A(n211), .B(n413), .Z(\ab[5][28] ) );
  AN2P U1485 ( .A(n211), .B(n409), .Z(\ab[5][27] ) );
  AN2P U1486 ( .A(n211), .B(n405), .Z(\ab[5][26] ) );
  AN2P U1487 ( .A(n211), .B(n401), .Z(\ab[5][25] ) );
  AN2P U1488 ( .A(n211), .B(n397), .Z(\ab[5][24] ) );
  AN2P U1489 ( .A(n211), .B(n393), .Z(\ab[5][23] ) );
  AN2P U1490 ( .A(n210), .B(n389), .Z(\ab[5][22] ) );
  AN2P U1491 ( .A(n210), .B(n385), .Z(\ab[5][21] ) );
  AN2P U1492 ( .A(n210), .B(n381), .Z(\ab[5][20] ) );
  AN2P U1493 ( .A(n210), .B(n377), .Z(\ab[5][19] ) );
  AN2P U1494 ( .A(n210), .B(n373), .Z(\ab[5][18] ) );
  AN2P U1495 ( .A(n210), .B(n369), .Z(\ab[5][17] ) );
  AN2P U1496 ( .A(n210), .B(n365), .Z(\ab[5][16] ) );
  AN2P U1497 ( .A(n210), .B(n361), .Z(\ab[5][15] ) );
  AN2P U1498 ( .A(n210), .B(n357), .Z(\ab[5][14] ) );
  AN2P U1499 ( .A(n210), .B(n353), .Z(\ab[5][13] ) );
  AN2P U1500 ( .A(n210), .B(n349), .Z(\ab[5][12] ) );
  AN2P U1501 ( .A(n210), .B(n345), .Z(\ab[5][11] ) );
  AN2P U1502 ( .A(n209), .B(n341), .Z(\ab[5][10] ) );
  AN2P U1503 ( .A(n209), .B(n337), .Z(\ab[5][9] ) );
  AN2P U1504 ( .A(n209), .B(n333), .Z(\ab[5][8] ) );
  AN2P U1505 ( .A(n209), .B(n329), .Z(\ab[5][7] ) );
  AN2P U1506 ( .A(n209), .B(n325), .Z(\ab[5][6] ) );
  AN2P U1507 ( .A(n209), .B(n321), .Z(\ab[5][5] ) );
  AN2P U1508 ( .A(n209), .B(n317), .Z(\ab[5][4] ) );
  AN2P U1509 ( .A(n209), .B(n313), .Z(\ab[5][3] ) );
  AN2P U1510 ( .A(n209), .B(n309), .Z(\ab[5][2] ) );
  AN2P U1511 ( .A(n209), .B(n305), .Z(\ab[5][1] ) );
  AN2P U1512 ( .A(n209), .B(n301), .Z(\ab[5][0] ) );
  AN2P U1513 ( .A(n225), .B(n455), .Z(\ab[6][94] ) );
  AN2P U1514 ( .A(n209), .B(n491), .Z(\ab[5][95] ) );
  AN2P U1515 ( .A(n225), .B(n456), .Z(\ab[6][93] ) );
  AN2P U1516 ( .A(n225), .B(n457), .Z(\ab[6][92] ) );
  AN2P U1517 ( .A(n225), .B(n458), .Z(\ab[6][91] ) );
  AN2P U1518 ( .A(n225), .B(n459), .Z(\ab[6][90] ) );
  AN2P U1519 ( .A(n225), .B(n460), .Z(\ab[6][89] ) );
  AN2P U1520 ( .A(n225), .B(n461), .Z(\ab[6][88] ) );
  AN2P U1521 ( .A(n225), .B(n462), .Z(\ab[6][87] ) );
  AN2P U1522 ( .A(n225), .B(n463), .Z(\ab[6][86] ) );
  AN2P U1523 ( .A(n225), .B(n464), .Z(\ab[6][85] ) );
  AN2P U1524 ( .A(n225), .B(n465), .Z(\ab[6][84] ) );
  AN2P U1525 ( .A(n225), .B(n466), .Z(\ab[6][83] ) );
  AN2P U1526 ( .A(n224), .B(n467), .Z(\ab[6][82] ) );
  AN2P U1527 ( .A(n224), .B(n468), .Z(\ab[6][81] ) );
  AN2P U1528 ( .A(n224), .B(n469), .Z(\ab[6][80] ) );
  AN2P U1529 ( .A(n224), .B(n470), .Z(\ab[6][79] ) );
  AN2P U1530 ( .A(n224), .B(n471), .Z(\ab[6][78] ) );
  AN2P U1531 ( .A(n224), .B(n472), .Z(\ab[6][77] ) );
  AN2P U1532 ( .A(n224), .B(n473), .Z(\ab[6][76] ) );
  AN2P U1533 ( .A(n224), .B(n474), .Z(\ab[6][75] ) );
  AN2P U1534 ( .A(n224), .B(n475), .Z(\ab[6][74] ) );
  AN2P U1535 ( .A(n224), .B(n476), .Z(\ab[6][73] ) );
  AN2P U1536 ( .A(n224), .B(n477), .Z(\ab[6][72] ) );
  AN2P U1537 ( .A(n224), .B(n478), .Z(\ab[6][71] ) );
  AN2P U1538 ( .A(n223), .B(n479), .Z(\ab[6][70] ) );
  AN2P U1539 ( .A(n223), .B(n480), .Z(\ab[6][69] ) );
  AN2P U1540 ( .A(n223), .B(n481), .Z(\ab[6][68] ) );
  AN2P U1541 ( .A(n223), .B(n482), .Z(\ab[6][67] ) );
  AN2P U1542 ( .A(n223), .B(n483), .Z(\ab[6][66] ) );
  AN2P U1543 ( .A(n223), .B(n484), .Z(\ab[6][65] ) );
  AN2P U1544 ( .A(n223), .B(n485), .Z(\ab[6][64] ) );
  AN2P U1545 ( .A(n223), .B(n486), .Z(\ab[6][63] ) );
  AN2P U1546 ( .A(n223), .B(n487), .Z(\ab[6][62] ) );
  AN2P U1547 ( .A(n223), .B(n488), .Z(\ab[6][61] ) );
  AN2P U1548 ( .A(n223), .B(n489), .Z(\ab[6][60] ) );
  AN2P U1549 ( .A(n223), .B(B[59]), .Z(\ab[6][59] ) );
  AN2P U1550 ( .A(n222), .B(B[58]), .Z(\ab[6][58] ) );
  AN2P U1551 ( .A(n222), .B(B[57]), .Z(\ab[6][57] ) );
  AN2P U1552 ( .A(n222), .B(B[56]), .Z(\ab[6][56] ) );
  AN2P U1553 ( .A(n222), .B(n490), .Z(\ab[6][55] ) );
  AN2P U1554 ( .A(n222), .B(B[54]), .Z(\ab[6][54] ) );
  AN2P U1555 ( .A(n222), .B(B[53]), .Z(\ab[6][53] ) );
  AN2P U1556 ( .A(n222), .B(B[52]), .Z(\ab[6][52] ) );
  AN2P U1557 ( .A(n222), .B(B[51]), .Z(\ab[6][51] ) );
  AN2P U1558 ( .A(n222), .B(B[50]), .Z(\ab[6][50] ) );
  AN2P U1559 ( .A(n222), .B(B[49]), .Z(\ab[6][49] ) );
  AN2P U1560 ( .A(n222), .B(B[48]), .Z(\ab[6][48] ) );
  AN2P U1561 ( .A(n222), .B(B[47]), .Z(\ab[6][47] ) );
  AN2P U1562 ( .A(n221), .B(B[46]), .Z(\ab[6][46] ) );
  AN2P U1563 ( .A(n221), .B(B[45]), .Z(\ab[6][45] ) );
  AN2P U1564 ( .A(n221), .B(B[44]), .Z(\ab[6][44] ) );
  AN2P U1565 ( .A(n221), .B(B[43]), .Z(\ab[6][43] ) );
  AN2P U1566 ( .A(n221), .B(B[42]), .Z(\ab[6][42] ) );
  AN2P U1567 ( .A(n221), .B(B[41]), .Z(\ab[6][41] ) );
  AN2P U1568 ( .A(n221), .B(B[40]), .Z(\ab[6][40] ) );
  AN2P U1569 ( .A(n221), .B(B[39]), .Z(\ab[6][39] ) );
  AN2P U1570 ( .A(n221), .B(n452), .Z(\ab[6][38] ) );
  AN2P U1571 ( .A(n221), .B(n448), .Z(\ab[6][37] ) );
  AN2P U1572 ( .A(n221), .B(n444), .Z(\ab[6][36] ) );
  AN2P U1573 ( .A(n221), .B(n440), .Z(\ab[6][35] ) );
  AN2P U1574 ( .A(n220), .B(n436), .Z(\ab[6][34] ) );
  AN2P U1575 ( .A(n220), .B(n432), .Z(\ab[6][33] ) );
  AN2P U1576 ( .A(n220), .B(n428), .Z(\ab[6][32] ) );
  AN2P U1577 ( .A(n220), .B(n424), .Z(\ab[6][31] ) );
  AN2P U1578 ( .A(n220), .B(n420), .Z(\ab[6][30] ) );
  AN2P U1579 ( .A(n220), .B(n416), .Z(\ab[6][29] ) );
  AN2P U1580 ( .A(n220), .B(n412), .Z(\ab[6][28] ) );
  AN2P U1581 ( .A(n220), .B(n408), .Z(\ab[6][27] ) );
  AN2P U1582 ( .A(n220), .B(n404), .Z(\ab[6][26] ) );
  AN2P U1583 ( .A(n220), .B(n400), .Z(\ab[6][25] ) );
  AN2P U1584 ( .A(n220), .B(n396), .Z(\ab[6][24] ) );
  AN2P U1585 ( .A(n220), .B(n392), .Z(\ab[6][23] ) );
  AN2P U1586 ( .A(n219), .B(n388), .Z(\ab[6][22] ) );
  AN2P U1587 ( .A(n219), .B(n384), .Z(\ab[6][21] ) );
  AN2P U1588 ( .A(n219), .B(n380), .Z(\ab[6][20] ) );
  AN2P U1589 ( .A(n219), .B(n376), .Z(\ab[6][19] ) );
  AN2P U1590 ( .A(n219), .B(n372), .Z(\ab[6][18] ) );
  AN2P U1591 ( .A(n219), .B(n368), .Z(\ab[6][17] ) );
  AN2P U1592 ( .A(n219), .B(n364), .Z(\ab[6][16] ) );
  AN2P U1593 ( .A(n219), .B(n360), .Z(\ab[6][15] ) );
  AN2P U1594 ( .A(n219), .B(n356), .Z(\ab[6][14] ) );
  AN2P U1595 ( .A(n219), .B(n352), .Z(\ab[6][13] ) );
  AN2P U1596 ( .A(n219), .B(n348), .Z(\ab[6][12] ) );
  AN2P U1597 ( .A(n219), .B(n344), .Z(\ab[6][11] ) );
  AN2P U1598 ( .A(n218), .B(n340), .Z(\ab[6][10] ) );
  AN2P U1599 ( .A(n218), .B(n336), .Z(\ab[6][9] ) );
  AN2P U1600 ( .A(n218), .B(n332), .Z(\ab[6][8] ) );
  AN2P U1601 ( .A(n218), .B(n328), .Z(\ab[6][7] ) );
  AN2P U1602 ( .A(n218), .B(n324), .Z(\ab[6][6] ) );
  AN2P U1603 ( .A(n218), .B(n320), .Z(\ab[6][5] ) );
  AN2P U1604 ( .A(n218), .B(n316), .Z(\ab[6][4] ) );
  AN2P U1605 ( .A(n218), .B(n312), .Z(\ab[6][3] ) );
  AN2P U1606 ( .A(n218), .B(n308), .Z(\ab[6][2] ) );
  AN2P U1607 ( .A(n218), .B(n304), .Z(\ab[6][1] ) );
  AN2P U1608 ( .A(n218), .B(n300), .Z(\ab[6][0] ) );
  AN2P U1609 ( .A(n234), .B(n455), .Z(\ab[7][94] ) );
  AN2P U1610 ( .A(n218), .B(n491), .Z(\ab[6][95] ) );
  AN2P U1611 ( .A(n234), .B(n456), .Z(\ab[7][93] ) );
  AN2P U1612 ( .A(n234), .B(n457), .Z(\ab[7][92] ) );
  AN2P U1613 ( .A(n234), .B(n458), .Z(\ab[7][91] ) );
  AN2P U1614 ( .A(n234), .B(n459), .Z(\ab[7][90] ) );
  AN2P U1615 ( .A(n234), .B(n460), .Z(\ab[7][89] ) );
  AN2P U1616 ( .A(n234), .B(n461), .Z(\ab[7][88] ) );
  AN2P U1617 ( .A(n234), .B(n462), .Z(\ab[7][87] ) );
  AN2P U1618 ( .A(n234), .B(n463), .Z(\ab[7][86] ) );
  AN2P U1619 ( .A(n234), .B(n464), .Z(\ab[7][85] ) );
  AN2P U1620 ( .A(n234), .B(n465), .Z(\ab[7][84] ) );
  AN2P U1621 ( .A(n234), .B(n466), .Z(\ab[7][83] ) );
  AN2P U1622 ( .A(n233), .B(n467), .Z(\ab[7][82] ) );
  AN2P U1623 ( .A(n233), .B(n468), .Z(\ab[7][81] ) );
  AN2P U1624 ( .A(n233), .B(n469), .Z(\ab[7][80] ) );
  AN2P U1625 ( .A(n233), .B(n470), .Z(\ab[7][79] ) );
  AN2P U1626 ( .A(n233), .B(n471), .Z(\ab[7][78] ) );
  AN2P U1627 ( .A(n233), .B(n472), .Z(\ab[7][77] ) );
  AN2P U1628 ( .A(n233), .B(n473), .Z(\ab[7][76] ) );
  AN2P U1629 ( .A(n233), .B(n474), .Z(\ab[7][75] ) );
  AN2P U1630 ( .A(n233), .B(n475), .Z(\ab[7][74] ) );
  AN2P U1631 ( .A(n233), .B(n476), .Z(\ab[7][73] ) );
  AN2P U1632 ( .A(n233), .B(n477), .Z(\ab[7][72] ) );
  AN2P U1633 ( .A(n233), .B(n478), .Z(\ab[7][71] ) );
  AN2P U1634 ( .A(n232), .B(n479), .Z(\ab[7][70] ) );
  AN2P U1635 ( .A(n232), .B(n480), .Z(\ab[7][69] ) );
  AN2P U1636 ( .A(n232), .B(n481), .Z(\ab[7][68] ) );
  AN2P U1637 ( .A(n232), .B(n482), .Z(\ab[7][67] ) );
  AN2P U1638 ( .A(n232), .B(n483), .Z(\ab[7][66] ) );
  AN2P U1639 ( .A(n232), .B(n484), .Z(\ab[7][65] ) );
  AN2P U1640 ( .A(n232), .B(n485), .Z(\ab[7][64] ) );
  AN2P U1641 ( .A(n232), .B(n486), .Z(\ab[7][63] ) );
  AN2P U1642 ( .A(n232), .B(n487), .Z(\ab[7][62] ) );
  AN2P U1643 ( .A(n232), .B(n488), .Z(\ab[7][61] ) );
  AN2P U1644 ( .A(n232), .B(n489), .Z(\ab[7][60] ) );
  AN2P U1645 ( .A(n232), .B(B[59]), .Z(\ab[7][59] ) );
  AN2P U1646 ( .A(n231), .B(B[58]), .Z(\ab[7][58] ) );
  AN2P U1647 ( .A(n231), .B(B[57]), .Z(\ab[7][57] ) );
  AN2P U1648 ( .A(n231), .B(B[56]), .Z(\ab[7][56] ) );
  AN2P U1649 ( .A(n231), .B(n490), .Z(\ab[7][55] ) );
  AN2P U1650 ( .A(n231), .B(B[54]), .Z(\ab[7][54] ) );
  AN2P U1651 ( .A(n231), .B(B[53]), .Z(\ab[7][53] ) );
  AN2P U1652 ( .A(n231), .B(B[52]), .Z(\ab[7][52] ) );
  AN2P U1653 ( .A(n231), .B(B[51]), .Z(\ab[7][51] ) );
  AN2P U1654 ( .A(n231), .B(B[50]), .Z(\ab[7][50] ) );
  AN2P U1655 ( .A(n231), .B(B[49]), .Z(\ab[7][49] ) );
  AN2P U1656 ( .A(n231), .B(B[48]), .Z(\ab[7][48] ) );
  AN2P U1657 ( .A(n231), .B(B[47]), .Z(\ab[7][47] ) );
  AN2P U1658 ( .A(n230), .B(B[46]), .Z(\ab[7][46] ) );
  AN2P U1659 ( .A(n230), .B(B[45]), .Z(\ab[7][45] ) );
  AN2P U1660 ( .A(n230), .B(B[44]), .Z(\ab[7][44] ) );
  AN2P U1661 ( .A(n230), .B(B[43]), .Z(\ab[7][43] ) );
  AN2P U1662 ( .A(n230), .B(B[42]), .Z(\ab[7][42] ) );
  AN2P U1663 ( .A(n230), .B(B[41]), .Z(\ab[7][41] ) );
  AN2P U1664 ( .A(n230), .B(B[40]), .Z(\ab[7][40] ) );
  AN2P U1665 ( .A(n230), .B(B[39]), .Z(\ab[7][39] ) );
  AN2P U1666 ( .A(n230), .B(n452), .Z(\ab[7][38] ) );
  AN2P U1667 ( .A(n230), .B(n448), .Z(\ab[7][37] ) );
  AN2P U1668 ( .A(n230), .B(n444), .Z(\ab[7][36] ) );
  AN2P U1669 ( .A(n230), .B(n440), .Z(\ab[7][35] ) );
  AN2P U1670 ( .A(n229), .B(n436), .Z(\ab[7][34] ) );
  AN2P U1671 ( .A(n229), .B(n432), .Z(\ab[7][33] ) );
  AN2P U1672 ( .A(n229), .B(n428), .Z(\ab[7][32] ) );
  AN2P U1673 ( .A(n229), .B(n424), .Z(\ab[7][31] ) );
  AN2P U1674 ( .A(n229), .B(n420), .Z(\ab[7][30] ) );
  AN2P U1675 ( .A(n229), .B(n416), .Z(\ab[7][29] ) );
  AN2P U1676 ( .A(n229), .B(n412), .Z(\ab[7][28] ) );
  AN2P U1677 ( .A(n229), .B(n408), .Z(\ab[7][27] ) );
  AN2P U1678 ( .A(n229), .B(n404), .Z(\ab[7][26] ) );
  AN2P U1679 ( .A(n229), .B(n400), .Z(\ab[7][25] ) );
  AN2P U1680 ( .A(n229), .B(n396), .Z(\ab[7][24] ) );
  AN2P U1681 ( .A(n229), .B(n392), .Z(\ab[7][23] ) );
  AN2P U1682 ( .A(n228), .B(n388), .Z(\ab[7][22] ) );
  AN2P U1683 ( .A(n228), .B(n384), .Z(\ab[7][21] ) );
  AN2P U1684 ( .A(n228), .B(n380), .Z(\ab[7][20] ) );
  AN2P U1685 ( .A(n228), .B(n376), .Z(\ab[7][19] ) );
  AN2P U1686 ( .A(n228), .B(n372), .Z(\ab[7][18] ) );
  AN2P U1687 ( .A(n228), .B(n368), .Z(\ab[7][17] ) );
  AN2P U1688 ( .A(n228), .B(n364), .Z(\ab[7][16] ) );
  AN2P U1689 ( .A(n228), .B(n360), .Z(\ab[7][15] ) );
  AN2P U1690 ( .A(n228), .B(n356), .Z(\ab[7][14] ) );
  AN2P U1691 ( .A(n228), .B(n352), .Z(\ab[7][13] ) );
  AN2P U1692 ( .A(n228), .B(n348), .Z(\ab[7][12] ) );
  AN2P U1693 ( .A(n228), .B(n344), .Z(\ab[7][11] ) );
  AN2P U1694 ( .A(n227), .B(n340), .Z(\ab[7][10] ) );
  AN2P U1695 ( .A(n227), .B(n336), .Z(\ab[7][9] ) );
  AN2P U1696 ( .A(n227), .B(n332), .Z(\ab[7][8] ) );
  AN2P U1697 ( .A(n227), .B(n328), .Z(\ab[7][7] ) );
  AN2P U1698 ( .A(n227), .B(n324), .Z(\ab[7][6] ) );
  AN2P U1699 ( .A(n227), .B(n320), .Z(\ab[7][5] ) );
  AN2P U1700 ( .A(n227), .B(n316), .Z(\ab[7][4] ) );
  AN2P U1701 ( .A(n227), .B(n312), .Z(\ab[7][3] ) );
  AN2P U1702 ( .A(n227), .B(n308), .Z(\ab[7][2] ) );
  AN2P U1703 ( .A(n227), .B(n304), .Z(\ab[7][1] ) );
  AN2P U1704 ( .A(n227), .B(n300), .Z(\ab[7][0] ) );
  AN2P U1705 ( .A(n243), .B(n455), .Z(\ab[8][94] ) );
  AN2P U1706 ( .A(n227), .B(n491), .Z(\ab[7][95] ) );
  AN2P U1707 ( .A(n243), .B(n456), .Z(\ab[8][93] ) );
  AN2P U1708 ( .A(n243), .B(n457), .Z(\ab[8][92] ) );
  AN2P U1709 ( .A(n243), .B(n458), .Z(\ab[8][91] ) );
  AN2P U1710 ( .A(n243), .B(n459), .Z(\ab[8][90] ) );
  AN2P U1711 ( .A(n243), .B(n460), .Z(\ab[8][89] ) );
  AN2P U1712 ( .A(n243), .B(n461), .Z(\ab[8][88] ) );
  AN2P U1713 ( .A(n243), .B(n462), .Z(\ab[8][87] ) );
  AN2P U1714 ( .A(n243), .B(n463), .Z(\ab[8][86] ) );
  AN2P U1715 ( .A(n243), .B(n464), .Z(\ab[8][85] ) );
  AN2P U1716 ( .A(n243), .B(n465), .Z(\ab[8][84] ) );
  AN2P U1717 ( .A(n243), .B(n466), .Z(\ab[8][83] ) );
  AN2P U1718 ( .A(n242), .B(n467), .Z(\ab[8][82] ) );
  AN2P U1719 ( .A(n242), .B(n468), .Z(\ab[8][81] ) );
  AN2P U1720 ( .A(n242), .B(n469), .Z(\ab[8][80] ) );
  AN2P U1721 ( .A(n242), .B(n470), .Z(\ab[8][79] ) );
  AN2P U1722 ( .A(n242), .B(n471), .Z(\ab[8][78] ) );
  AN2P U1723 ( .A(n242), .B(n472), .Z(\ab[8][77] ) );
  AN2P U1724 ( .A(n242), .B(n473), .Z(\ab[8][76] ) );
  AN2P U1725 ( .A(n242), .B(n474), .Z(\ab[8][75] ) );
  AN2P U1726 ( .A(n242), .B(n475), .Z(\ab[8][74] ) );
  AN2P U1727 ( .A(n242), .B(n476), .Z(\ab[8][73] ) );
  AN2P U1728 ( .A(n242), .B(n477), .Z(\ab[8][72] ) );
  AN2P U1729 ( .A(n242), .B(n478), .Z(\ab[8][71] ) );
  AN2P U1730 ( .A(n241), .B(n479), .Z(\ab[8][70] ) );
  AN2P U1731 ( .A(n241), .B(n480), .Z(\ab[8][69] ) );
  AN2P U1732 ( .A(n241), .B(n481), .Z(\ab[8][68] ) );
  AN2P U1733 ( .A(n241), .B(n482), .Z(\ab[8][67] ) );
  AN2P U1734 ( .A(n241), .B(n483), .Z(\ab[8][66] ) );
  AN2P U1735 ( .A(n241), .B(n484), .Z(\ab[8][65] ) );
  AN2P U1736 ( .A(n241), .B(n485), .Z(\ab[8][64] ) );
  AN2P U1737 ( .A(n241), .B(n486), .Z(\ab[8][63] ) );
  AN2P U1738 ( .A(n241), .B(n487), .Z(\ab[8][62] ) );
  AN2P U1739 ( .A(n241), .B(n488), .Z(\ab[8][61] ) );
  AN2P U1740 ( .A(n241), .B(n489), .Z(\ab[8][60] ) );
  AN2P U1741 ( .A(n241), .B(B[59]), .Z(\ab[8][59] ) );
  AN2P U1742 ( .A(n240), .B(B[58]), .Z(\ab[8][58] ) );
  AN2P U1743 ( .A(n240), .B(B[57]), .Z(\ab[8][57] ) );
  AN2P U1744 ( .A(n240), .B(B[56]), .Z(\ab[8][56] ) );
  AN2P U1745 ( .A(n240), .B(n490), .Z(\ab[8][55] ) );
  AN2P U1746 ( .A(n240), .B(B[54]), .Z(\ab[8][54] ) );
  AN2P U1747 ( .A(n240), .B(B[53]), .Z(\ab[8][53] ) );
  AN2P U1748 ( .A(n240), .B(B[52]), .Z(\ab[8][52] ) );
  AN2P U1749 ( .A(n240), .B(B[51]), .Z(\ab[8][51] ) );
  AN2P U1750 ( .A(n240), .B(B[50]), .Z(\ab[8][50] ) );
  AN2P U1751 ( .A(n240), .B(B[49]), .Z(\ab[8][49] ) );
  AN2P U1752 ( .A(n240), .B(B[48]), .Z(\ab[8][48] ) );
  AN2P U1753 ( .A(n240), .B(B[47]), .Z(\ab[8][47] ) );
  AN2P U1754 ( .A(n239), .B(B[46]), .Z(\ab[8][46] ) );
  AN2P U1755 ( .A(n239), .B(B[45]), .Z(\ab[8][45] ) );
  AN2P U1756 ( .A(n239), .B(B[44]), .Z(\ab[8][44] ) );
  AN2P U1757 ( .A(n239), .B(B[43]), .Z(\ab[8][43] ) );
  AN2P U1758 ( .A(n239), .B(B[42]), .Z(\ab[8][42] ) );
  AN2P U1759 ( .A(n239), .B(B[41]), .Z(\ab[8][41] ) );
  AN2P U1760 ( .A(n239), .B(B[40]), .Z(\ab[8][40] ) );
  AN2P U1761 ( .A(n239), .B(B[39]), .Z(\ab[8][39] ) );
  AN2P U1762 ( .A(n239), .B(n452), .Z(\ab[8][38] ) );
  AN2P U1763 ( .A(n239), .B(n448), .Z(\ab[8][37] ) );
  AN2P U1764 ( .A(n239), .B(n444), .Z(\ab[8][36] ) );
  AN2P U1765 ( .A(n239), .B(n440), .Z(\ab[8][35] ) );
  AN2P U1766 ( .A(n238), .B(n436), .Z(\ab[8][34] ) );
  AN2P U1767 ( .A(n238), .B(n432), .Z(\ab[8][33] ) );
  AN2P U1768 ( .A(n238), .B(n428), .Z(\ab[8][32] ) );
  AN2P U1769 ( .A(n238), .B(n424), .Z(\ab[8][31] ) );
  AN2P U1770 ( .A(n238), .B(n420), .Z(\ab[8][30] ) );
  AN2P U1771 ( .A(n238), .B(n416), .Z(\ab[8][29] ) );
  AN2P U1772 ( .A(n238), .B(n412), .Z(\ab[8][28] ) );
  AN2P U1773 ( .A(n238), .B(n408), .Z(\ab[8][27] ) );
  AN2P U1774 ( .A(n238), .B(n404), .Z(\ab[8][26] ) );
  AN2P U1775 ( .A(n238), .B(n400), .Z(\ab[8][25] ) );
  AN2P U1776 ( .A(n238), .B(n396), .Z(\ab[8][24] ) );
  AN2P U1777 ( .A(n238), .B(n392), .Z(\ab[8][23] ) );
  AN2P U1778 ( .A(n237), .B(n388), .Z(\ab[8][22] ) );
  AN2P U1779 ( .A(n237), .B(n384), .Z(\ab[8][21] ) );
  AN2P U1780 ( .A(n237), .B(n380), .Z(\ab[8][20] ) );
  AN2P U1781 ( .A(n237), .B(n376), .Z(\ab[8][19] ) );
  AN2P U1782 ( .A(n237), .B(n372), .Z(\ab[8][18] ) );
  AN2P U1783 ( .A(n237), .B(n368), .Z(\ab[8][17] ) );
  AN2P U1784 ( .A(n237), .B(n364), .Z(\ab[8][16] ) );
  AN2P U1785 ( .A(n237), .B(n360), .Z(\ab[8][15] ) );
  AN2P U1786 ( .A(n237), .B(n356), .Z(\ab[8][14] ) );
  AN2P U1787 ( .A(n237), .B(n352), .Z(\ab[8][13] ) );
  AN2P U1788 ( .A(n237), .B(n348), .Z(\ab[8][12] ) );
  AN2P U1789 ( .A(n237), .B(n344), .Z(\ab[8][11] ) );
  AN2P U1790 ( .A(n236), .B(n340), .Z(\ab[8][10] ) );
  AN2P U1791 ( .A(n236), .B(n336), .Z(\ab[8][9] ) );
  AN2P U1792 ( .A(n236), .B(n332), .Z(\ab[8][8] ) );
  AN2P U1793 ( .A(n236), .B(n328), .Z(\ab[8][7] ) );
  AN2P U1794 ( .A(n236), .B(n324), .Z(\ab[8][6] ) );
  AN2P U1795 ( .A(n236), .B(n320), .Z(\ab[8][5] ) );
  AN2P U1796 ( .A(n236), .B(n316), .Z(\ab[8][4] ) );
  AN2P U1797 ( .A(n236), .B(n312), .Z(\ab[8][3] ) );
  AN2P U1798 ( .A(n236), .B(n308), .Z(\ab[8][2] ) );
  AN2P U1799 ( .A(n236), .B(n304), .Z(\ab[8][1] ) );
  AN2P U1800 ( .A(n236), .B(n300), .Z(\ab[8][0] ) );
  AN2P U1801 ( .A(n252), .B(n455), .Z(\ab[9][94] ) );
  AN2P U1802 ( .A(n236), .B(n491), .Z(\ab[8][95] ) );
  AN2P U1803 ( .A(n252), .B(n456), .Z(\ab[9][93] ) );
  AN2P U1804 ( .A(n252), .B(n457), .Z(\ab[9][92] ) );
  AN2P U1805 ( .A(n252), .B(n458), .Z(\ab[9][91] ) );
  AN2P U1806 ( .A(n252), .B(n459), .Z(\ab[9][90] ) );
  AN2P U1807 ( .A(n252), .B(n460), .Z(\ab[9][89] ) );
  AN2P U1808 ( .A(n252), .B(n461), .Z(\ab[9][88] ) );
  AN2P U1809 ( .A(n252), .B(n462), .Z(\ab[9][87] ) );
  AN2P U1810 ( .A(n252), .B(n463), .Z(\ab[9][86] ) );
  AN2P U1811 ( .A(n252), .B(n464), .Z(\ab[9][85] ) );
  AN2P U1812 ( .A(n252), .B(n465), .Z(\ab[9][84] ) );
  AN2P U1813 ( .A(n252), .B(n466), .Z(\ab[9][83] ) );
  AN2P U1814 ( .A(n251), .B(n467), .Z(\ab[9][82] ) );
  AN2P U1815 ( .A(n251), .B(n468), .Z(\ab[9][81] ) );
  AN2P U1816 ( .A(n251), .B(n469), .Z(\ab[9][80] ) );
  AN2P U1817 ( .A(n251), .B(n470), .Z(\ab[9][79] ) );
  AN2P U1818 ( .A(n251), .B(n471), .Z(\ab[9][78] ) );
  AN2P U1819 ( .A(n251), .B(n472), .Z(\ab[9][77] ) );
  AN2P U1820 ( .A(n251), .B(n473), .Z(\ab[9][76] ) );
  AN2P U1821 ( .A(n251), .B(n474), .Z(\ab[9][75] ) );
  AN2P U1822 ( .A(n251), .B(n475), .Z(\ab[9][74] ) );
  AN2P U1823 ( .A(n251), .B(n476), .Z(\ab[9][73] ) );
  AN2P U1824 ( .A(n251), .B(n477), .Z(\ab[9][72] ) );
  AN2P U1825 ( .A(n251), .B(n478), .Z(\ab[9][71] ) );
  AN2P U1826 ( .A(n250), .B(n479), .Z(\ab[9][70] ) );
  AN2P U1827 ( .A(n250), .B(n480), .Z(\ab[9][69] ) );
  AN2P U1828 ( .A(n250), .B(n481), .Z(\ab[9][68] ) );
  AN2P U1829 ( .A(n250), .B(n482), .Z(\ab[9][67] ) );
  AN2P U1830 ( .A(n250), .B(n483), .Z(\ab[9][66] ) );
  AN2P U1831 ( .A(n250), .B(n484), .Z(\ab[9][65] ) );
  AN2P U1832 ( .A(n250), .B(n485), .Z(\ab[9][64] ) );
  AN2P U1833 ( .A(n250), .B(n486), .Z(\ab[9][63] ) );
  AN2P U1834 ( .A(n250), .B(n487), .Z(\ab[9][62] ) );
  AN2P U1835 ( .A(n250), .B(n488), .Z(\ab[9][61] ) );
  AN2P U1836 ( .A(n250), .B(n489), .Z(\ab[9][60] ) );
  AN2P U1837 ( .A(n250), .B(B[59]), .Z(\ab[9][59] ) );
  AN2P U1838 ( .A(n249), .B(B[58]), .Z(\ab[9][58] ) );
  AN2P U1839 ( .A(n249), .B(B[57]), .Z(\ab[9][57] ) );
  AN2P U1840 ( .A(n249), .B(B[56]), .Z(\ab[9][56] ) );
  AN2P U1841 ( .A(n249), .B(n490), .Z(\ab[9][55] ) );
  AN2P U1842 ( .A(n249), .B(B[54]), .Z(\ab[9][54] ) );
  AN2P U1843 ( .A(n249), .B(B[53]), .Z(\ab[9][53] ) );
  AN2P U1844 ( .A(n249), .B(B[52]), .Z(\ab[9][52] ) );
  AN2P U1845 ( .A(n249), .B(B[51]), .Z(\ab[9][51] ) );
  AN2P U1846 ( .A(n249), .B(B[50]), .Z(\ab[9][50] ) );
  AN2P U1847 ( .A(n249), .B(B[49]), .Z(\ab[9][49] ) );
  AN2P U1848 ( .A(n249), .B(B[48]), .Z(\ab[9][48] ) );
  AN2P U1849 ( .A(n249), .B(B[47]), .Z(\ab[9][47] ) );
  AN2P U1850 ( .A(n248), .B(B[46]), .Z(\ab[9][46] ) );
  AN2P U1851 ( .A(n248), .B(B[45]), .Z(\ab[9][45] ) );
  AN2P U1852 ( .A(n248), .B(B[44]), .Z(\ab[9][44] ) );
  AN2P U1853 ( .A(n248), .B(B[43]), .Z(\ab[9][43] ) );
  AN2P U1854 ( .A(n248), .B(B[42]), .Z(\ab[9][42] ) );
  AN2P U1855 ( .A(n248), .B(B[41]), .Z(\ab[9][41] ) );
  AN2P U1856 ( .A(n248), .B(B[40]), .Z(\ab[9][40] ) );
  AN2P U1857 ( .A(n248), .B(B[39]), .Z(\ab[9][39] ) );
  AN2P U1858 ( .A(n248), .B(n452), .Z(\ab[9][38] ) );
  AN2P U1859 ( .A(n248), .B(n448), .Z(\ab[9][37] ) );
  AN2P U1860 ( .A(n248), .B(n444), .Z(\ab[9][36] ) );
  AN2P U1861 ( .A(n248), .B(n440), .Z(\ab[9][35] ) );
  AN2P U1862 ( .A(n247), .B(n436), .Z(\ab[9][34] ) );
  AN2P U1863 ( .A(n247), .B(n432), .Z(\ab[9][33] ) );
  AN2P U1864 ( .A(n247), .B(n428), .Z(\ab[9][32] ) );
  AN2P U1865 ( .A(n247), .B(n424), .Z(\ab[9][31] ) );
  AN2P U1866 ( .A(n247), .B(n420), .Z(\ab[9][30] ) );
  AN2P U1867 ( .A(n247), .B(n416), .Z(\ab[9][29] ) );
  AN2P U1868 ( .A(n247), .B(n412), .Z(\ab[9][28] ) );
  AN2P U1869 ( .A(n247), .B(n408), .Z(\ab[9][27] ) );
  AN2P U1870 ( .A(n247), .B(n404), .Z(\ab[9][26] ) );
  AN2P U1871 ( .A(n247), .B(n400), .Z(\ab[9][25] ) );
  AN2P U1872 ( .A(n247), .B(n396), .Z(\ab[9][24] ) );
  AN2P U1873 ( .A(n247), .B(n392), .Z(\ab[9][23] ) );
  AN2P U1874 ( .A(n246), .B(n388), .Z(\ab[9][22] ) );
  AN2P U1875 ( .A(n246), .B(n384), .Z(\ab[9][21] ) );
  AN2P U1876 ( .A(n246), .B(n380), .Z(\ab[9][20] ) );
  AN2P U1877 ( .A(n246), .B(n376), .Z(\ab[9][19] ) );
  AN2P U1878 ( .A(n246), .B(n372), .Z(\ab[9][18] ) );
  AN2P U1879 ( .A(n246), .B(n368), .Z(\ab[9][17] ) );
  AN2P U1880 ( .A(n246), .B(n364), .Z(\ab[9][16] ) );
  AN2P U1881 ( .A(n246), .B(n360), .Z(\ab[9][15] ) );
  AN2P U1882 ( .A(n246), .B(n356), .Z(\ab[9][14] ) );
  AN2P U1883 ( .A(n246), .B(n352), .Z(\ab[9][13] ) );
  AN2P U1884 ( .A(n246), .B(n348), .Z(\ab[9][12] ) );
  AN2P U1885 ( .A(n246), .B(n344), .Z(\ab[9][11] ) );
  AN2P U1886 ( .A(n245), .B(n340), .Z(\ab[9][10] ) );
  AN2P U1887 ( .A(n245), .B(n336), .Z(\ab[9][9] ) );
  AN2P U1888 ( .A(n245), .B(n332), .Z(\ab[9][8] ) );
  AN2P U1889 ( .A(n245), .B(n328), .Z(\ab[9][7] ) );
  AN2P U1890 ( .A(n245), .B(n324), .Z(\ab[9][6] ) );
  AN2P U1891 ( .A(n245), .B(n320), .Z(\ab[9][5] ) );
  AN2P U1892 ( .A(n245), .B(n316), .Z(\ab[9][4] ) );
  AN2P U1893 ( .A(n245), .B(n312), .Z(\ab[9][3] ) );
  AN2P U1894 ( .A(n245), .B(n308), .Z(\ab[9][2] ) );
  AN2P U1895 ( .A(n245), .B(n304), .Z(\ab[9][1] ) );
  AN2P U1896 ( .A(n245), .B(n300), .Z(\ab[9][0] ) );
  AN2P U1897 ( .A(n261), .B(n455), .Z(\ab[10][94] ) );
  AN2P U1898 ( .A(n245), .B(n491), .Z(\ab[9][95] ) );
  AN2P U1899 ( .A(n261), .B(n456), .Z(\ab[10][93] ) );
  AN2P U1900 ( .A(n261), .B(n457), .Z(\ab[10][92] ) );
  AN2P U1901 ( .A(n261), .B(n458), .Z(\ab[10][91] ) );
  AN2P U1902 ( .A(n261), .B(n459), .Z(\ab[10][90] ) );
  AN2P U1903 ( .A(n261), .B(n460), .Z(\ab[10][89] ) );
  AN2P U1904 ( .A(n261), .B(n461), .Z(\ab[10][88] ) );
  AN2P U1905 ( .A(n261), .B(n462), .Z(\ab[10][87] ) );
  AN2P U1906 ( .A(n261), .B(n463), .Z(\ab[10][86] ) );
  AN2P U1907 ( .A(n261), .B(n464), .Z(\ab[10][85] ) );
  AN2P U1908 ( .A(n261), .B(n465), .Z(\ab[10][84] ) );
  AN2P U1909 ( .A(n261), .B(n466), .Z(\ab[10][83] ) );
  AN2P U1910 ( .A(n260), .B(n467), .Z(\ab[10][82] ) );
  AN2P U1911 ( .A(n260), .B(n468), .Z(\ab[10][81] ) );
  AN2P U1912 ( .A(n260), .B(n469), .Z(\ab[10][80] ) );
  AN2P U1913 ( .A(n260), .B(n470), .Z(\ab[10][79] ) );
  AN2P U1914 ( .A(n260), .B(n471), .Z(\ab[10][78] ) );
  AN2P U1915 ( .A(n260), .B(n472), .Z(\ab[10][77] ) );
  AN2P U1916 ( .A(n260), .B(n473), .Z(\ab[10][76] ) );
  AN2P U1917 ( .A(n260), .B(n474), .Z(\ab[10][75] ) );
  AN2P U1918 ( .A(n260), .B(n475), .Z(\ab[10][74] ) );
  AN2P U1919 ( .A(n260), .B(n476), .Z(\ab[10][73] ) );
  AN2P U1920 ( .A(n260), .B(n477), .Z(\ab[10][72] ) );
  AN2P U1921 ( .A(n260), .B(n478), .Z(\ab[10][71] ) );
  AN2P U1922 ( .A(n259), .B(n479), .Z(\ab[10][70] ) );
  AN2P U1923 ( .A(n259), .B(n480), .Z(\ab[10][69] ) );
  AN2P U1924 ( .A(n259), .B(n481), .Z(\ab[10][68] ) );
  AN2P U1925 ( .A(n259), .B(n482), .Z(\ab[10][67] ) );
  AN2P U1926 ( .A(n259), .B(n483), .Z(\ab[10][66] ) );
  AN2P U1927 ( .A(n259), .B(n484), .Z(\ab[10][65] ) );
  AN2P U1928 ( .A(n259), .B(n485), .Z(\ab[10][64] ) );
  AN2P U1929 ( .A(n259), .B(n486), .Z(\ab[10][63] ) );
  AN2P U1930 ( .A(n259), .B(n487), .Z(\ab[10][62] ) );
  AN2P U1931 ( .A(n259), .B(n488), .Z(\ab[10][61] ) );
  AN2P U1932 ( .A(n259), .B(n489), .Z(\ab[10][60] ) );
  AN2P U1933 ( .A(n259), .B(B[59]), .Z(\ab[10][59] ) );
  AN2P U1934 ( .A(n258), .B(B[58]), .Z(\ab[10][58] ) );
  AN2P U1935 ( .A(n258), .B(B[57]), .Z(\ab[10][57] ) );
  AN2P U1936 ( .A(n258), .B(B[56]), .Z(\ab[10][56] ) );
  AN2P U1937 ( .A(n258), .B(n490), .Z(\ab[10][55] ) );
  AN2P U1938 ( .A(n258), .B(B[54]), .Z(\ab[10][54] ) );
  AN2P U1939 ( .A(n258), .B(B[53]), .Z(\ab[10][53] ) );
  AN2P U1940 ( .A(n258), .B(B[52]), .Z(\ab[10][52] ) );
  AN2P U1941 ( .A(n258), .B(B[51]), .Z(\ab[10][51] ) );
  AN2P U1942 ( .A(n258), .B(B[50]), .Z(\ab[10][50] ) );
  AN2P U1943 ( .A(n258), .B(B[49]), .Z(\ab[10][49] ) );
  AN2P U1944 ( .A(n258), .B(B[48]), .Z(\ab[10][48] ) );
  AN2P U1945 ( .A(n258), .B(B[47]), .Z(\ab[10][47] ) );
  AN2P U1946 ( .A(n257), .B(B[46]), .Z(\ab[10][46] ) );
  AN2P U1947 ( .A(n257), .B(B[45]), .Z(\ab[10][45] ) );
  AN2P U1948 ( .A(n257), .B(B[44]), .Z(\ab[10][44] ) );
  AN2P U1949 ( .A(n257), .B(B[43]), .Z(\ab[10][43] ) );
  AN2P U1950 ( .A(n257), .B(B[42]), .Z(\ab[10][42] ) );
  AN2P U1951 ( .A(n257), .B(B[41]), .Z(\ab[10][41] ) );
  AN2P U1952 ( .A(n257), .B(B[40]), .Z(\ab[10][40] ) );
  AN2P U1953 ( .A(n257), .B(B[39]), .Z(\ab[10][39] ) );
  AN2P U1954 ( .A(n257), .B(n452), .Z(\ab[10][38] ) );
  AN2P U1955 ( .A(n257), .B(n448), .Z(\ab[10][37] ) );
  AN2P U1956 ( .A(n257), .B(n444), .Z(\ab[10][36] ) );
  AN2P U1957 ( .A(n257), .B(n440), .Z(\ab[10][35] ) );
  AN2P U1958 ( .A(n256), .B(n436), .Z(\ab[10][34] ) );
  AN2P U1959 ( .A(n256), .B(n432), .Z(\ab[10][33] ) );
  AN2P U1960 ( .A(n256), .B(n428), .Z(\ab[10][32] ) );
  AN2P U1961 ( .A(n256), .B(n424), .Z(\ab[10][31] ) );
  AN2P U1962 ( .A(n256), .B(n420), .Z(\ab[10][30] ) );
  AN2P U1963 ( .A(n256), .B(n416), .Z(\ab[10][29] ) );
  AN2P U1964 ( .A(n256), .B(n412), .Z(\ab[10][28] ) );
  AN2P U1965 ( .A(n256), .B(n408), .Z(\ab[10][27] ) );
  AN2P U1966 ( .A(n256), .B(n404), .Z(\ab[10][26] ) );
  AN2P U1967 ( .A(n256), .B(n400), .Z(\ab[10][25] ) );
  AN2P U1968 ( .A(n256), .B(n396), .Z(\ab[10][24] ) );
  AN2P U1969 ( .A(n256), .B(n392), .Z(\ab[10][23] ) );
  AN2P U1970 ( .A(n255), .B(n388), .Z(\ab[10][22] ) );
  AN2P U1971 ( .A(n255), .B(n384), .Z(\ab[10][21] ) );
  AN2P U1972 ( .A(n255), .B(n380), .Z(\ab[10][20] ) );
  AN2P U1973 ( .A(n255), .B(n376), .Z(\ab[10][19] ) );
  AN2P U1974 ( .A(n255), .B(n372), .Z(\ab[10][18] ) );
  AN2P U1975 ( .A(n255), .B(n368), .Z(\ab[10][17] ) );
  AN2P U1976 ( .A(n255), .B(n364), .Z(\ab[10][16] ) );
  AN2P U1977 ( .A(n255), .B(n360), .Z(\ab[10][15] ) );
  AN2P U1978 ( .A(n255), .B(n356), .Z(\ab[10][14] ) );
  AN2P U1979 ( .A(n255), .B(n352), .Z(\ab[10][13] ) );
  AN2P U1980 ( .A(n255), .B(n348), .Z(\ab[10][12] ) );
  AN2P U1981 ( .A(n255), .B(n344), .Z(\ab[10][11] ) );
  AN2P U1982 ( .A(n254), .B(n340), .Z(\ab[10][10] ) );
  AN2P U1983 ( .A(n254), .B(n336), .Z(\ab[10][9] ) );
  AN2P U1984 ( .A(n254), .B(n332), .Z(\ab[10][8] ) );
  AN2P U1985 ( .A(n254), .B(n328), .Z(\ab[10][7] ) );
  AN2P U1986 ( .A(n254), .B(n324), .Z(\ab[10][6] ) );
  AN2P U1987 ( .A(n254), .B(n320), .Z(\ab[10][5] ) );
  AN2P U1988 ( .A(n254), .B(n316), .Z(\ab[10][4] ) );
  AN2P U1989 ( .A(n254), .B(n312), .Z(\ab[10][3] ) );
  AN2P U1990 ( .A(n254), .B(n308), .Z(\ab[10][2] ) );
  AN2P U1991 ( .A(n254), .B(n304), .Z(\ab[10][1] ) );
  AN2P U1992 ( .A(n254), .B(n300), .Z(\ab[10][0] ) );
  AN2P U1993 ( .A(n270), .B(n455), .Z(\ab[11][94] ) );
  AN2P U1994 ( .A(n254), .B(n491), .Z(\ab[10][95] ) );
  AN2P U1995 ( .A(n270), .B(n456), .Z(\ab[11][93] ) );
  AN2P U1996 ( .A(n270), .B(n457), .Z(\ab[11][92] ) );
  AN2P U1997 ( .A(n270), .B(n458), .Z(\ab[11][91] ) );
  AN2P U1998 ( .A(n270), .B(n459), .Z(\ab[11][90] ) );
  AN2P U1999 ( .A(n270), .B(n460), .Z(\ab[11][89] ) );
  AN2P U2000 ( .A(n270), .B(n461), .Z(\ab[11][88] ) );
  AN2P U2001 ( .A(n270), .B(n462), .Z(\ab[11][87] ) );
  AN2P U2002 ( .A(n270), .B(n463), .Z(\ab[11][86] ) );
  AN2P U2003 ( .A(n270), .B(n464), .Z(\ab[11][85] ) );
  AN2P U2004 ( .A(n270), .B(n465), .Z(\ab[11][84] ) );
  AN2P U2005 ( .A(n270), .B(n466), .Z(\ab[11][83] ) );
  AN2P U2006 ( .A(n269), .B(n467), .Z(\ab[11][82] ) );
  AN2P U2007 ( .A(n269), .B(n468), .Z(\ab[11][81] ) );
  AN2P U2008 ( .A(n269), .B(n469), .Z(\ab[11][80] ) );
  AN2P U2009 ( .A(n269), .B(n470), .Z(\ab[11][79] ) );
  AN2P U2010 ( .A(n269), .B(n471), .Z(\ab[11][78] ) );
  AN2P U2011 ( .A(n269), .B(n472), .Z(\ab[11][77] ) );
  AN2P U2012 ( .A(n269), .B(n473), .Z(\ab[11][76] ) );
  AN2P U2013 ( .A(n269), .B(n474), .Z(\ab[11][75] ) );
  AN2P U2014 ( .A(n269), .B(n475), .Z(\ab[11][74] ) );
  AN2P U2015 ( .A(n269), .B(n476), .Z(\ab[11][73] ) );
  AN2P U2016 ( .A(n269), .B(n477), .Z(\ab[11][72] ) );
  AN2P U2017 ( .A(n269), .B(n478), .Z(\ab[11][71] ) );
  AN2P U2018 ( .A(n268), .B(n479), .Z(\ab[11][70] ) );
  AN2P U2019 ( .A(n268), .B(n480), .Z(\ab[11][69] ) );
  AN2P U2020 ( .A(n268), .B(n481), .Z(\ab[11][68] ) );
  AN2P U2021 ( .A(n268), .B(n482), .Z(\ab[11][67] ) );
  AN2P U2022 ( .A(n268), .B(n483), .Z(\ab[11][66] ) );
  AN2P U2023 ( .A(n268), .B(n484), .Z(\ab[11][65] ) );
  AN2P U2024 ( .A(n268), .B(n485), .Z(\ab[11][64] ) );
  AN2P U2025 ( .A(n268), .B(n486), .Z(\ab[11][63] ) );
  AN2P U2026 ( .A(n268), .B(n487), .Z(\ab[11][62] ) );
  AN2P U2027 ( .A(n268), .B(n488), .Z(\ab[11][61] ) );
  AN2P U2028 ( .A(n268), .B(n489), .Z(\ab[11][60] ) );
  AN2P U2029 ( .A(n268), .B(B[59]), .Z(\ab[11][59] ) );
  AN2P U2030 ( .A(n267), .B(B[58]), .Z(\ab[11][58] ) );
  AN2P U2031 ( .A(n267), .B(B[57]), .Z(\ab[11][57] ) );
  AN2P U2032 ( .A(n267), .B(B[56]), .Z(\ab[11][56] ) );
  AN2P U2033 ( .A(n267), .B(n490), .Z(\ab[11][55] ) );
  AN2P U2034 ( .A(n267), .B(B[54]), .Z(\ab[11][54] ) );
  AN2P U2035 ( .A(n267), .B(B[53]), .Z(\ab[11][53] ) );
  AN2P U2036 ( .A(n267), .B(B[52]), .Z(\ab[11][52] ) );
  AN2P U2037 ( .A(n267), .B(B[51]), .Z(\ab[11][51] ) );
  AN2P U2038 ( .A(n267), .B(B[50]), .Z(\ab[11][50] ) );
  AN2P U2039 ( .A(n267), .B(B[49]), .Z(\ab[11][49] ) );
  AN2P U2040 ( .A(n267), .B(B[48]), .Z(\ab[11][48] ) );
  AN2P U2041 ( .A(n267), .B(B[47]), .Z(\ab[11][47] ) );
  AN2P U2042 ( .A(n266), .B(B[46]), .Z(\ab[11][46] ) );
  AN2P U2043 ( .A(n266), .B(B[45]), .Z(\ab[11][45] ) );
  AN2P U2044 ( .A(n266), .B(B[44]), .Z(\ab[11][44] ) );
  AN2P U2045 ( .A(n266), .B(B[43]), .Z(\ab[11][43] ) );
  AN2P U2046 ( .A(n266), .B(B[42]), .Z(\ab[11][42] ) );
  AN2P U2047 ( .A(n266), .B(B[41]), .Z(\ab[11][41] ) );
  AN2P U2048 ( .A(n266), .B(B[40]), .Z(\ab[11][40] ) );
  AN2P U2049 ( .A(n266), .B(B[39]), .Z(\ab[11][39] ) );
  AN2P U2050 ( .A(n266), .B(n452), .Z(\ab[11][38] ) );
  AN2P U2051 ( .A(n266), .B(n448), .Z(\ab[11][37] ) );
  AN2P U2052 ( .A(n266), .B(n444), .Z(\ab[11][36] ) );
  AN2P U2053 ( .A(n266), .B(n440), .Z(\ab[11][35] ) );
  AN2P U2054 ( .A(n265), .B(n436), .Z(\ab[11][34] ) );
  AN2P U2055 ( .A(n265), .B(n432), .Z(\ab[11][33] ) );
  AN2P U2056 ( .A(n265), .B(n428), .Z(\ab[11][32] ) );
  AN2P U2057 ( .A(n265), .B(n424), .Z(\ab[11][31] ) );
  AN2P U2058 ( .A(n265), .B(n420), .Z(\ab[11][30] ) );
  AN2P U2059 ( .A(n265), .B(n416), .Z(\ab[11][29] ) );
  AN2P U2060 ( .A(n265), .B(n412), .Z(\ab[11][28] ) );
  AN2P U2061 ( .A(n265), .B(n408), .Z(\ab[11][27] ) );
  AN2P U2062 ( .A(n265), .B(n404), .Z(\ab[11][26] ) );
  AN2P U2063 ( .A(n265), .B(n400), .Z(\ab[11][25] ) );
  AN2P U2064 ( .A(n265), .B(n396), .Z(\ab[11][24] ) );
  AN2P U2065 ( .A(n265), .B(n392), .Z(\ab[11][23] ) );
  AN2P U2066 ( .A(n264), .B(n388), .Z(\ab[11][22] ) );
  AN2P U2067 ( .A(n264), .B(n384), .Z(\ab[11][21] ) );
  AN2P U2068 ( .A(n264), .B(n380), .Z(\ab[11][20] ) );
  AN2P U2069 ( .A(n264), .B(n376), .Z(\ab[11][19] ) );
  AN2P U2070 ( .A(n264), .B(n372), .Z(\ab[11][18] ) );
  AN2P U2071 ( .A(n264), .B(n368), .Z(\ab[11][17] ) );
  AN2P U2072 ( .A(n264), .B(n364), .Z(\ab[11][16] ) );
  AN2P U2073 ( .A(n264), .B(n360), .Z(\ab[11][15] ) );
  AN2P U2074 ( .A(n264), .B(n356), .Z(\ab[11][14] ) );
  AN2P U2075 ( .A(n264), .B(n352), .Z(\ab[11][13] ) );
  AN2P U2076 ( .A(n264), .B(n348), .Z(\ab[11][12] ) );
  AN2P U2077 ( .A(n264), .B(n344), .Z(\ab[11][11] ) );
  AN2P U2078 ( .A(n263), .B(n340), .Z(\ab[11][10] ) );
  AN2P U2079 ( .A(n263), .B(n336), .Z(\ab[11][9] ) );
  AN2P U2080 ( .A(n263), .B(n332), .Z(\ab[11][8] ) );
  AN2P U2081 ( .A(n263), .B(n328), .Z(\ab[11][7] ) );
  AN2P U2082 ( .A(n263), .B(n324), .Z(\ab[11][6] ) );
  AN2P U2083 ( .A(n263), .B(n320), .Z(\ab[11][5] ) );
  AN2P U2084 ( .A(n263), .B(n316), .Z(\ab[11][4] ) );
  AN2P U2085 ( .A(n263), .B(n312), .Z(\ab[11][3] ) );
  AN2P U2086 ( .A(n263), .B(n308), .Z(\ab[11][2] ) );
  AN2P U2087 ( .A(n263), .B(n304), .Z(\ab[11][1] ) );
  AN2P U2088 ( .A(n263), .B(n300), .Z(\ab[11][0] ) );
  AN2P U2089 ( .A(n279), .B(n455), .Z(\ab[12][94] ) );
  AN2P U2090 ( .A(n263), .B(n491), .Z(\ab[11][95] ) );
  AN2P U2091 ( .A(n279), .B(n456), .Z(\ab[12][93] ) );
  AN2P U2092 ( .A(n279), .B(n457), .Z(\ab[12][92] ) );
  AN2P U2093 ( .A(n279), .B(n458), .Z(\ab[12][91] ) );
  AN2P U2094 ( .A(n279), .B(n459), .Z(\ab[12][90] ) );
  AN2P U2095 ( .A(n279), .B(n460), .Z(\ab[12][89] ) );
  AN2P U2096 ( .A(n279), .B(n461), .Z(\ab[12][88] ) );
  AN2P U2097 ( .A(n279), .B(n462), .Z(\ab[12][87] ) );
  AN2P U2098 ( .A(n279), .B(n463), .Z(\ab[12][86] ) );
  AN2P U2099 ( .A(n279), .B(n464), .Z(\ab[12][85] ) );
  AN2P U2100 ( .A(n279), .B(n465), .Z(\ab[12][84] ) );
  AN2P U2101 ( .A(n279), .B(n466), .Z(\ab[12][83] ) );
  AN2P U2102 ( .A(n278), .B(n467), .Z(\ab[12][82] ) );
  AN2P U2103 ( .A(n278), .B(n468), .Z(\ab[12][81] ) );
  AN2P U2104 ( .A(n278), .B(n469), .Z(\ab[12][80] ) );
  AN2P U2105 ( .A(n278), .B(n470), .Z(\ab[12][79] ) );
  AN2P U2106 ( .A(n278), .B(n471), .Z(\ab[12][78] ) );
  AN2P U2107 ( .A(n278), .B(n472), .Z(\ab[12][77] ) );
  AN2P U2108 ( .A(n278), .B(n473), .Z(\ab[12][76] ) );
  AN2P U2109 ( .A(n278), .B(n474), .Z(\ab[12][75] ) );
  AN2P U2110 ( .A(n278), .B(n475), .Z(\ab[12][74] ) );
  AN2P U2111 ( .A(n278), .B(n476), .Z(\ab[12][73] ) );
  AN2P U2112 ( .A(n278), .B(n477), .Z(\ab[12][72] ) );
  AN2P U2113 ( .A(n278), .B(n478), .Z(\ab[12][71] ) );
  AN2P U2114 ( .A(n277), .B(n479), .Z(\ab[12][70] ) );
  AN2P U2115 ( .A(n277), .B(n480), .Z(\ab[12][69] ) );
  AN2P U2116 ( .A(n277), .B(n481), .Z(\ab[12][68] ) );
  AN2P U2117 ( .A(n277), .B(n482), .Z(\ab[12][67] ) );
  AN2P U2118 ( .A(n277), .B(n483), .Z(\ab[12][66] ) );
  AN2P U2119 ( .A(n277), .B(n484), .Z(\ab[12][65] ) );
  AN2P U2120 ( .A(n277), .B(n485), .Z(\ab[12][64] ) );
  AN2P U2121 ( .A(n277), .B(n486), .Z(\ab[12][63] ) );
  AN2P U2122 ( .A(n277), .B(n487), .Z(\ab[12][62] ) );
  AN2P U2123 ( .A(n277), .B(n488), .Z(\ab[12][61] ) );
  AN2P U2124 ( .A(n277), .B(n489), .Z(\ab[12][60] ) );
  AN2P U2125 ( .A(n277), .B(B[59]), .Z(\ab[12][59] ) );
  AN2P U2126 ( .A(n276), .B(B[58]), .Z(\ab[12][58] ) );
  AN2P U2127 ( .A(n276), .B(B[57]), .Z(\ab[12][57] ) );
  AN2P U2128 ( .A(n276), .B(B[56]), .Z(\ab[12][56] ) );
  AN2P U2129 ( .A(n276), .B(n490), .Z(\ab[12][55] ) );
  AN2P U2130 ( .A(n276), .B(B[54]), .Z(\ab[12][54] ) );
  AN2P U2131 ( .A(n276), .B(B[53]), .Z(\ab[12][53] ) );
  AN2P U2132 ( .A(n276), .B(B[52]), .Z(\ab[12][52] ) );
  AN2P U2133 ( .A(n276), .B(B[51]), .Z(\ab[12][51] ) );
  AN2P U2134 ( .A(n276), .B(B[50]), .Z(\ab[12][50] ) );
  AN2P U2135 ( .A(n276), .B(B[49]), .Z(\ab[12][49] ) );
  AN2P U2136 ( .A(n276), .B(B[48]), .Z(\ab[12][48] ) );
  AN2P U2137 ( .A(n276), .B(B[47]), .Z(\ab[12][47] ) );
  AN2P U2138 ( .A(n275), .B(B[46]), .Z(\ab[12][46] ) );
  AN2P U2139 ( .A(n275), .B(B[45]), .Z(\ab[12][45] ) );
  AN2P U2140 ( .A(n275), .B(B[44]), .Z(\ab[12][44] ) );
  AN2P U2141 ( .A(n275), .B(B[43]), .Z(\ab[12][43] ) );
  AN2P U2142 ( .A(n275), .B(B[42]), .Z(\ab[12][42] ) );
  AN2P U2143 ( .A(n275), .B(B[41]), .Z(\ab[12][41] ) );
  AN2P U2144 ( .A(n275), .B(B[40]), .Z(\ab[12][40] ) );
  AN2P U2145 ( .A(n275), .B(B[39]), .Z(\ab[12][39] ) );
  AN2P U2146 ( .A(n275), .B(n452), .Z(\ab[12][38] ) );
  AN2P U2147 ( .A(n275), .B(n448), .Z(\ab[12][37] ) );
  AN2P U2148 ( .A(n275), .B(n444), .Z(\ab[12][36] ) );
  AN2P U2149 ( .A(n275), .B(n440), .Z(\ab[12][35] ) );
  AN2P U2150 ( .A(n274), .B(n436), .Z(\ab[12][34] ) );
  AN2P U2151 ( .A(n274), .B(n432), .Z(\ab[12][33] ) );
  AN2P U2152 ( .A(n274), .B(n428), .Z(\ab[12][32] ) );
  AN2P U2153 ( .A(n274), .B(n424), .Z(\ab[12][31] ) );
  AN2P U2154 ( .A(n274), .B(n420), .Z(\ab[12][30] ) );
  AN2P U2155 ( .A(n274), .B(n416), .Z(\ab[12][29] ) );
  AN2P U2156 ( .A(n274), .B(n412), .Z(\ab[12][28] ) );
  AN2P U2157 ( .A(n274), .B(n408), .Z(\ab[12][27] ) );
  AN2P U2158 ( .A(n274), .B(n404), .Z(\ab[12][26] ) );
  AN2P U2159 ( .A(n274), .B(n400), .Z(\ab[12][25] ) );
  AN2P U2160 ( .A(n274), .B(n396), .Z(\ab[12][24] ) );
  AN2P U2161 ( .A(n274), .B(n392), .Z(\ab[12][23] ) );
  AN2P U2162 ( .A(n273), .B(n388), .Z(\ab[12][22] ) );
  AN2P U2163 ( .A(n273), .B(n384), .Z(\ab[12][21] ) );
  AN2P U2164 ( .A(n273), .B(n380), .Z(\ab[12][20] ) );
  AN2P U2165 ( .A(n273), .B(n376), .Z(\ab[12][19] ) );
  AN2P U2166 ( .A(n273), .B(n372), .Z(\ab[12][18] ) );
  AN2P U2167 ( .A(n273), .B(n368), .Z(\ab[12][17] ) );
  AN2P U2168 ( .A(n273), .B(n364), .Z(\ab[12][16] ) );
  AN2P U2169 ( .A(n273), .B(n360), .Z(\ab[12][15] ) );
  AN2P U2170 ( .A(n273), .B(n356), .Z(\ab[12][14] ) );
  AN2P U2171 ( .A(n273), .B(n352), .Z(\ab[12][13] ) );
  AN2P U2172 ( .A(n273), .B(n348), .Z(\ab[12][12] ) );
  AN2P U2173 ( .A(n273), .B(n344), .Z(\ab[12][11] ) );
  AN2P U2174 ( .A(n272), .B(n340), .Z(\ab[12][10] ) );
  AN2P U2175 ( .A(n272), .B(n336), .Z(\ab[12][9] ) );
  AN2P U2176 ( .A(n272), .B(n332), .Z(\ab[12][8] ) );
  AN2P U2177 ( .A(n272), .B(n328), .Z(\ab[12][7] ) );
  AN2P U2178 ( .A(n272), .B(n324), .Z(\ab[12][6] ) );
  AN2P U2179 ( .A(n272), .B(n320), .Z(\ab[12][5] ) );
  AN2P U2180 ( .A(n272), .B(n316), .Z(\ab[12][4] ) );
  AN2P U2181 ( .A(n272), .B(n312), .Z(\ab[12][3] ) );
  AN2P U2182 ( .A(n272), .B(n308), .Z(\ab[12][2] ) );
  AN2P U2183 ( .A(n272), .B(n304), .Z(\ab[12][1] ) );
  AN2P U2184 ( .A(n272), .B(n300), .Z(\ab[12][0] ) );
  AN2P U2185 ( .A(n288), .B(n455), .Z(\ab[13][94] ) );
  AN2P U2186 ( .A(n272), .B(n491), .Z(\ab[12][95] ) );
  AN2P U2187 ( .A(n288), .B(n456), .Z(\ab[13][93] ) );
  AN2P U2188 ( .A(n288), .B(n457), .Z(\ab[13][92] ) );
  AN2P U2189 ( .A(n288), .B(n458), .Z(\ab[13][91] ) );
  AN2P U2190 ( .A(n288), .B(n459), .Z(\ab[13][90] ) );
  AN2P U2191 ( .A(n288), .B(n460), .Z(\ab[13][89] ) );
  AN2P U2192 ( .A(n288), .B(n461), .Z(\ab[13][88] ) );
  AN2P U2193 ( .A(n288), .B(n462), .Z(\ab[13][87] ) );
  AN2P U2194 ( .A(n288), .B(n463), .Z(\ab[13][86] ) );
  AN2P U2195 ( .A(n288), .B(n464), .Z(\ab[13][85] ) );
  AN2P U2196 ( .A(n288), .B(n465), .Z(\ab[13][84] ) );
  AN2P U2197 ( .A(n288), .B(n466), .Z(\ab[13][83] ) );
  AN2P U2198 ( .A(n287), .B(n467), .Z(\ab[13][82] ) );
  AN2P U2199 ( .A(n287), .B(n468), .Z(\ab[13][81] ) );
  AN2P U2200 ( .A(n287), .B(n469), .Z(\ab[13][80] ) );
  AN2P U2201 ( .A(n287), .B(n470), .Z(\ab[13][79] ) );
  AN2P U2202 ( .A(n287), .B(n471), .Z(\ab[13][78] ) );
  AN2P U2203 ( .A(n287), .B(n472), .Z(\ab[13][77] ) );
  AN2P U2204 ( .A(n287), .B(n473), .Z(\ab[13][76] ) );
  AN2P U2205 ( .A(n287), .B(n474), .Z(\ab[13][75] ) );
  AN2P U2206 ( .A(n287), .B(n475), .Z(\ab[13][74] ) );
  AN2P U2207 ( .A(n287), .B(n476), .Z(\ab[13][73] ) );
  AN2P U2208 ( .A(n287), .B(n477), .Z(\ab[13][72] ) );
  AN2P U2209 ( .A(n287), .B(n478), .Z(\ab[13][71] ) );
  AN2P U2210 ( .A(n286), .B(n479), .Z(\ab[13][70] ) );
  AN2P U2211 ( .A(n286), .B(n480), .Z(\ab[13][69] ) );
  AN2P U2212 ( .A(n286), .B(n481), .Z(\ab[13][68] ) );
  AN2P U2213 ( .A(n286), .B(n482), .Z(\ab[13][67] ) );
  AN2P U2214 ( .A(n286), .B(n483), .Z(\ab[13][66] ) );
  AN2P U2215 ( .A(n286), .B(n484), .Z(\ab[13][65] ) );
  AN2P U2216 ( .A(n286), .B(n485), .Z(\ab[13][64] ) );
  AN2P U2217 ( .A(n286), .B(n486), .Z(\ab[13][63] ) );
  AN2P U2218 ( .A(n286), .B(n487), .Z(\ab[13][62] ) );
  AN2P U2219 ( .A(n286), .B(n488), .Z(\ab[13][61] ) );
  AN2P U2220 ( .A(n286), .B(n489), .Z(\ab[13][60] ) );
  AN2P U2221 ( .A(n286), .B(B[59]), .Z(\ab[13][59] ) );
  AN2P U2222 ( .A(n285), .B(B[58]), .Z(\ab[13][58] ) );
  AN2P U2223 ( .A(n285), .B(B[57]), .Z(\ab[13][57] ) );
  AN2P U2224 ( .A(n285), .B(B[56]), .Z(\ab[13][56] ) );
  AN2P U2225 ( .A(n285), .B(n490), .Z(\ab[13][55] ) );
  AN2P U2226 ( .A(n285), .B(B[54]), .Z(\ab[13][54] ) );
  AN2P U2227 ( .A(n285), .B(B[53]), .Z(\ab[13][53] ) );
  AN2P U2228 ( .A(n285), .B(B[52]), .Z(\ab[13][52] ) );
  AN2P U2229 ( .A(n285), .B(B[51]), .Z(\ab[13][51] ) );
  AN2P U2230 ( .A(n285), .B(B[50]), .Z(\ab[13][50] ) );
  AN2P U2231 ( .A(n285), .B(B[49]), .Z(\ab[13][49] ) );
  AN2P U2232 ( .A(n285), .B(B[48]), .Z(\ab[13][48] ) );
  AN2P U2233 ( .A(n285), .B(B[47]), .Z(\ab[13][47] ) );
  AN2P U2234 ( .A(n284), .B(B[46]), .Z(\ab[13][46] ) );
  AN2P U2235 ( .A(n284), .B(B[45]), .Z(\ab[13][45] ) );
  AN2P U2236 ( .A(n284), .B(B[44]), .Z(\ab[13][44] ) );
  AN2P U2237 ( .A(n284), .B(B[43]), .Z(\ab[13][43] ) );
  AN2P U2238 ( .A(n284), .B(B[42]), .Z(\ab[13][42] ) );
  AN2P U2239 ( .A(n284), .B(B[41]), .Z(\ab[13][41] ) );
  AN2P U2240 ( .A(n284), .B(B[40]), .Z(\ab[13][40] ) );
  AN2P U2241 ( .A(n284), .B(B[39]), .Z(\ab[13][39] ) );
  AN2P U2242 ( .A(n284), .B(n452), .Z(\ab[13][38] ) );
  AN2P U2243 ( .A(n284), .B(n448), .Z(\ab[13][37] ) );
  AN2P U2244 ( .A(n284), .B(n444), .Z(\ab[13][36] ) );
  AN2P U2245 ( .A(n284), .B(n440), .Z(\ab[13][35] ) );
  AN2P U2246 ( .A(n283), .B(n436), .Z(\ab[13][34] ) );
  AN2P U2247 ( .A(n283), .B(n432), .Z(\ab[13][33] ) );
  AN2P U2248 ( .A(n283), .B(n428), .Z(\ab[13][32] ) );
  AN2P U2249 ( .A(n283), .B(n424), .Z(\ab[13][31] ) );
  AN2P U2250 ( .A(n283), .B(n420), .Z(\ab[13][30] ) );
  AN2P U2251 ( .A(n283), .B(n416), .Z(\ab[13][29] ) );
  AN2P U2252 ( .A(n283), .B(n412), .Z(\ab[13][28] ) );
  AN2P U2253 ( .A(n283), .B(n408), .Z(\ab[13][27] ) );
  AN2P U2254 ( .A(n283), .B(n404), .Z(\ab[13][26] ) );
  AN2P U2255 ( .A(n283), .B(n400), .Z(\ab[13][25] ) );
  AN2P U2256 ( .A(n283), .B(n396), .Z(\ab[13][24] ) );
  AN2P U2257 ( .A(n283), .B(n392), .Z(\ab[13][23] ) );
  AN2P U2258 ( .A(n282), .B(n388), .Z(\ab[13][22] ) );
  AN2P U2259 ( .A(n282), .B(n384), .Z(\ab[13][21] ) );
  AN2P U2260 ( .A(n282), .B(n380), .Z(\ab[13][20] ) );
  AN2P U2261 ( .A(n282), .B(n376), .Z(\ab[13][19] ) );
  AN2P U2262 ( .A(n282), .B(n372), .Z(\ab[13][18] ) );
  AN2P U2263 ( .A(n282), .B(n368), .Z(\ab[13][17] ) );
  AN2P U2264 ( .A(n282), .B(n364), .Z(\ab[13][16] ) );
  AN2P U2265 ( .A(n282), .B(n360), .Z(\ab[13][15] ) );
  AN2P U2266 ( .A(n282), .B(n356), .Z(\ab[13][14] ) );
  AN2P U2267 ( .A(n282), .B(n352), .Z(\ab[13][13] ) );
  AN2P U2268 ( .A(n282), .B(n348), .Z(\ab[13][12] ) );
  AN2P U2269 ( .A(n282), .B(n344), .Z(\ab[13][11] ) );
  AN2P U2270 ( .A(n281), .B(n340), .Z(\ab[13][10] ) );
  AN2P U2271 ( .A(n281), .B(n336), .Z(\ab[13][9] ) );
  AN2P U2272 ( .A(n281), .B(n332), .Z(\ab[13][8] ) );
  AN2P U2273 ( .A(n281), .B(n328), .Z(\ab[13][7] ) );
  AN2P U2274 ( .A(n281), .B(n324), .Z(\ab[13][6] ) );
  AN2P U2275 ( .A(n281), .B(n320), .Z(\ab[13][5] ) );
  AN2P U2276 ( .A(n281), .B(n316), .Z(\ab[13][4] ) );
  AN2P U2277 ( .A(n281), .B(n312), .Z(\ab[13][3] ) );
  AN2P U2278 ( .A(n281), .B(n308), .Z(\ab[13][2] ) );
  AN2P U2279 ( .A(n281), .B(n304), .Z(\ab[13][1] ) );
  AN2P U2280 ( .A(n281), .B(n300), .Z(\ab[13][0] ) );
  AN2P U2281 ( .A(n297), .B(n455), .Z(\ab[14][94] ) );
  AN2P U2282 ( .A(n281), .B(n491), .Z(\ab[13][95] ) );
  AN2P U2283 ( .A(n297), .B(n456), .Z(\ab[14][93] ) );
  AN2P U2284 ( .A(n297), .B(n457), .Z(\ab[14][92] ) );
  AN2P U2285 ( .A(n297), .B(n458), .Z(\ab[14][91] ) );
  AN2P U2286 ( .A(n297), .B(n459), .Z(\ab[14][90] ) );
  AN2P U2287 ( .A(n297), .B(n460), .Z(\ab[14][89] ) );
  AN2P U2288 ( .A(n297), .B(n461), .Z(\ab[14][88] ) );
  AN2P U2289 ( .A(n297), .B(n462), .Z(\ab[14][87] ) );
  AN2P U2290 ( .A(n297), .B(n463), .Z(\ab[14][86] ) );
  AN2P U2291 ( .A(n297), .B(n464), .Z(\ab[14][85] ) );
  AN2P U2292 ( .A(n297), .B(n465), .Z(\ab[14][84] ) );
  AN2P U2293 ( .A(n297), .B(n466), .Z(\ab[14][83] ) );
  AN2P U2294 ( .A(n296), .B(n467), .Z(\ab[14][82] ) );
  AN2P U2295 ( .A(n296), .B(n468), .Z(\ab[14][81] ) );
  AN2P U2296 ( .A(n296), .B(n469), .Z(\ab[14][80] ) );
  AN2P U2297 ( .A(n296), .B(n470), .Z(\ab[14][79] ) );
  AN2P U2298 ( .A(n296), .B(n471), .Z(\ab[14][78] ) );
  AN2P U2299 ( .A(n296), .B(n472), .Z(\ab[14][77] ) );
  AN2P U2300 ( .A(n296), .B(n473), .Z(\ab[14][76] ) );
  AN2P U2301 ( .A(n296), .B(n474), .Z(\ab[14][75] ) );
  AN2P U2302 ( .A(n296), .B(n475), .Z(\ab[14][74] ) );
  AN2P U2303 ( .A(n296), .B(n476), .Z(\ab[14][73] ) );
  AN2P U2304 ( .A(n296), .B(n477), .Z(\ab[14][72] ) );
  AN2P U2305 ( .A(n296), .B(n478), .Z(\ab[14][71] ) );
  AN2P U2306 ( .A(n295), .B(n479), .Z(\ab[14][70] ) );
  AN2P U2307 ( .A(n295), .B(n480), .Z(\ab[14][69] ) );
  AN2P U2308 ( .A(n295), .B(n481), .Z(\ab[14][68] ) );
  AN2P U2309 ( .A(n295), .B(n482), .Z(\ab[14][67] ) );
  AN2P U2310 ( .A(n295), .B(n483), .Z(\ab[14][66] ) );
  AN2P U2311 ( .A(n295), .B(n484), .Z(\ab[14][65] ) );
  AN2P U2312 ( .A(n295), .B(n485), .Z(\ab[14][64] ) );
  AN2P U2313 ( .A(n295), .B(n486), .Z(\ab[14][63] ) );
  AN2P U2314 ( .A(n295), .B(n487), .Z(\ab[14][62] ) );
  AN2P U2315 ( .A(n295), .B(n488), .Z(\ab[14][61] ) );
  AN2P U2316 ( .A(n295), .B(n489), .Z(\ab[14][60] ) );
  AN2P U2317 ( .A(n295), .B(B[59]), .Z(\ab[14][59] ) );
  AN2P U2318 ( .A(n294), .B(B[58]), .Z(\ab[14][58] ) );
  AN2P U2319 ( .A(n294), .B(B[57]), .Z(\ab[14][57] ) );
  AN2P U2320 ( .A(n294), .B(B[56]), .Z(\ab[14][56] ) );
  AN2P U2321 ( .A(n294), .B(n490), .Z(\ab[14][55] ) );
  AN2P U2322 ( .A(n294), .B(B[54]), .Z(\ab[14][54] ) );
  AN2P U2323 ( .A(n294), .B(B[53]), .Z(\ab[14][53] ) );
  AN2P U2324 ( .A(n294), .B(B[52]), .Z(\ab[14][52] ) );
  AN2P U2325 ( .A(n294), .B(B[51]), .Z(\ab[14][51] ) );
  AN2P U2326 ( .A(n294), .B(B[50]), .Z(\ab[14][50] ) );
  AN2P U2327 ( .A(n294), .B(B[49]), .Z(\ab[14][49] ) );
  AN2P U2328 ( .A(n294), .B(B[48]), .Z(\ab[14][48] ) );
  AN2P U2329 ( .A(n294), .B(B[47]), .Z(\ab[14][47] ) );
  AN2P U2330 ( .A(n293), .B(B[46]), .Z(\ab[14][46] ) );
  AN2P U2331 ( .A(n293), .B(B[45]), .Z(\ab[14][45] ) );
  AN2P U2332 ( .A(n293), .B(B[44]), .Z(\ab[14][44] ) );
  AN2P U2333 ( .A(n293), .B(B[43]), .Z(\ab[14][43] ) );
  AN2P U2334 ( .A(n293), .B(B[42]), .Z(\ab[14][42] ) );
  AN2P U2335 ( .A(n293), .B(B[41]), .Z(\ab[14][41] ) );
  AN2P U2336 ( .A(n293), .B(B[40]), .Z(\ab[14][40] ) );
  AN2P U2337 ( .A(n293), .B(B[39]), .Z(\ab[14][39] ) );
  AN2P U2338 ( .A(n293), .B(n452), .Z(\ab[14][38] ) );
  AN2P U2339 ( .A(n293), .B(n448), .Z(\ab[14][37] ) );
  AN2P U2340 ( .A(n293), .B(n444), .Z(\ab[14][36] ) );
  AN2P U2341 ( .A(n293), .B(n440), .Z(\ab[14][35] ) );
  AN2P U2342 ( .A(n292), .B(n436), .Z(\ab[14][34] ) );
  AN2P U2343 ( .A(n292), .B(n432), .Z(\ab[14][33] ) );
  AN2P U2344 ( .A(n292), .B(n428), .Z(\ab[14][32] ) );
  AN2P U2345 ( .A(n292), .B(n424), .Z(\ab[14][31] ) );
  AN2P U2346 ( .A(n292), .B(n420), .Z(\ab[14][30] ) );
  AN2P U2347 ( .A(n292), .B(n416), .Z(\ab[14][29] ) );
  AN2P U2348 ( .A(n292), .B(n412), .Z(\ab[14][28] ) );
  AN2P U2349 ( .A(n292), .B(n408), .Z(\ab[14][27] ) );
  AN2P U2350 ( .A(n292), .B(n404), .Z(\ab[14][26] ) );
  AN2P U2351 ( .A(n292), .B(n400), .Z(\ab[14][25] ) );
  AN2P U2352 ( .A(n292), .B(n396), .Z(\ab[14][24] ) );
  AN2P U2353 ( .A(n292), .B(n392), .Z(\ab[14][23] ) );
  AN2P U2354 ( .A(n291), .B(n388), .Z(\ab[14][22] ) );
  AN2P U2355 ( .A(n291), .B(n384), .Z(\ab[14][21] ) );
  AN2P U2356 ( .A(n291), .B(n380), .Z(\ab[14][20] ) );
  AN2P U2357 ( .A(n291), .B(n376), .Z(\ab[14][19] ) );
  AN2P U2358 ( .A(n291), .B(n372), .Z(\ab[14][18] ) );
  AN2P U2359 ( .A(n291), .B(n368), .Z(\ab[14][17] ) );
  AN2P U2360 ( .A(n291), .B(n364), .Z(\ab[14][16] ) );
  AN2P U2361 ( .A(n291), .B(n360), .Z(\ab[14][15] ) );
  AN2P U2362 ( .A(n291), .B(n356), .Z(\ab[14][14] ) );
  AN2P U2363 ( .A(n291), .B(n352), .Z(\ab[14][13] ) );
  AN2P U2364 ( .A(n291), .B(n348), .Z(\ab[14][12] ) );
  AN2P U2365 ( .A(n291), .B(n344), .Z(\ab[14][11] ) );
  AN2P U2366 ( .A(n290), .B(n340), .Z(\ab[14][10] ) );
  AN2P U2367 ( .A(n290), .B(n336), .Z(\ab[14][9] ) );
  AN2P U2368 ( .A(n290), .B(n332), .Z(\ab[14][8] ) );
  AN2P U2369 ( .A(n290), .B(n328), .Z(\ab[14][7] ) );
  AN2P U2370 ( .A(n290), .B(n324), .Z(\ab[14][6] ) );
  AN2P U2371 ( .A(n290), .B(n320), .Z(\ab[14][5] ) );
  AN2P U2372 ( .A(n290), .B(n316), .Z(\ab[14][4] ) );
  AN2P U2373 ( .A(n290), .B(n312), .Z(\ab[14][3] ) );
  AN2P U2374 ( .A(n290), .B(n308), .Z(\ab[14][2] ) );
  AN2P U2375 ( .A(n290), .B(n304), .Z(\ab[14][1] ) );
  AN2P U2376 ( .A(n290), .B(n300), .Z(\ab[14][0] ) );
  AN2P U2377 ( .A(n290), .B(n491), .Z(\ab[14][95] ) );
  AN2P U2378 ( .A(n452), .B(n11), .Z(\ab[15][38] ) );
  AN2P U2379 ( .A(n448), .B(n11), .Z(\ab[15][37] ) );
  AN2P U2380 ( .A(n444), .B(n11), .Z(\ab[15][36] ) );
  AN2P U2381 ( .A(n440), .B(n11), .Z(\ab[15][35] ) );
  AN2P U2382 ( .A(n436), .B(n11), .Z(\ab[15][34] ) );
  AN2P U2383 ( .A(n432), .B(n11), .Z(\ab[15][33] ) );
  AN2P U2384 ( .A(n428), .B(n11), .Z(\ab[15][32] ) );
  AN2P U2385 ( .A(n424), .B(n11), .Z(\ab[15][31] ) );
  AN2P U2386 ( .A(n420), .B(n12), .Z(\ab[15][30] ) );
  AN2P U2387 ( .A(n416), .B(n12), .Z(\ab[15][29] ) );
  AN2P U2388 ( .A(n412), .B(n12), .Z(\ab[15][28] ) );
  AN2P U2389 ( .A(n408), .B(n12), .Z(\ab[15][27] ) );
  AN2P U2390 ( .A(n404), .B(n12), .Z(\ab[15][26] ) );
  AN2P U2391 ( .A(n400), .B(n12), .Z(\ab[15][25] ) );
  AN2P U2392 ( .A(n396), .B(n12), .Z(\ab[15][24] ) );
  AN2P U2393 ( .A(n392), .B(n12), .Z(\ab[15][23] ) );
  AN2P U2394 ( .A(n388), .B(n13), .Z(\ab[15][22] ) );
  AN2P U2395 ( .A(n384), .B(n13), .Z(\ab[15][21] ) );
  AN2P U2396 ( .A(n380), .B(n13), .Z(\ab[15][20] ) );
  AN2P U2397 ( .A(n376), .B(n13), .Z(\ab[15][19] ) );
  AN2P U2398 ( .A(n372), .B(n13), .Z(\ab[15][18] ) );
  AN2P U2399 ( .A(n368), .B(n13), .Z(\ab[15][17] ) );
  AN2P U2400 ( .A(n364), .B(n13), .Z(\ab[15][16] ) );
  AN2P U2401 ( .A(n360), .B(n13), .Z(\ab[15][15] ) );
  AN2P U2402 ( .A(n356), .B(n14), .Z(\ab[15][14] ) );
  AN2P U2403 ( .A(n352), .B(n14), .Z(\ab[15][13] ) );
  AN2P U2404 ( .A(n348), .B(n14), .Z(\ab[15][12] ) );
  AN2P U2405 ( .A(n344), .B(n14), .Z(\ab[15][11] ) );
  AN2P U2406 ( .A(n340), .B(n14), .Z(\ab[15][10] ) );
  AN2P U2407 ( .A(n336), .B(n14), .Z(\ab[15][9] ) );
  AN2P U2408 ( .A(n332), .B(n14), .Z(\ab[15][8] ) );
  AN2P U2409 ( .A(n328), .B(n14), .Z(\ab[15][7] ) );
  AN2P U2410 ( .A(n324), .B(n15), .Z(\ab[15][6] ) );
  AN2P U2411 ( .A(n320), .B(n15), .Z(\ab[15][5] ) );
  AN2P U2412 ( .A(n316), .B(n15), .Z(\ab[15][4] ) );
  AN2P U2413 ( .A(n312), .B(n15), .Z(\ab[15][3] ) );
  AN2P U2414 ( .A(n308), .B(n15), .Z(\ab[15][2] ) );
  AN2P U2415 ( .A(n304), .B(n15), .Z(\ab[15][1] ) );
  AN2P U2416 ( .A(n300), .B(n15), .Z(\ab[15][0] ) );
  AN2P U2417 ( .A(n452), .B(n159), .Z(\ab[16][38] ) );
  AN2P U2418 ( .A(n448), .B(n159), .Z(\ab[16][37] ) );
  AN2P U2419 ( .A(n444), .B(n159), .Z(\ab[16][36] ) );
  AN2P U2420 ( .A(n440), .B(n159), .Z(\ab[16][35] ) );
  AN2P U2421 ( .A(n436), .B(n159), .Z(\ab[16][34] ) );
  AN2P U2422 ( .A(n432), .B(n159), .Z(\ab[16][33] ) );
  AN2P U2423 ( .A(n428), .B(n159), .Z(\ab[16][32] ) );
  AN2P U2424 ( .A(n424), .B(n159), .Z(\ab[16][31] ) );
  AN2P U2425 ( .A(n420), .B(n160), .Z(\ab[16][30] ) );
  AN2P U2426 ( .A(n416), .B(n160), .Z(\ab[16][29] ) );
  AN2P U2427 ( .A(n412), .B(n160), .Z(\ab[16][28] ) );
  AN2P U2428 ( .A(n408), .B(n160), .Z(\ab[16][27] ) );
  AN2P U2429 ( .A(n404), .B(n160), .Z(\ab[16][26] ) );
  AN2P U2430 ( .A(n400), .B(n160), .Z(\ab[16][25] ) );
  AN2P U2431 ( .A(n396), .B(n160), .Z(\ab[16][24] ) );
  AN2P U2432 ( .A(n392), .B(n160), .Z(\ab[16][23] ) );
  AN2P U2433 ( .A(n388), .B(n161), .Z(\ab[16][22] ) );
  AN2P U2434 ( .A(n384), .B(n161), .Z(\ab[16][21] ) );
  AN2P U2435 ( .A(n380), .B(n161), .Z(\ab[16][20] ) );
  AN2P U2436 ( .A(n376), .B(n161), .Z(\ab[16][19] ) );
  AN2P U2437 ( .A(n372), .B(n161), .Z(\ab[16][18] ) );
  AN2P U2438 ( .A(n368), .B(n161), .Z(\ab[16][17] ) );
  AN2P U2439 ( .A(n364), .B(n161), .Z(\ab[16][16] ) );
  AN2P U2440 ( .A(n360), .B(n161), .Z(\ab[16][15] ) );
  AN2P U2441 ( .A(n356), .B(n162), .Z(\ab[16][14] ) );
  AN2P U2442 ( .A(n352), .B(n162), .Z(\ab[16][13] ) );
  AN2P U2443 ( .A(n348), .B(n162), .Z(\ab[16][12] ) );
  AN2P U2444 ( .A(n344), .B(n162), .Z(\ab[16][11] ) );
  AN2P U2445 ( .A(n340), .B(n162), .Z(\ab[16][10] ) );
  AN2P U2446 ( .A(n336), .B(n162), .Z(\ab[16][9] ) );
  AN2P U2447 ( .A(n332), .B(n162), .Z(\ab[16][8] ) );
  AN2P U2448 ( .A(n328), .B(n162), .Z(\ab[16][7] ) );
  AN2P U2449 ( .A(n324), .B(n163), .Z(\ab[16][6] ) );
  AN2P U2450 ( .A(n320), .B(n163), .Z(\ab[16][5] ) );
  AN2P U2451 ( .A(n316), .B(n163), .Z(\ab[16][4] ) );
  AN2P U2452 ( .A(n312), .B(n163), .Z(\ab[16][3] ) );
  AN2P U2453 ( .A(n308), .B(n163), .Z(\ab[16][2] ) );
  AN2P U2454 ( .A(n304), .B(n163), .Z(\ab[16][1] ) );
  AN2P U2455 ( .A(n300), .B(n163), .Z(\ab[16][0] ) );
  AN2P U2456 ( .A(n452), .B(n148), .Z(\ab[17][38] ) );
  AN2P U2457 ( .A(n448), .B(n148), .Z(\ab[17][37] ) );
  AN2P U2458 ( .A(n444), .B(n148), .Z(\ab[17][36] ) );
  AN2P U2459 ( .A(n440), .B(n148), .Z(\ab[17][35] ) );
  AN2P U2460 ( .A(n436), .B(n148), .Z(\ab[17][34] ) );
  AN2P U2461 ( .A(n432), .B(n148), .Z(\ab[17][33] ) );
  AN2P U2462 ( .A(n428), .B(n148), .Z(\ab[17][32] ) );
  AN2P U2463 ( .A(n424), .B(n148), .Z(\ab[17][31] ) );
  AN2P U2464 ( .A(n420), .B(n149), .Z(\ab[17][30] ) );
  AN2P U2465 ( .A(n416), .B(n149), .Z(\ab[17][29] ) );
  AN2P U2466 ( .A(n412), .B(n149), .Z(\ab[17][28] ) );
  AN2P U2467 ( .A(n408), .B(n149), .Z(\ab[17][27] ) );
  AN2P U2468 ( .A(n404), .B(n149), .Z(\ab[17][26] ) );
  AN2P U2469 ( .A(n400), .B(n149), .Z(\ab[17][25] ) );
  AN2P U2470 ( .A(n396), .B(n149), .Z(\ab[17][24] ) );
  AN2P U2471 ( .A(n392), .B(n149), .Z(\ab[17][23] ) );
  AN2P U2472 ( .A(n388), .B(n150), .Z(\ab[17][22] ) );
  AN2P U2473 ( .A(n384), .B(n150), .Z(\ab[17][21] ) );
  AN2P U2474 ( .A(n380), .B(n150), .Z(\ab[17][20] ) );
  AN2P U2475 ( .A(n376), .B(n150), .Z(\ab[17][19] ) );
  AN2P U2476 ( .A(n372), .B(n150), .Z(\ab[17][18] ) );
  AN2P U2477 ( .A(n368), .B(n150), .Z(\ab[17][17] ) );
  AN2P U2478 ( .A(n364), .B(n150), .Z(\ab[17][16] ) );
  AN2P U2479 ( .A(n360), .B(n150), .Z(\ab[17][15] ) );
  AN2P U2480 ( .A(n356), .B(n151), .Z(\ab[17][14] ) );
  AN2P U2481 ( .A(n352), .B(n151), .Z(\ab[17][13] ) );
  AN2P U2482 ( .A(n348), .B(n151), .Z(\ab[17][12] ) );
  AN2P U2483 ( .A(n344), .B(n151), .Z(\ab[17][11] ) );
  AN2P U2484 ( .A(n340), .B(n151), .Z(\ab[17][10] ) );
  AN2P U2485 ( .A(n336), .B(n151), .Z(\ab[17][9] ) );
  AN2P U2486 ( .A(n332), .B(n151), .Z(\ab[17][8] ) );
  AN2P U2487 ( .A(n328), .B(n151), .Z(\ab[17][7] ) );
  AN2P U2488 ( .A(n324), .B(n152), .Z(\ab[17][6] ) );
  AN2P U2489 ( .A(n320), .B(n152), .Z(\ab[17][5] ) );
  AN2P U2490 ( .A(n316), .B(n152), .Z(\ab[17][4] ) );
  AN2P U2491 ( .A(n312), .B(n152), .Z(\ab[17][3] ) );
  AN2P U2492 ( .A(n308), .B(n152), .Z(\ab[17][2] ) );
  AN2P U2493 ( .A(n304), .B(n152), .Z(\ab[17][1] ) );
  AN2P U2494 ( .A(n300), .B(n152), .Z(\ab[17][0] ) );
  AN2P U2495 ( .A(n451), .B(n137), .Z(\ab[18][38] ) );
  AN2P U2496 ( .A(n447), .B(n137), .Z(\ab[18][37] ) );
  AN2P U2497 ( .A(n443), .B(n137), .Z(\ab[18][36] ) );
  AN2P U2498 ( .A(n439), .B(n137), .Z(\ab[18][35] ) );
  AN2P U2499 ( .A(n435), .B(n137), .Z(\ab[18][34] ) );
  AN2P U2500 ( .A(n431), .B(n137), .Z(\ab[18][33] ) );
  AN2P U2501 ( .A(n427), .B(n137), .Z(\ab[18][32] ) );
  AN2P U2502 ( .A(n423), .B(n137), .Z(\ab[18][31] ) );
  AN2P U2503 ( .A(n419), .B(n138), .Z(\ab[18][30] ) );
  AN2P U2504 ( .A(n415), .B(n138), .Z(\ab[18][29] ) );
  AN2P U2505 ( .A(n411), .B(n138), .Z(\ab[18][28] ) );
  AN2P U2506 ( .A(n407), .B(n138), .Z(\ab[18][27] ) );
  AN2P U2507 ( .A(n403), .B(n138), .Z(\ab[18][26] ) );
  AN2P U2508 ( .A(n399), .B(n138), .Z(\ab[18][25] ) );
  AN2P U2509 ( .A(n395), .B(n138), .Z(\ab[18][24] ) );
  AN2P U2510 ( .A(n391), .B(n138), .Z(\ab[18][23] ) );
  AN2P U2511 ( .A(n387), .B(n139), .Z(\ab[18][22] ) );
  AN2P U2512 ( .A(n383), .B(n139), .Z(\ab[18][21] ) );
  AN2P U2513 ( .A(n379), .B(n139), .Z(\ab[18][20] ) );
  AN2P U2514 ( .A(n375), .B(n139), .Z(\ab[18][19] ) );
  AN2P U2515 ( .A(n371), .B(n139), .Z(\ab[18][18] ) );
  AN2P U2516 ( .A(n367), .B(n139), .Z(\ab[18][17] ) );
  AN2P U2517 ( .A(n363), .B(n139), .Z(\ab[18][16] ) );
  AN2P U2518 ( .A(n359), .B(n139), .Z(\ab[18][15] ) );
  AN2P U2519 ( .A(n355), .B(n140), .Z(\ab[18][14] ) );
  AN2P U2520 ( .A(n351), .B(n140), .Z(\ab[18][13] ) );
  AN2P U2521 ( .A(n347), .B(n140), .Z(\ab[18][12] ) );
  AN2P U2522 ( .A(n343), .B(n140), .Z(\ab[18][11] ) );
  AN2P U2523 ( .A(n339), .B(n140), .Z(\ab[18][10] ) );
  AN2P U2524 ( .A(n335), .B(n140), .Z(\ab[18][9] ) );
  AN2P U2525 ( .A(n331), .B(n140), .Z(\ab[18][8] ) );
  AN2P U2526 ( .A(n327), .B(n140), .Z(\ab[18][7] ) );
  AN2P U2527 ( .A(n323), .B(n141), .Z(\ab[18][6] ) );
  AN2P U2528 ( .A(n319), .B(n141), .Z(\ab[18][5] ) );
  AN2P U2529 ( .A(n315), .B(n141), .Z(\ab[18][4] ) );
  AN2P U2530 ( .A(n311), .B(n141), .Z(\ab[18][3] ) );
  AN2P U2531 ( .A(n307), .B(n141), .Z(\ab[18][2] ) );
  AN2P U2532 ( .A(n303), .B(n141), .Z(\ab[18][1] ) );
  AN2P U2533 ( .A(n299), .B(n141), .Z(\ab[18][0] ) );
  AN2P U2534 ( .A(n451), .B(n126), .Z(\ab[19][38] ) );
  AN2P U2535 ( .A(n447), .B(n126), .Z(\ab[19][37] ) );
  AN2P U2536 ( .A(n443), .B(n126), .Z(\ab[19][36] ) );
  AN2P U2537 ( .A(n439), .B(n126), .Z(\ab[19][35] ) );
  AN2P U2538 ( .A(n435), .B(n126), .Z(\ab[19][34] ) );
  AN2P U2539 ( .A(n431), .B(n126), .Z(\ab[19][33] ) );
  AN2P U2540 ( .A(n427), .B(n126), .Z(\ab[19][32] ) );
  AN2P U2541 ( .A(n423), .B(n126), .Z(\ab[19][31] ) );
  AN2P U2542 ( .A(n419), .B(n127), .Z(\ab[19][30] ) );
  AN2P U2543 ( .A(n415), .B(n127), .Z(\ab[19][29] ) );
  AN2P U2544 ( .A(n411), .B(n127), .Z(\ab[19][28] ) );
  AN2P U2545 ( .A(n407), .B(n127), .Z(\ab[19][27] ) );
  AN2P U2546 ( .A(n403), .B(n127), .Z(\ab[19][26] ) );
  AN2P U2547 ( .A(n399), .B(n127), .Z(\ab[19][25] ) );
  AN2P U2548 ( .A(n395), .B(n127), .Z(\ab[19][24] ) );
  AN2P U2549 ( .A(n391), .B(n127), .Z(\ab[19][23] ) );
  AN2P U2550 ( .A(n387), .B(n128), .Z(\ab[19][22] ) );
  AN2P U2551 ( .A(n383), .B(n128), .Z(\ab[19][21] ) );
  AN2P U2552 ( .A(n379), .B(n128), .Z(\ab[19][20] ) );
  AN2P U2553 ( .A(n375), .B(n128), .Z(\ab[19][19] ) );
  AN2P U2554 ( .A(n371), .B(n128), .Z(\ab[19][18] ) );
  AN2P U2555 ( .A(n367), .B(n128), .Z(\ab[19][17] ) );
  AN2P U2556 ( .A(n363), .B(n128), .Z(\ab[19][16] ) );
  AN2P U2557 ( .A(n359), .B(n128), .Z(\ab[19][15] ) );
  AN2P U2558 ( .A(n355), .B(n129), .Z(\ab[19][14] ) );
  AN2P U2559 ( .A(n351), .B(n129), .Z(\ab[19][13] ) );
  AN2P U2560 ( .A(n347), .B(n129), .Z(\ab[19][12] ) );
  AN2P U2561 ( .A(n343), .B(n129), .Z(\ab[19][11] ) );
  AN2P U2562 ( .A(n339), .B(n129), .Z(\ab[19][10] ) );
  AN2P U2563 ( .A(n335), .B(n129), .Z(\ab[19][9] ) );
  AN2P U2564 ( .A(n331), .B(n129), .Z(\ab[19][8] ) );
  AN2P U2565 ( .A(n327), .B(n129), .Z(\ab[19][7] ) );
  AN2P U2566 ( .A(n323), .B(n130), .Z(\ab[19][6] ) );
  AN2P U2567 ( .A(n319), .B(n130), .Z(\ab[19][5] ) );
  AN2P U2568 ( .A(n315), .B(n130), .Z(\ab[19][4] ) );
  AN2P U2569 ( .A(n311), .B(n130), .Z(\ab[19][3] ) );
  AN2P U2570 ( .A(n307), .B(n130), .Z(\ab[19][2] ) );
  AN2P U2571 ( .A(n303), .B(n130), .Z(\ab[19][1] ) );
  AN2P U2572 ( .A(n299), .B(n130), .Z(\ab[19][0] ) );
  AN2P U2573 ( .A(n451), .B(n115), .Z(\ab[20][38] ) );
  AN2P U2574 ( .A(n447), .B(n115), .Z(\ab[20][37] ) );
  AN2P U2575 ( .A(n443), .B(n115), .Z(\ab[20][36] ) );
  AN2P U2576 ( .A(n439), .B(n115), .Z(\ab[20][35] ) );
  AN2P U2577 ( .A(n435), .B(n115), .Z(\ab[20][34] ) );
  AN2P U2578 ( .A(n431), .B(n115), .Z(\ab[20][33] ) );
  AN2P U2579 ( .A(n427), .B(n115), .Z(\ab[20][32] ) );
  AN2P U2580 ( .A(n423), .B(n115), .Z(\ab[20][31] ) );
  AN2P U2581 ( .A(n419), .B(n116), .Z(\ab[20][30] ) );
  AN2P U2582 ( .A(n415), .B(n116), .Z(\ab[20][29] ) );
  AN2P U2583 ( .A(n411), .B(n116), .Z(\ab[20][28] ) );
  AN2P U2584 ( .A(n407), .B(n116), .Z(\ab[20][27] ) );
  AN2P U2585 ( .A(n403), .B(n116), .Z(\ab[20][26] ) );
  AN2P U2586 ( .A(n399), .B(n116), .Z(\ab[20][25] ) );
  AN2P U2587 ( .A(n395), .B(n116), .Z(\ab[20][24] ) );
  AN2P U2588 ( .A(n391), .B(n116), .Z(\ab[20][23] ) );
  AN2P U2589 ( .A(n387), .B(n117), .Z(\ab[20][22] ) );
  AN2P U2590 ( .A(n383), .B(n117), .Z(\ab[20][21] ) );
  AN2P U2591 ( .A(n379), .B(n117), .Z(\ab[20][20] ) );
  AN2P U2592 ( .A(n375), .B(n117), .Z(\ab[20][19] ) );
  AN2P U2593 ( .A(n371), .B(n117), .Z(\ab[20][18] ) );
  AN2P U2594 ( .A(n367), .B(n117), .Z(\ab[20][17] ) );
  AN2P U2595 ( .A(n363), .B(n117), .Z(\ab[20][16] ) );
  AN2P U2596 ( .A(n359), .B(n117), .Z(\ab[20][15] ) );
  AN2P U2597 ( .A(n355), .B(n118), .Z(\ab[20][14] ) );
  AN2P U2598 ( .A(n351), .B(n118), .Z(\ab[20][13] ) );
  AN2P U2599 ( .A(n347), .B(n118), .Z(\ab[20][12] ) );
  AN2P U2600 ( .A(n343), .B(n118), .Z(\ab[20][11] ) );
  AN2P U2601 ( .A(n339), .B(n118), .Z(\ab[20][10] ) );
  AN2P U2602 ( .A(n335), .B(n118), .Z(\ab[20][9] ) );
  AN2P U2603 ( .A(n331), .B(n118), .Z(\ab[20][8] ) );
  AN2P U2604 ( .A(n327), .B(n118), .Z(\ab[20][7] ) );
  AN2P U2605 ( .A(n323), .B(n119), .Z(\ab[20][6] ) );
  AN2P U2606 ( .A(n319), .B(n119), .Z(\ab[20][5] ) );
  AN2P U2607 ( .A(n315), .B(n119), .Z(\ab[20][4] ) );
  AN2P U2608 ( .A(n311), .B(n119), .Z(\ab[20][3] ) );
  AN2P U2609 ( .A(n307), .B(n119), .Z(\ab[20][2] ) );
  AN2P U2610 ( .A(n303), .B(n119), .Z(\ab[20][1] ) );
  AN2P U2611 ( .A(n299), .B(n119), .Z(\ab[20][0] ) );
  AN2P U2612 ( .A(n451), .B(n104), .Z(\ab[21][38] ) );
  AN2P U2613 ( .A(n447), .B(n104), .Z(\ab[21][37] ) );
  AN2P U2614 ( .A(n443), .B(n104), .Z(\ab[21][36] ) );
  AN2P U2615 ( .A(n439), .B(n104), .Z(\ab[21][35] ) );
  AN2P U2616 ( .A(n435), .B(n104), .Z(\ab[21][34] ) );
  AN2P U2617 ( .A(n431), .B(n104), .Z(\ab[21][33] ) );
  AN2P U2618 ( .A(n427), .B(n104), .Z(\ab[21][32] ) );
  AN2P U2619 ( .A(n423), .B(n104), .Z(\ab[21][31] ) );
  AN2P U2620 ( .A(n419), .B(n105), .Z(\ab[21][30] ) );
  AN2P U2621 ( .A(n415), .B(n105), .Z(\ab[21][29] ) );
  AN2P U2622 ( .A(n411), .B(n105), .Z(\ab[21][28] ) );
  AN2P U2623 ( .A(n407), .B(n105), .Z(\ab[21][27] ) );
  AN2P U2624 ( .A(n403), .B(n105), .Z(\ab[21][26] ) );
  AN2P U2625 ( .A(n399), .B(n105), .Z(\ab[21][25] ) );
  AN2P U2626 ( .A(n395), .B(n105), .Z(\ab[21][24] ) );
  AN2P U2627 ( .A(n391), .B(n105), .Z(\ab[21][23] ) );
  AN2P U2628 ( .A(n387), .B(n106), .Z(\ab[21][22] ) );
  AN2P U2629 ( .A(n383), .B(n106), .Z(\ab[21][21] ) );
  AN2P U2630 ( .A(n379), .B(n106), .Z(\ab[21][20] ) );
  AN2P U2631 ( .A(n375), .B(n106), .Z(\ab[21][19] ) );
  AN2P U2632 ( .A(n371), .B(n106), .Z(\ab[21][18] ) );
  AN2P U2633 ( .A(n367), .B(n106), .Z(\ab[21][17] ) );
  AN2P U2634 ( .A(n363), .B(n106), .Z(\ab[21][16] ) );
  AN2P U2635 ( .A(n359), .B(n106), .Z(\ab[21][15] ) );
  AN2P U2636 ( .A(n355), .B(n107), .Z(\ab[21][14] ) );
  AN2P U2637 ( .A(n351), .B(n107), .Z(\ab[21][13] ) );
  AN2P U2638 ( .A(n347), .B(n107), .Z(\ab[21][12] ) );
  AN2P U2639 ( .A(n343), .B(n107), .Z(\ab[21][11] ) );
  AN2P U2640 ( .A(n339), .B(n107), .Z(\ab[21][10] ) );
  AN2P U2641 ( .A(n335), .B(n107), .Z(\ab[21][9] ) );
  AN2P U2642 ( .A(n331), .B(n107), .Z(\ab[21][8] ) );
  AN2P U2643 ( .A(n327), .B(n107), .Z(\ab[21][7] ) );
  AN2P U2644 ( .A(n323), .B(n108), .Z(\ab[21][6] ) );
  AN2P U2645 ( .A(n319), .B(n108), .Z(\ab[21][5] ) );
  AN2P U2646 ( .A(n315), .B(n108), .Z(\ab[21][4] ) );
  AN2P U2647 ( .A(n311), .B(n108), .Z(\ab[21][3] ) );
  AN2P U2648 ( .A(n307), .B(n108), .Z(\ab[21][2] ) );
  AN2P U2649 ( .A(n303), .B(n108), .Z(\ab[21][1] ) );
  AN2P U2650 ( .A(n299), .B(n108), .Z(\ab[21][0] ) );
  AN2P U2651 ( .A(n451), .B(n93), .Z(\ab[22][38] ) );
  AN2P U2652 ( .A(n447), .B(n93), .Z(\ab[22][37] ) );
  AN2P U2653 ( .A(n443), .B(n93), .Z(\ab[22][36] ) );
  AN2P U2654 ( .A(n439), .B(n93), .Z(\ab[22][35] ) );
  AN2P U2655 ( .A(n435), .B(n93), .Z(\ab[22][34] ) );
  AN2P U2656 ( .A(n431), .B(n93), .Z(\ab[22][33] ) );
  AN2P U2657 ( .A(n427), .B(n93), .Z(\ab[22][32] ) );
  AN2P U2658 ( .A(n423), .B(n93), .Z(\ab[22][31] ) );
  AN2P U2659 ( .A(n419), .B(n94), .Z(\ab[22][30] ) );
  AN2P U2660 ( .A(n415), .B(n94), .Z(\ab[22][29] ) );
  AN2P U2661 ( .A(n411), .B(n94), .Z(\ab[22][28] ) );
  AN2P U2662 ( .A(n407), .B(n94), .Z(\ab[22][27] ) );
  AN2P U2663 ( .A(n403), .B(n94), .Z(\ab[22][26] ) );
  AN2P U2664 ( .A(n399), .B(n94), .Z(\ab[22][25] ) );
  AN2P U2665 ( .A(n395), .B(n94), .Z(\ab[22][24] ) );
  AN2P U2666 ( .A(n391), .B(n94), .Z(\ab[22][23] ) );
  AN2P U2667 ( .A(n387), .B(n95), .Z(\ab[22][22] ) );
  AN2P U2668 ( .A(n383), .B(n95), .Z(\ab[22][21] ) );
  AN2P U2669 ( .A(n379), .B(n95), .Z(\ab[22][20] ) );
  AN2P U2670 ( .A(n375), .B(n95), .Z(\ab[22][19] ) );
  AN2P U2671 ( .A(n371), .B(n95), .Z(\ab[22][18] ) );
  AN2P U2672 ( .A(n367), .B(n95), .Z(\ab[22][17] ) );
  AN2P U2673 ( .A(n363), .B(n95), .Z(\ab[22][16] ) );
  AN2P U2674 ( .A(n359), .B(n95), .Z(\ab[22][15] ) );
  AN2P U2675 ( .A(n355), .B(n96), .Z(\ab[22][14] ) );
  AN2P U2676 ( .A(n351), .B(n96), .Z(\ab[22][13] ) );
  AN2P U2677 ( .A(n347), .B(n96), .Z(\ab[22][12] ) );
  AN2P U2678 ( .A(n343), .B(n96), .Z(\ab[22][11] ) );
  AN2P U2679 ( .A(n339), .B(n96), .Z(\ab[22][10] ) );
  AN2P U2680 ( .A(n335), .B(n96), .Z(\ab[22][9] ) );
  AN2P U2681 ( .A(n331), .B(n96), .Z(\ab[22][8] ) );
  AN2P U2682 ( .A(n327), .B(n96), .Z(\ab[22][7] ) );
  AN2P U2683 ( .A(n323), .B(n97), .Z(\ab[22][6] ) );
  AN2P U2684 ( .A(n319), .B(n97), .Z(\ab[22][5] ) );
  AN2P U2685 ( .A(n315), .B(n97), .Z(\ab[22][4] ) );
  AN2P U2686 ( .A(n311), .B(n97), .Z(\ab[22][3] ) );
  AN2P U2687 ( .A(n307), .B(n97), .Z(\ab[22][2] ) );
  AN2P U2688 ( .A(n303), .B(n97), .Z(\ab[22][1] ) );
  AN2P U2689 ( .A(n299), .B(n97), .Z(\ab[22][0] ) );
  AN2P U2690 ( .A(n451), .B(n88), .Z(\ab[23][38] ) );
  AN2P U2691 ( .A(n447), .B(n88), .Z(\ab[23][37] ) );
  AN2P U2692 ( .A(n443), .B(n88), .Z(\ab[23][36] ) );
  AN2P U2693 ( .A(n439), .B(n88), .Z(\ab[23][35] ) );
  AN2P U2694 ( .A(n435), .B(n88), .Z(\ab[23][34] ) );
  AN2P U2695 ( .A(n431), .B(n88), .Z(\ab[23][33] ) );
  AN2P U2696 ( .A(n427), .B(n88), .Z(\ab[23][32] ) );
  AN2P U2697 ( .A(n423), .B(n88), .Z(\ab[23][31] ) );
  AN2P U2698 ( .A(n419), .B(n89), .Z(\ab[23][30] ) );
  AN2P U2699 ( .A(n415), .B(n89), .Z(\ab[23][29] ) );
  AN2P U2700 ( .A(n411), .B(n89), .Z(\ab[23][28] ) );
  AN2P U2701 ( .A(n407), .B(n89), .Z(\ab[23][27] ) );
  AN2P U2702 ( .A(n403), .B(n89), .Z(\ab[23][26] ) );
  AN2P U2703 ( .A(n399), .B(n89), .Z(\ab[23][25] ) );
  AN2P U2704 ( .A(n395), .B(n89), .Z(\ab[23][24] ) );
  AN2P U2705 ( .A(n391), .B(n89), .Z(\ab[23][23] ) );
  AN2P U2706 ( .A(n387), .B(n90), .Z(\ab[23][22] ) );
  AN2P U2707 ( .A(n383), .B(n90), .Z(\ab[23][21] ) );
  AN2P U2708 ( .A(n379), .B(n90), .Z(\ab[23][20] ) );
  AN2P U2709 ( .A(n375), .B(n90), .Z(\ab[23][19] ) );
  AN2P U2710 ( .A(n371), .B(n90), .Z(\ab[23][18] ) );
  AN2P U2711 ( .A(n367), .B(n90), .Z(\ab[23][17] ) );
  AN2P U2712 ( .A(n363), .B(n90), .Z(\ab[23][16] ) );
  AN2P U2713 ( .A(n359), .B(n90), .Z(\ab[23][15] ) );
  AN2P U2714 ( .A(n355), .B(n91), .Z(\ab[23][14] ) );
  AN2P U2715 ( .A(n351), .B(n91), .Z(\ab[23][13] ) );
  AN2P U2716 ( .A(n347), .B(n91), .Z(\ab[23][12] ) );
  AN2P U2717 ( .A(n343), .B(n91), .Z(\ab[23][11] ) );
  AN2P U2718 ( .A(n339), .B(n91), .Z(\ab[23][10] ) );
  AN2P U2719 ( .A(n335), .B(n91), .Z(\ab[23][9] ) );
  AN2P U2720 ( .A(n331), .B(n91), .Z(\ab[23][8] ) );
  AN2P U2721 ( .A(n327), .B(n91), .Z(\ab[23][7] ) );
  AN2P U2722 ( .A(n323), .B(n92), .Z(\ab[23][6] ) );
  AN2P U2723 ( .A(n319), .B(n92), .Z(\ab[23][5] ) );
  AN2P U2724 ( .A(n315), .B(n92), .Z(\ab[23][4] ) );
  AN2P U2725 ( .A(n311), .B(n92), .Z(\ab[23][3] ) );
  AN2P U2726 ( .A(n307), .B(n92), .Z(\ab[23][2] ) );
  AN2P U2727 ( .A(n303), .B(n92), .Z(\ab[23][1] ) );
  AN2P U2728 ( .A(n299), .B(n92), .Z(\ab[23][0] ) );
  AN2P U2729 ( .A(n451), .B(n77), .Z(\ab[24][38] ) );
  AN2P U2730 ( .A(n447), .B(n77), .Z(\ab[24][37] ) );
  AN2P U2731 ( .A(n443), .B(n77), .Z(\ab[24][36] ) );
  AN2P U2732 ( .A(n439), .B(n77), .Z(\ab[24][35] ) );
  AN2P U2733 ( .A(n435), .B(n77), .Z(\ab[24][34] ) );
  AN2P U2734 ( .A(n431), .B(n77), .Z(\ab[24][33] ) );
  AN2P U2735 ( .A(n427), .B(n77), .Z(\ab[24][32] ) );
  AN2P U2736 ( .A(n423), .B(n77), .Z(\ab[24][31] ) );
  AN2P U2737 ( .A(n419), .B(n78), .Z(\ab[24][30] ) );
  AN2P U2738 ( .A(n415), .B(n78), .Z(\ab[24][29] ) );
  AN2P U2739 ( .A(n411), .B(n78), .Z(\ab[24][28] ) );
  AN2P U2740 ( .A(n407), .B(n78), .Z(\ab[24][27] ) );
  AN2P U2741 ( .A(n403), .B(n78), .Z(\ab[24][26] ) );
  AN2P U2742 ( .A(n399), .B(n78), .Z(\ab[24][25] ) );
  AN2P U2743 ( .A(n395), .B(n78), .Z(\ab[24][24] ) );
  AN2P U2744 ( .A(n391), .B(n78), .Z(\ab[24][23] ) );
  AN2P U2745 ( .A(n387), .B(n79), .Z(\ab[24][22] ) );
  AN2P U2746 ( .A(n383), .B(n79), .Z(\ab[24][21] ) );
  AN2P U2747 ( .A(n379), .B(n79), .Z(\ab[24][20] ) );
  AN2P U2748 ( .A(n375), .B(n79), .Z(\ab[24][19] ) );
  AN2P U2749 ( .A(n371), .B(n79), .Z(\ab[24][18] ) );
  AN2P U2750 ( .A(n367), .B(n79), .Z(\ab[24][17] ) );
  AN2P U2751 ( .A(n363), .B(n79), .Z(\ab[24][16] ) );
  AN2P U2752 ( .A(n359), .B(n79), .Z(\ab[24][15] ) );
  AN2P U2753 ( .A(n355), .B(n80), .Z(\ab[24][14] ) );
  AN2P U2754 ( .A(n351), .B(n80), .Z(\ab[24][13] ) );
  AN2P U2755 ( .A(n347), .B(n80), .Z(\ab[24][12] ) );
  AN2P U2756 ( .A(n343), .B(n80), .Z(\ab[24][11] ) );
  AN2P U2757 ( .A(n339), .B(n80), .Z(\ab[24][10] ) );
  AN2P U2758 ( .A(n335), .B(n80), .Z(\ab[24][9] ) );
  AN2P U2759 ( .A(n331), .B(n80), .Z(\ab[24][8] ) );
  AN2P U2760 ( .A(n327), .B(n80), .Z(\ab[24][7] ) );
  AN2P U2761 ( .A(n323), .B(n81), .Z(\ab[24][6] ) );
  AN2P U2762 ( .A(n319), .B(n81), .Z(\ab[24][5] ) );
  AN2P U2763 ( .A(n315), .B(n81), .Z(\ab[24][4] ) );
  AN2P U2764 ( .A(n311), .B(n81), .Z(\ab[24][3] ) );
  AN2P U2765 ( .A(n307), .B(n81), .Z(\ab[24][2] ) );
  AN2P U2766 ( .A(n303), .B(n81), .Z(\ab[24][1] ) );
  AN2P U2767 ( .A(n299), .B(n81), .Z(\ab[24][0] ) );
  AN2P U2768 ( .A(n451), .B(n66), .Z(\ab[25][38] ) );
  AN2P U2769 ( .A(n447), .B(n66), .Z(\ab[25][37] ) );
  AN2P U2770 ( .A(n443), .B(n66), .Z(\ab[25][36] ) );
  AN2P U2771 ( .A(n439), .B(n66), .Z(\ab[25][35] ) );
  AN2P U2772 ( .A(n435), .B(n66), .Z(\ab[25][34] ) );
  AN2P U2773 ( .A(n431), .B(n66), .Z(\ab[25][33] ) );
  AN2P U2774 ( .A(n427), .B(n66), .Z(\ab[25][32] ) );
  AN2P U2775 ( .A(n423), .B(n66), .Z(\ab[25][31] ) );
  AN2P U2776 ( .A(n419), .B(n67), .Z(\ab[25][30] ) );
  AN2P U2777 ( .A(n415), .B(n67), .Z(\ab[25][29] ) );
  AN2P U2778 ( .A(n411), .B(n67), .Z(\ab[25][28] ) );
  AN2P U2779 ( .A(n407), .B(n67), .Z(\ab[25][27] ) );
  AN2P U2780 ( .A(n403), .B(n67), .Z(\ab[25][26] ) );
  AN2P U2781 ( .A(n399), .B(n67), .Z(\ab[25][25] ) );
  AN2P U2782 ( .A(n395), .B(n67), .Z(\ab[25][24] ) );
  AN2P U2783 ( .A(n391), .B(n67), .Z(\ab[25][23] ) );
  AN2P U2784 ( .A(n387), .B(n68), .Z(\ab[25][22] ) );
  AN2P U2785 ( .A(n383), .B(n68), .Z(\ab[25][21] ) );
  AN2P U2786 ( .A(n379), .B(n68), .Z(\ab[25][20] ) );
  AN2P U2787 ( .A(n375), .B(n68), .Z(\ab[25][19] ) );
  AN2P U2788 ( .A(n371), .B(n68), .Z(\ab[25][18] ) );
  AN2P U2789 ( .A(n367), .B(n68), .Z(\ab[25][17] ) );
  AN2P U2790 ( .A(n363), .B(n68), .Z(\ab[25][16] ) );
  AN2P U2791 ( .A(n359), .B(n68), .Z(\ab[25][15] ) );
  AN2P U2792 ( .A(n355), .B(n69), .Z(\ab[25][14] ) );
  AN2P U2793 ( .A(n351), .B(n69), .Z(\ab[25][13] ) );
  AN2P U2794 ( .A(n347), .B(n69), .Z(\ab[25][12] ) );
  AN2P U2795 ( .A(n343), .B(n69), .Z(\ab[25][11] ) );
  AN2P U2796 ( .A(n339), .B(n69), .Z(\ab[25][10] ) );
  AN2P U2797 ( .A(n335), .B(n69), .Z(\ab[25][9] ) );
  AN2P U2798 ( .A(n331), .B(n69), .Z(\ab[25][8] ) );
  AN2P U2799 ( .A(n327), .B(n69), .Z(\ab[25][7] ) );
  AN2P U2800 ( .A(n323), .B(n70), .Z(\ab[25][6] ) );
  AN2P U2801 ( .A(n319), .B(n70), .Z(\ab[25][5] ) );
  AN2P U2802 ( .A(n315), .B(n70), .Z(\ab[25][4] ) );
  AN2P U2803 ( .A(n311), .B(n70), .Z(\ab[25][3] ) );
  AN2P U2804 ( .A(n307), .B(n70), .Z(\ab[25][2] ) );
  AN2P U2805 ( .A(n303), .B(n70), .Z(\ab[25][1] ) );
  AN2P U2806 ( .A(n299), .B(n70), .Z(\ab[25][0] ) );
  AN2P U2807 ( .A(n451), .B(n55), .Z(\ab[26][38] ) );
  AN2P U2808 ( .A(n447), .B(n55), .Z(\ab[26][37] ) );
  AN2P U2809 ( .A(n443), .B(n55), .Z(\ab[26][36] ) );
  AN2P U2810 ( .A(n439), .B(n55), .Z(\ab[26][35] ) );
  AN2P U2811 ( .A(n435), .B(n55), .Z(\ab[26][34] ) );
  AN2P U2812 ( .A(n431), .B(n55), .Z(\ab[26][33] ) );
  AN2P U2813 ( .A(n427), .B(n55), .Z(\ab[26][32] ) );
  AN2P U2814 ( .A(n423), .B(n55), .Z(\ab[26][31] ) );
  AN2P U2815 ( .A(n419), .B(n56), .Z(\ab[26][30] ) );
  AN2P U2816 ( .A(n415), .B(n56), .Z(\ab[26][29] ) );
  AN2P U2817 ( .A(n411), .B(n56), .Z(\ab[26][28] ) );
  AN2P U2818 ( .A(n407), .B(n56), .Z(\ab[26][27] ) );
  AN2P U2819 ( .A(n403), .B(n56), .Z(\ab[26][26] ) );
  AN2P U2820 ( .A(n399), .B(n56), .Z(\ab[26][25] ) );
  AN2P U2821 ( .A(n395), .B(n56), .Z(\ab[26][24] ) );
  AN2P U2822 ( .A(n391), .B(n56), .Z(\ab[26][23] ) );
  AN2P U2823 ( .A(n387), .B(n57), .Z(\ab[26][22] ) );
  AN2P U2824 ( .A(n383), .B(n57), .Z(\ab[26][21] ) );
  AN2P U2825 ( .A(n379), .B(n57), .Z(\ab[26][20] ) );
  AN2P U2826 ( .A(n375), .B(n57), .Z(\ab[26][19] ) );
  AN2P U2827 ( .A(n371), .B(n57), .Z(\ab[26][18] ) );
  AN2P U2828 ( .A(n367), .B(n57), .Z(\ab[26][17] ) );
  AN2P U2829 ( .A(n363), .B(n57), .Z(\ab[26][16] ) );
  AN2P U2830 ( .A(n359), .B(n57), .Z(\ab[26][15] ) );
  AN2P U2831 ( .A(n355), .B(n58), .Z(\ab[26][14] ) );
  AN2P U2832 ( .A(n351), .B(n58), .Z(\ab[26][13] ) );
  AN2P U2833 ( .A(n347), .B(n58), .Z(\ab[26][12] ) );
  AN2P U2834 ( .A(n343), .B(n58), .Z(\ab[26][11] ) );
  AN2P U2835 ( .A(n339), .B(n58), .Z(\ab[26][10] ) );
  AN2P U2836 ( .A(n335), .B(n58), .Z(\ab[26][9] ) );
  AN2P U2837 ( .A(n331), .B(n58), .Z(\ab[26][8] ) );
  AN2P U2838 ( .A(n327), .B(n58), .Z(\ab[26][7] ) );
  AN2P U2839 ( .A(n323), .B(n59), .Z(\ab[26][6] ) );
  AN2P U2840 ( .A(n319), .B(n59), .Z(\ab[26][5] ) );
  AN2P U2841 ( .A(n315), .B(n59), .Z(\ab[26][4] ) );
  AN2P U2842 ( .A(n311), .B(n59), .Z(\ab[26][3] ) );
  AN2P U2843 ( .A(n307), .B(n59), .Z(\ab[26][2] ) );
  AN2P U2844 ( .A(n303), .B(n59), .Z(\ab[26][1] ) );
  AN2P U2845 ( .A(n299), .B(n59), .Z(\ab[26][0] ) );
  AN2P U2846 ( .A(n451), .B(n44), .Z(\ab[27][38] ) );
  AN2P U2847 ( .A(n447), .B(n44), .Z(\ab[27][37] ) );
  AN2P U2848 ( .A(n443), .B(n44), .Z(\ab[27][36] ) );
  AN2P U2849 ( .A(n439), .B(n44), .Z(\ab[27][35] ) );
  AN2P U2850 ( .A(n435), .B(n44), .Z(\ab[27][34] ) );
  AN2P U2851 ( .A(n431), .B(n44), .Z(\ab[27][33] ) );
  AN2P U2852 ( .A(n427), .B(n44), .Z(\ab[27][32] ) );
  AN2P U2853 ( .A(n423), .B(n44), .Z(\ab[27][31] ) );
  AN2P U2854 ( .A(n419), .B(n45), .Z(\ab[27][30] ) );
  AN2P U2855 ( .A(n415), .B(n45), .Z(\ab[27][29] ) );
  AN2P U2856 ( .A(n411), .B(n45), .Z(\ab[27][28] ) );
  AN2P U2857 ( .A(n407), .B(n45), .Z(\ab[27][27] ) );
  AN2P U2858 ( .A(n403), .B(n45), .Z(\ab[27][26] ) );
  AN2P U2859 ( .A(n399), .B(n45), .Z(\ab[27][25] ) );
  AN2P U2860 ( .A(n395), .B(n45), .Z(\ab[27][24] ) );
  AN2P U2861 ( .A(n391), .B(n45), .Z(\ab[27][23] ) );
  AN2P U2862 ( .A(n387), .B(n46), .Z(\ab[27][22] ) );
  AN2P U2863 ( .A(n383), .B(n46), .Z(\ab[27][21] ) );
  AN2P U2864 ( .A(n379), .B(n46), .Z(\ab[27][20] ) );
  AN2P U2865 ( .A(n375), .B(n46), .Z(\ab[27][19] ) );
  AN2P U2866 ( .A(n371), .B(n46), .Z(\ab[27][18] ) );
  AN2P U2867 ( .A(n367), .B(n46), .Z(\ab[27][17] ) );
  AN2P U2868 ( .A(n363), .B(n46), .Z(\ab[27][16] ) );
  AN2P U2869 ( .A(n359), .B(n46), .Z(\ab[27][15] ) );
  AN2P U2870 ( .A(n355), .B(n47), .Z(\ab[27][14] ) );
  AN2P U2871 ( .A(n351), .B(n47), .Z(\ab[27][13] ) );
  AN2P U2872 ( .A(n347), .B(n47), .Z(\ab[27][12] ) );
  AN2P U2873 ( .A(n343), .B(n47), .Z(\ab[27][11] ) );
  AN2P U2874 ( .A(n339), .B(n47), .Z(\ab[27][10] ) );
  AN2P U2875 ( .A(n335), .B(n47), .Z(\ab[27][9] ) );
  AN2P U2876 ( .A(n331), .B(n47), .Z(\ab[27][8] ) );
  AN2P U2877 ( .A(n327), .B(n47), .Z(\ab[27][7] ) );
  AN2P U2878 ( .A(n323), .B(n48), .Z(\ab[27][6] ) );
  AN2P U2879 ( .A(n319), .B(n48), .Z(\ab[27][5] ) );
  AN2P U2880 ( .A(n315), .B(n48), .Z(\ab[27][4] ) );
  AN2P U2881 ( .A(n311), .B(n48), .Z(\ab[27][3] ) );
  AN2P U2882 ( .A(n307), .B(n48), .Z(\ab[27][2] ) );
  AN2P U2883 ( .A(n303), .B(n48), .Z(\ab[27][1] ) );
  AN2P U2884 ( .A(n299), .B(n48), .Z(\ab[27][0] ) );
  AN2P U2885 ( .A(n451), .B(n33), .Z(\ab[28][38] ) );
  AN2P U2886 ( .A(n447), .B(n33), .Z(\ab[28][37] ) );
  AN2P U2887 ( .A(n443), .B(n33), .Z(\ab[28][36] ) );
  AN2P U2888 ( .A(n439), .B(n33), .Z(\ab[28][35] ) );
  AN2P U2889 ( .A(n435), .B(n33), .Z(\ab[28][34] ) );
  AN2P U2890 ( .A(n431), .B(n33), .Z(\ab[28][33] ) );
  AN2P U2891 ( .A(n427), .B(n33), .Z(\ab[28][32] ) );
  AN2P U2892 ( .A(n423), .B(n33), .Z(\ab[28][31] ) );
  AN2P U2893 ( .A(n419), .B(n34), .Z(\ab[28][30] ) );
  AN2P U2894 ( .A(n415), .B(n34), .Z(\ab[28][29] ) );
  AN2P U2895 ( .A(n411), .B(n34), .Z(\ab[28][28] ) );
  AN2P U2896 ( .A(n407), .B(n34), .Z(\ab[28][27] ) );
  AN2P U2897 ( .A(n403), .B(n34), .Z(\ab[28][26] ) );
  AN2P U2898 ( .A(n399), .B(n34), .Z(\ab[28][25] ) );
  AN2P U2899 ( .A(n395), .B(n34), .Z(\ab[28][24] ) );
  AN2P U2900 ( .A(n391), .B(n34), .Z(\ab[28][23] ) );
  AN2P U2901 ( .A(n387), .B(n35), .Z(\ab[28][22] ) );
  AN2P U2902 ( .A(n383), .B(n35), .Z(\ab[28][21] ) );
  AN2P U2903 ( .A(n379), .B(n35), .Z(\ab[28][20] ) );
  AN2P U2904 ( .A(n375), .B(n35), .Z(\ab[28][19] ) );
  AN2P U2905 ( .A(n371), .B(n35), .Z(\ab[28][18] ) );
  AN2P U2906 ( .A(n367), .B(n35), .Z(\ab[28][17] ) );
  AN2P U2907 ( .A(n363), .B(n35), .Z(\ab[28][16] ) );
  AN2P U2908 ( .A(n359), .B(n35), .Z(\ab[28][15] ) );
  AN2P U2909 ( .A(n355), .B(n36), .Z(\ab[28][14] ) );
  AN2P U2910 ( .A(n351), .B(n36), .Z(\ab[28][13] ) );
  AN2P U2911 ( .A(n347), .B(n36), .Z(\ab[28][12] ) );
  AN2P U2912 ( .A(n343), .B(n36), .Z(\ab[28][11] ) );
  AN2P U2913 ( .A(n339), .B(n36), .Z(\ab[28][10] ) );
  AN2P U2914 ( .A(n335), .B(n36), .Z(\ab[28][9] ) );
  AN2P U2915 ( .A(n331), .B(n36), .Z(\ab[28][8] ) );
  AN2P U2916 ( .A(n327), .B(n36), .Z(\ab[28][7] ) );
  AN2P U2917 ( .A(n323), .B(n37), .Z(\ab[28][6] ) );
  AN2P U2918 ( .A(n319), .B(n37), .Z(\ab[28][5] ) );
  AN2P U2919 ( .A(n315), .B(n37), .Z(\ab[28][4] ) );
  AN2P U2920 ( .A(n311), .B(n37), .Z(\ab[28][3] ) );
  AN2P U2921 ( .A(n307), .B(n37), .Z(\ab[28][2] ) );
  AN2P U2922 ( .A(n303), .B(n37), .Z(\ab[28][1] ) );
  AN2P U2923 ( .A(n299), .B(n37), .Z(\ab[28][0] ) );
  AN2P U2924 ( .A(n451), .B(n22), .Z(\ab[29][38] ) );
  AN2P U2925 ( .A(n447), .B(n22), .Z(\ab[29][37] ) );
  AN2P U2926 ( .A(n443), .B(n22), .Z(\ab[29][36] ) );
  AN2P U2927 ( .A(n439), .B(n22), .Z(\ab[29][35] ) );
  AN2P U2928 ( .A(n435), .B(n22), .Z(\ab[29][34] ) );
  AN2P U2929 ( .A(n431), .B(n22), .Z(\ab[29][33] ) );
  AN2P U2930 ( .A(n427), .B(n22), .Z(\ab[29][32] ) );
  AN2P U2931 ( .A(n423), .B(n22), .Z(\ab[29][31] ) );
  AN2P U2932 ( .A(n419), .B(n23), .Z(\ab[29][30] ) );
  AN2P U2933 ( .A(n415), .B(n23), .Z(\ab[29][29] ) );
  AN2P U2934 ( .A(n411), .B(n23), .Z(\ab[29][28] ) );
  AN2P U2935 ( .A(n407), .B(n23), .Z(\ab[29][27] ) );
  AN2P U2936 ( .A(n403), .B(n23), .Z(\ab[29][26] ) );
  AN2P U2937 ( .A(n399), .B(n23), .Z(\ab[29][25] ) );
  AN2P U2938 ( .A(n395), .B(n23), .Z(\ab[29][24] ) );
  AN2P U2939 ( .A(n391), .B(n23), .Z(\ab[29][23] ) );
  AN2P U2940 ( .A(n387), .B(n24), .Z(\ab[29][22] ) );
  AN2P U2941 ( .A(n383), .B(n24), .Z(\ab[29][21] ) );
  AN2P U2942 ( .A(n379), .B(n24), .Z(\ab[29][20] ) );
  AN2P U2943 ( .A(n375), .B(n24), .Z(\ab[29][19] ) );
  AN2P U2944 ( .A(n371), .B(n24), .Z(\ab[29][18] ) );
  AN2P U2945 ( .A(n367), .B(n24), .Z(\ab[29][17] ) );
  AN2P U2946 ( .A(n363), .B(n24), .Z(\ab[29][16] ) );
  AN2P U2947 ( .A(n359), .B(n24), .Z(\ab[29][15] ) );
  AN2P U2948 ( .A(n355), .B(n25), .Z(\ab[29][14] ) );
  AN2P U2949 ( .A(n351), .B(n25), .Z(\ab[29][13] ) );
  AN2P U2950 ( .A(n347), .B(n25), .Z(\ab[29][12] ) );
  AN2P U2951 ( .A(n343), .B(n25), .Z(\ab[29][11] ) );
  AN2P U2952 ( .A(n339), .B(n25), .Z(\ab[29][10] ) );
  AN2P U2953 ( .A(n335), .B(n25), .Z(\ab[29][9] ) );
  AN2P U2954 ( .A(n331), .B(n25), .Z(\ab[29][8] ) );
  AN2P U2955 ( .A(n327), .B(n25), .Z(\ab[29][7] ) );
  AN2P U2956 ( .A(n323), .B(n26), .Z(\ab[29][6] ) );
  AN2P U2957 ( .A(n319), .B(n26), .Z(\ab[29][5] ) );
  AN2P U2958 ( .A(n315), .B(n26), .Z(\ab[29][4] ) );
  AN2P U2959 ( .A(n311), .B(n26), .Z(\ab[29][3] ) );
  AN2P U2960 ( .A(n307), .B(n26), .Z(\ab[29][2] ) );
  AN2P U2961 ( .A(n303), .B(n26), .Z(\ab[29][1] ) );
  AN2P U2962 ( .A(n299), .B(n26), .Z(\ab[29][0] ) );
  NR2 U2964 ( .A(n492), .B(n16), .Z(\ab[29][95] ) );
  NR2 U2965 ( .A(n493), .B(n16), .Z(\ab[29][94] ) );
  NR2 U2966 ( .A(n494), .B(n16), .Z(\ab[29][93] ) );
  NR2 U2967 ( .A(n495), .B(n16), .Z(\ab[29][92] ) );
  NR2 U2968 ( .A(n496), .B(n16), .Z(\ab[29][91] ) );
  NR2 U2969 ( .A(n497), .B(n16), .Z(\ab[29][90] ) );
  NR2 U2970 ( .A(n498), .B(n16), .Z(\ab[29][89] ) );
  NR2 U2971 ( .A(n499), .B(n16), .Z(\ab[29][88] ) );
  NR2 U2972 ( .A(n500), .B(n16), .Z(\ab[29][87] ) );
  NR2 U2973 ( .A(n501), .B(n16), .Z(\ab[29][86] ) );
  NR2 U2974 ( .A(n502), .B(n16), .Z(\ab[29][85] ) );
  NR2 U2975 ( .A(n503), .B(n16), .Z(\ab[29][84] ) );
  NR2 U2976 ( .A(n504), .B(n17), .Z(\ab[29][83] ) );
  NR2 U2977 ( .A(n505), .B(n17), .Z(\ab[29][82] ) );
  NR2 U2978 ( .A(n506), .B(n17), .Z(\ab[29][81] ) );
  NR2 U2979 ( .A(n507), .B(n17), .Z(\ab[29][80] ) );
  NR2 U2980 ( .A(n508), .B(n17), .Z(\ab[29][79] ) );
  NR2 U2981 ( .A(n509), .B(n17), .Z(\ab[29][78] ) );
  NR2 U2982 ( .A(n510), .B(n17), .Z(\ab[29][77] ) );
  NR2 U2983 ( .A(n511), .B(n17), .Z(\ab[29][76] ) );
  NR2 U2984 ( .A(n512), .B(n17), .Z(\ab[29][75] ) );
  NR2 U2985 ( .A(n513), .B(n17), .Z(\ab[29][74] ) );
  NR2 U2986 ( .A(n514), .B(n17), .Z(\ab[29][73] ) );
  NR2 U2987 ( .A(n515), .B(n17), .Z(\ab[29][72] ) );
  NR2 U2988 ( .A(n516), .B(n18), .Z(\ab[29][71] ) );
  NR2 U2989 ( .A(n517), .B(n18), .Z(\ab[29][70] ) );
  NR2 U2990 ( .A(n518), .B(n18), .Z(\ab[29][69] ) );
  NR2 U2991 ( .A(n519), .B(n18), .Z(\ab[29][68] ) );
  NR2 U2992 ( .A(n520), .B(n18), .Z(\ab[29][67] ) );
  NR2 U2993 ( .A(n521), .B(n18), .Z(\ab[29][66] ) );
  NR2 U2994 ( .A(n522), .B(n18), .Z(\ab[29][65] ) );
  NR2 U2995 ( .A(n523), .B(n18), .Z(\ab[29][64] ) );
  NR2 U2996 ( .A(n524), .B(n18), .Z(\ab[29][63] ) );
  NR2 U2997 ( .A(n525), .B(n18), .Z(\ab[29][62] ) );
  NR2 U2998 ( .A(n526), .B(n18), .Z(\ab[29][61] ) );
  NR2 U2999 ( .A(n527), .B(n18), .Z(\ab[29][60] ) );
  NR2 U3000 ( .A(n528), .B(n19), .Z(\ab[29][59] ) );
  NR2 U3001 ( .A(n529), .B(n19), .Z(\ab[29][58] ) );
  NR2 U3002 ( .A(n530), .B(n19), .Z(\ab[29][57] ) );
  NR2 U3003 ( .A(n531), .B(n19), .Z(\ab[29][56] ) );
  NR2 U3004 ( .A(n532), .B(n19), .Z(\ab[29][55] ) );
  NR2 U3005 ( .A(n533), .B(n19), .Z(\ab[29][54] ) );
  NR2 U3006 ( .A(n534), .B(n19), .Z(\ab[29][53] ) );
  NR2 U3007 ( .A(n535), .B(n19), .Z(\ab[29][52] ) );
  NR2 U3008 ( .A(n536), .B(n19), .Z(\ab[29][51] ) );
  NR2 U3009 ( .A(n537), .B(n19), .Z(\ab[29][50] ) );
  NR2 U3010 ( .A(n538), .B(n19), .Z(\ab[29][49] ) );
  NR2 U3011 ( .A(n539), .B(n19), .Z(\ab[29][48] ) );
  NR2 U3012 ( .A(n540), .B(n20), .Z(\ab[29][47] ) );
  NR2 U3013 ( .A(n541), .B(n20), .Z(\ab[29][46] ) );
  NR2 U3014 ( .A(n542), .B(n20), .Z(\ab[29][45] ) );
  NR2 U3015 ( .A(n543), .B(n20), .Z(\ab[29][44] ) );
  NR2 U3016 ( .A(n544), .B(n20), .Z(\ab[29][43] ) );
  NR2 U3017 ( .A(n545), .B(n20), .Z(\ab[29][42] ) );
  NR2 U3018 ( .A(n546), .B(n20), .Z(\ab[29][41] ) );
  NR2 U3019 ( .A(n547), .B(n20), .Z(\ab[29][40] ) );
  NR2 U3020 ( .A(n548), .B(n20), .Z(\ab[29][39] ) );
  NR2 U3021 ( .A(n492), .B(n27), .Z(\ab[28][95] ) );
  NR2 U3022 ( .A(n493), .B(n27), .Z(\ab[28][94] ) );
  NR2 U3023 ( .A(n494), .B(n27), .Z(\ab[28][93] ) );
  NR2 U3024 ( .A(n495), .B(n27), .Z(\ab[28][92] ) );
  NR2 U3025 ( .A(n496), .B(n27), .Z(\ab[28][91] ) );
  NR2 U3026 ( .A(n497), .B(n27), .Z(\ab[28][90] ) );
  NR2 U3027 ( .A(n498), .B(n27), .Z(\ab[28][89] ) );
  NR2 U3028 ( .A(n499), .B(n27), .Z(\ab[28][88] ) );
  NR2 U3029 ( .A(n500), .B(n27), .Z(\ab[28][87] ) );
  NR2 U3030 ( .A(n501), .B(n27), .Z(\ab[28][86] ) );
  NR2 U3031 ( .A(n502), .B(n27), .Z(\ab[28][85] ) );
  NR2 U3032 ( .A(n503), .B(n27), .Z(\ab[28][84] ) );
  NR2 U3033 ( .A(n504), .B(n28), .Z(\ab[28][83] ) );
  NR2 U3034 ( .A(n505), .B(n28), .Z(\ab[28][82] ) );
  NR2 U3035 ( .A(n506), .B(n28), .Z(\ab[28][81] ) );
  NR2 U3036 ( .A(n507), .B(n28), .Z(\ab[28][80] ) );
  NR2 U3037 ( .A(n508), .B(n28), .Z(\ab[28][79] ) );
  NR2 U3038 ( .A(n509), .B(n28), .Z(\ab[28][78] ) );
  NR2 U3039 ( .A(n510), .B(n28), .Z(\ab[28][77] ) );
  NR2 U3040 ( .A(n511), .B(n28), .Z(\ab[28][76] ) );
  NR2 U3041 ( .A(n512), .B(n28), .Z(\ab[28][75] ) );
  NR2 U3042 ( .A(n513), .B(n28), .Z(\ab[28][74] ) );
  NR2 U3043 ( .A(n514), .B(n28), .Z(\ab[28][73] ) );
  NR2 U3044 ( .A(n515), .B(n28), .Z(\ab[28][72] ) );
  NR2 U3045 ( .A(n516), .B(n29), .Z(\ab[28][71] ) );
  NR2 U3046 ( .A(n517), .B(n29), .Z(\ab[28][70] ) );
  NR2 U3047 ( .A(n518), .B(n29), .Z(\ab[28][69] ) );
  NR2 U3048 ( .A(n519), .B(n29), .Z(\ab[28][68] ) );
  NR2 U3049 ( .A(n520), .B(n29), .Z(\ab[28][67] ) );
  NR2 U3050 ( .A(n521), .B(n29), .Z(\ab[28][66] ) );
  NR2 U3051 ( .A(n522), .B(n29), .Z(\ab[28][65] ) );
  NR2 U3052 ( .A(n523), .B(n29), .Z(\ab[28][64] ) );
  NR2 U3053 ( .A(n524), .B(n29), .Z(\ab[28][63] ) );
  NR2 U3054 ( .A(n525), .B(n29), .Z(\ab[28][62] ) );
  NR2 U3055 ( .A(n526), .B(n29), .Z(\ab[28][61] ) );
  NR2 U3056 ( .A(n527), .B(n29), .Z(\ab[28][60] ) );
  NR2 U3057 ( .A(n528), .B(n30), .Z(\ab[28][59] ) );
  NR2 U3058 ( .A(n529), .B(n30), .Z(\ab[28][58] ) );
  NR2 U3059 ( .A(n530), .B(n30), .Z(\ab[28][57] ) );
  NR2 U3060 ( .A(n531), .B(n30), .Z(\ab[28][56] ) );
  NR2 U3061 ( .A(n532), .B(n30), .Z(\ab[28][55] ) );
  NR2 U3062 ( .A(n533), .B(n30), .Z(\ab[28][54] ) );
  NR2 U3063 ( .A(n534), .B(n30), .Z(\ab[28][53] ) );
  NR2 U3064 ( .A(n535), .B(n30), .Z(\ab[28][52] ) );
  NR2 U3065 ( .A(n536), .B(n30), .Z(\ab[28][51] ) );
  NR2 U3066 ( .A(n537), .B(n30), .Z(\ab[28][50] ) );
  NR2 U3067 ( .A(n538), .B(n30), .Z(\ab[28][49] ) );
  NR2 U3068 ( .A(n539), .B(n30), .Z(\ab[28][48] ) );
  NR2 U3069 ( .A(n540), .B(n31), .Z(\ab[28][47] ) );
  NR2 U3070 ( .A(n541), .B(n31), .Z(\ab[28][46] ) );
  NR2 U3071 ( .A(n542), .B(n31), .Z(\ab[28][45] ) );
  NR2 U3072 ( .A(n543), .B(n31), .Z(\ab[28][44] ) );
  NR2 U3073 ( .A(n544), .B(n31), .Z(\ab[28][43] ) );
  NR2 U3074 ( .A(n545), .B(n31), .Z(\ab[28][42] ) );
  NR2 U3075 ( .A(n546), .B(n31), .Z(\ab[28][41] ) );
  NR2 U3076 ( .A(n547), .B(n31), .Z(\ab[28][40] ) );
  NR2 U3077 ( .A(n548), .B(n31), .Z(\ab[28][39] ) );
  NR2 U3078 ( .A(n492), .B(n38), .Z(\ab[27][95] ) );
  NR2 U3079 ( .A(n493), .B(n38), .Z(\ab[27][94] ) );
  NR2 U3080 ( .A(n494), .B(n38), .Z(\ab[27][93] ) );
  NR2 U3081 ( .A(n495), .B(n38), .Z(\ab[27][92] ) );
  NR2 U3082 ( .A(n496), .B(n38), .Z(\ab[27][91] ) );
  NR2 U3083 ( .A(n497), .B(n38), .Z(\ab[27][90] ) );
  NR2 U3084 ( .A(n498), .B(n38), .Z(\ab[27][89] ) );
  NR2 U3085 ( .A(n499), .B(n38), .Z(\ab[27][88] ) );
  NR2 U3086 ( .A(n500), .B(n38), .Z(\ab[27][87] ) );
  NR2 U3087 ( .A(n501), .B(n38), .Z(\ab[27][86] ) );
  NR2 U3088 ( .A(n502), .B(n38), .Z(\ab[27][85] ) );
  NR2 U3089 ( .A(n503), .B(n38), .Z(\ab[27][84] ) );
  NR2 U3090 ( .A(n504), .B(n39), .Z(\ab[27][83] ) );
  NR2 U3091 ( .A(n505), .B(n39), .Z(\ab[27][82] ) );
  NR2 U3092 ( .A(n506), .B(n39), .Z(\ab[27][81] ) );
  NR2 U3093 ( .A(n507), .B(n39), .Z(\ab[27][80] ) );
  NR2 U3094 ( .A(n508), .B(n39), .Z(\ab[27][79] ) );
  NR2 U3095 ( .A(n509), .B(n39), .Z(\ab[27][78] ) );
  NR2 U3096 ( .A(n510), .B(n39), .Z(\ab[27][77] ) );
  NR2 U3097 ( .A(n511), .B(n39), .Z(\ab[27][76] ) );
  NR2 U3098 ( .A(n512), .B(n39), .Z(\ab[27][75] ) );
  NR2 U3099 ( .A(n513), .B(n39), .Z(\ab[27][74] ) );
  NR2 U3100 ( .A(n514), .B(n39), .Z(\ab[27][73] ) );
  NR2 U3101 ( .A(n515), .B(n39), .Z(\ab[27][72] ) );
  NR2 U3102 ( .A(n516), .B(n40), .Z(\ab[27][71] ) );
  NR2 U3103 ( .A(n517), .B(n40), .Z(\ab[27][70] ) );
  NR2 U3104 ( .A(n518), .B(n40), .Z(\ab[27][69] ) );
  NR2 U3105 ( .A(n519), .B(n40), .Z(\ab[27][68] ) );
  NR2 U3106 ( .A(n520), .B(n40), .Z(\ab[27][67] ) );
  NR2 U3107 ( .A(n521), .B(n40), .Z(\ab[27][66] ) );
  NR2 U3108 ( .A(n522), .B(n40), .Z(\ab[27][65] ) );
  NR2 U3109 ( .A(n523), .B(n40), .Z(\ab[27][64] ) );
  NR2 U3110 ( .A(n524), .B(n40), .Z(\ab[27][63] ) );
  NR2 U3111 ( .A(n525), .B(n40), .Z(\ab[27][62] ) );
  NR2 U3112 ( .A(n526), .B(n40), .Z(\ab[27][61] ) );
  NR2 U3113 ( .A(n527), .B(n40), .Z(\ab[27][60] ) );
  NR2 U3114 ( .A(n528), .B(n41), .Z(\ab[27][59] ) );
  NR2 U3115 ( .A(n529), .B(n41), .Z(\ab[27][58] ) );
  NR2 U3116 ( .A(n530), .B(n41), .Z(\ab[27][57] ) );
  NR2 U3117 ( .A(n531), .B(n41), .Z(\ab[27][56] ) );
  NR2 U3118 ( .A(n532), .B(n41), .Z(\ab[27][55] ) );
  NR2 U3119 ( .A(n533), .B(n41), .Z(\ab[27][54] ) );
  NR2 U3120 ( .A(n534), .B(n41), .Z(\ab[27][53] ) );
  NR2 U3121 ( .A(n535), .B(n41), .Z(\ab[27][52] ) );
  NR2 U3122 ( .A(n536), .B(n41), .Z(\ab[27][51] ) );
  NR2 U3123 ( .A(n537), .B(n41), .Z(\ab[27][50] ) );
  NR2 U3124 ( .A(n538), .B(n41), .Z(\ab[27][49] ) );
  NR2 U3125 ( .A(n539), .B(n41), .Z(\ab[27][48] ) );
  NR2 U3126 ( .A(n540), .B(n42), .Z(\ab[27][47] ) );
  NR2 U3127 ( .A(n541), .B(n42), .Z(\ab[27][46] ) );
  NR2 U3128 ( .A(n542), .B(n42), .Z(\ab[27][45] ) );
  NR2 U3129 ( .A(n543), .B(n42), .Z(\ab[27][44] ) );
  NR2 U3130 ( .A(n544), .B(n42), .Z(\ab[27][43] ) );
  NR2 U3131 ( .A(n545), .B(n42), .Z(\ab[27][42] ) );
  NR2 U3132 ( .A(n546), .B(n42), .Z(\ab[27][41] ) );
  NR2 U3133 ( .A(n547), .B(n42), .Z(\ab[27][40] ) );
  NR2 U3134 ( .A(n548), .B(n42), .Z(\ab[27][39] ) );
  NR2 U3135 ( .A(n492), .B(n49), .Z(\ab[26][95] ) );
  NR2 U3136 ( .A(n493), .B(n49), .Z(\ab[26][94] ) );
  NR2 U3137 ( .A(n494), .B(n49), .Z(\ab[26][93] ) );
  NR2 U3138 ( .A(n495), .B(n49), .Z(\ab[26][92] ) );
  NR2 U3139 ( .A(n496), .B(n49), .Z(\ab[26][91] ) );
  NR2 U3140 ( .A(n497), .B(n49), .Z(\ab[26][90] ) );
  NR2 U3141 ( .A(n498), .B(n49), .Z(\ab[26][89] ) );
  NR2 U3142 ( .A(n499), .B(n49), .Z(\ab[26][88] ) );
  NR2 U3143 ( .A(n500), .B(n49), .Z(\ab[26][87] ) );
  NR2 U3144 ( .A(n501), .B(n49), .Z(\ab[26][86] ) );
  NR2 U3145 ( .A(n502), .B(n49), .Z(\ab[26][85] ) );
  NR2 U3146 ( .A(n503), .B(n49), .Z(\ab[26][84] ) );
  NR2 U3147 ( .A(n504), .B(n50), .Z(\ab[26][83] ) );
  NR2 U3148 ( .A(n505), .B(n50), .Z(\ab[26][82] ) );
  NR2 U3149 ( .A(n506), .B(n50), .Z(\ab[26][81] ) );
  NR2 U3150 ( .A(n507), .B(n50), .Z(\ab[26][80] ) );
  NR2 U3151 ( .A(n508), .B(n50), .Z(\ab[26][79] ) );
  NR2 U3152 ( .A(n509), .B(n50), .Z(\ab[26][78] ) );
  NR2 U3153 ( .A(n510), .B(n50), .Z(\ab[26][77] ) );
  NR2 U3154 ( .A(n511), .B(n50), .Z(\ab[26][76] ) );
  NR2 U3155 ( .A(n512), .B(n50), .Z(\ab[26][75] ) );
  NR2 U3156 ( .A(n513), .B(n50), .Z(\ab[26][74] ) );
  NR2 U3157 ( .A(n514), .B(n50), .Z(\ab[26][73] ) );
  NR2 U3158 ( .A(n515), .B(n50), .Z(\ab[26][72] ) );
  NR2 U3159 ( .A(n516), .B(n51), .Z(\ab[26][71] ) );
  NR2 U3160 ( .A(n517), .B(n51), .Z(\ab[26][70] ) );
  NR2 U3161 ( .A(n518), .B(n51), .Z(\ab[26][69] ) );
  NR2 U3162 ( .A(n519), .B(n51), .Z(\ab[26][68] ) );
  NR2 U3163 ( .A(n520), .B(n51), .Z(\ab[26][67] ) );
  NR2 U3164 ( .A(n521), .B(n51), .Z(\ab[26][66] ) );
  NR2 U3165 ( .A(n522), .B(n51), .Z(\ab[26][65] ) );
  NR2 U3166 ( .A(n523), .B(n51), .Z(\ab[26][64] ) );
  NR2 U3167 ( .A(n524), .B(n51), .Z(\ab[26][63] ) );
  NR2 U3168 ( .A(n525), .B(n51), .Z(\ab[26][62] ) );
  NR2 U3169 ( .A(n526), .B(n51), .Z(\ab[26][61] ) );
  NR2 U3170 ( .A(n527), .B(n51), .Z(\ab[26][60] ) );
  NR2 U3171 ( .A(n528), .B(n52), .Z(\ab[26][59] ) );
  NR2 U3172 ( .A(n529), .B(n52), .Z(\ab[26][58] ) );
  NR2 U3173 ( .A(n530), .B(n52), .Z(\ab[26][57] ) );
  NR2 U3174 ( .A(n531), .B(n52), .Z(\ab[26][56] ) );
  NR2 U3175 ( .A(n532), .B(n52), .Z(\ab[26][55] ) );
  NR2 U3176 ( .A(n533), .B(n52), .Z(\ab[26][54] ) );
  NR2 U3177 ( .A(n534), .B(n52), .Z(\ab[26][53] ) );
  NR2 U3178 ( .A(n535), .B(n52), .Z(\ab[26][52] ) );
  NR2 U3179 ( .A(n536), .B(n52), .Z(\ab[26][51] ) );
  NR2 U3180 ( .A(n537), .B(n52), .Z(\ab[26][50] ) );
  NR2 U3181 ( .A(n538), .B(n52), .Z(\ab[26][49] ) );
  NR2 U3182 ( .A(n539), .B(n52), .Z(\ab[26][48] ) );
  NR2 U3183 ( .A(n540), .B(n53), .Z(\ab[26][47] ) );
  NR2 U3184 ( .A(n541), .B(n53), .Z(\ab[26][46] ) );
  NR2 U3185 ( .A(n542), .B(n53), .Z(\ab[26][45] ) );
  NR2 U3186 ( .A(n543), .B(n53), .Z(\ab[26][44] ) );
  NR2 U3187 ( .A(n544), .B(n53), .Z(\ab[26][43] ) );
  NR2 U3188 ( .A(n545), .B(n53), .Z(\ab[26][42] ) );
  NR2 U3189 ( .A(n546), .B(n53), .Z(\ab[26][41] ) );
  NR2 U3190 ( .A(n547), .B(n53), .Z(\ab[26][40] ) );
  NR2 U3191 ( .A(n548), .B(n53), .Z(\ab[26][39] ) );
  NR2 U3192 ( .A(n492), .B(n60), .Z(\ab[25][95] ) );
  NR2 U3193 ( .A(n493), .B(n60), .Z(\ab[25][94] ) );
  NR2 U3194 ( .A(n494), .B(n60), .Z(\ab[25][93] ) );
  NR2 U3195 ( .A(n495), .B(n60), .Z(\ab[25][92] ) );
  NR2 U3196 ( .A(n496), .B(n60), .Z(\ab[25][91] ) );
  NR2 U3197 ( .A(n497), .B(n60), .Z(\ab[25][90] ) );
  NR2 U3198 ( .A(n498), .B(n60), .Z(\ab[25][89] ) );
  NR2 U3199 ( .A(n499), .B(n60), .Z(\ab[25][88] ) );
  NR2 U3200 ( .A(n500), .B(n60), .Z(\ab[25][87] ) );
  NR2 U3201 ( .A(n501), .B(n60), .Z(\ab[25][86] ) );
  NR2 U3202 ( .A(n502), .B(n60), .Z(\ab[25][85] ) );
  NR2 U3203 ( .A(n503), .B(n60), .Z(\ab[25][84] ) );
  NR2 U3204 ( .A(n504), .B(n61), .Z(\ab[25][83] ) );
  NR2 U3205 ( .A(n505), .B(n61), .Z(\ab[25][82] ) );
  NR2 U3206 ( .A(n506), .B(n61), .Z(\ab[25][81] ) );
  NR2 U3207 ( .A(n507), .B(n61), .Z(\ab[25][80] ) );
  NR2 U3208 ( .A(n508), .B(n61), .Z(\ab[25][79] ) );
  NR2 U3209 ( .A(n509), .B(n61), .Z(\ab[25][78] ) );
  NR2 U3210 ( .A(n510), .B(n61), .Z(\ab[25][77] ) );
  NR2 U3211 ( .A(n511), .B(n61), .Z(\ab[25][76] ) );
  NR2 U3212 ( .A(n512), .B(n61), .Z(\ab[25][75] ) );
  NR2 U3213 ( .A(n513), .B(n61), .Z(\ab[25][74] ) );
  NR2 U3214 ( .A(n514), .B(n61), .Z(\ab[25][73] ) );
  NR2 U3215 ( .A(n515), .B(n61), .Z(\ab[25][72] ) );
  NR2 U3216 ( .A(n516), .B(n62), .Z(\ab[25][71] ) );
  NR2 U3217 ( .A(n517), .B(n62), .Z(\ab[25][70] ) );
  NR2 U3218 ( .A(n518), .B(n62), .Z(\ab[25][69] ) );
  NR2 U3219 ( .A(n519), .B(n62), .Z(\ab[25][68] ) );
  NR2 U3220 ( .A(n520), .B(n62), .Z(\ab[25][67] ) );
  NR2 U3221 ( .A(n521), .B(n62), .Z(\ab[25][66] ) );
  NR2 U3222 ( .A(n522), .B(n62), .Z(\ab[25][65] ) );
  NR2 U3223 ( .A(n523), .B(n62), .Z(\ab[25][64] ) );
  NR2 U3224 ( .A(n524), .B(n62), .Z(\ab[25][63] ) );
  NR2 U3225 ( .A(n525), .B(n62), .Z(\ab[25][62] ) );
  NR2 U3226 ( .A(n526), .B(n62), .Z(\ab[25][61] ) );
  NR2 U3227 ( .A(n527), .B(n62), .Z(\ab[25][60] ) );
  NR2 U3228 ( .A(n528), .B(n63), .Z(\ab[25][59] ) );
  NR2 U3229 ( .A(n529), .B(n63), .Z(\ab[25][58] ) );
  NR2 U3230 ( .A(n530), .B(n63), .Z(\ab[25][57] ) );
  NR2 U3231 ( .A(n531), .B(n63), .Z(\ab[25][56] ) );
  NR2 U3232 ( .A(n532), .B(n63), .Z(\ab[25][55] ) );
  NR2 U3233 ( .A(n533), .B(n63), .Z(\ab[25][54] ) );
  NR2 U3234 ( .A(n534), .B(n63), .Z(\ab[25][53] ) );
  NR2 U3235 ( .A(n535), .B(n63), .Z(\ab[25][52] ) );
  NR2 U3236 ( .A(n536), .B(n63), .Z(\ab[25][51] ) );
  NR2 U3237 ( .A(n537), .B(n63), .Z(\ab[25][50] ) );
  NR2 U3238 ( .A(n538), .B(n63), .Z(\ab[25][49] ) );
  NR2 U3239 ( .A(n539), .B(n63), .Z(\ab[25][48] ) );
  NR2 U3240 ( .A(n540), .B(n64), .Z(\ab[25][47] ) );
  NR2 U3241 ( .A(n541), .B(n64), .Z(\ab[25][46] ) );
  NR2 U3242 ( .A(n542), .B(n64), .Z(\ab[25][45] ) );
  NR2 U3243 ( .A(n543), .B(n64), .Z(\ab[25][44] ) );
  NR2 U3244 ( .A(n544), .B(n64), .Z(\ab[25][43] ) );
  NR2 U3245 ( .A(n545), .B(n64), .Z(\ab[25][42] ) );
  NR2 U3246 ( .A(n546), .B(n64), .Z(\ab[25][41] ) );
  NR2 U3247 ( .A(n547), .B(n64), .Z(\ab[25][40] ) );
  NR2 U3248 ( .A(n548), .B(n64), .Z(\ab[25][39] ) );
  NR2 U3249 ( .A(n492), .B(n71), .Z(\ab[24][95] ) );
  NR2 U3250 ( .A(n493), .B(n71), .Z(\ab[24][94] ) );
  NR2 U3251 ( .A(n494), .B(n71), .Z(\ab[24][93] ) );
  NR2 U3252 ( .A(n495), .B(n71), .Z(\ab[24][92] ) );
  NR2 U3253 ( .A(n496), .B(n71), .Z(\ab[24][91] ) );
  NR2 U3254 ( .A(n497), .B(n71), .Z(\ab[24][90] ) );
  NR2 U3255 ( .A(n498), .B(n71), .Z(\ab[24][89] ) );
  NR2 U3256 ( .A(n499), .B(n71), .Z(\ab[24][88] ) );
  NR2 U3257 ( .A(n500), .B(n71), .Z(\ab[24][87] ) );
  NR2 U3258 ( .A(n501), .B(n71), .Z(\ab[24][86] ) );
  NR2 U3259 ( .A(n502), .B(n71), .Z(\ab[24][85] ) );
  NR2 U3260 ( .A(n503), .B(n71), .Z(\ab[24][84] ) );
  NR2 U3261 ( .A(n504), .B(n72), .Z(\ab[24][83] ) );
  NR2 U3262 ( .A(n505), .B(n72), .Z(\ab[24][82] ) );
  NR2 U3263 ( .A(n506), .B(n72), .Z(\ab[24][81] ) );
  NR2 U3264 ( .A(n507), .B(n72), .Z(\ab[24][80] ) );
  NR2 U3265 ( .A(n508), .B(n72), .Z(\ab[24][79] ) );
  NR2 U3266 ( .A(n509), .B(n72), .Z(\ab[24][78] ) );
  NR2 U3267 ( .A(n510), .B(n72), .Z(\ab[24][77] ) );
  NR2 U3268 ( .A(n511), .B(n72), .Z(\ab[24][76] ) );
  NR2 U3269 ( .A(n512), .B(n72), .Z(\ab[24][75] ) );
  NR2 U3270 ( .A(n513), .B(n72), .Z(\ab[24][74] ) );
  NR2 U3271 ( .A(n514), .B(n72), .Z(\ab[24][73] ) );
  NR2 U3272 ( .A(n515), .B(n72), .Z(\ab[24][72] ) );
  NR2 U3273 ( .A(n516), .B(n73), .Z(\ab[24][71] ) );
  NR2 U3274 ( .A(n517), .B(n73), .Z(\ab[24][70] ) );
  NR2 U3275 ( .A(n518), .B(n73), .Z(\ab[24][69] ) );
  NR2 U3276 ( .A(n519), .B(n73), .Z(\ab[24][68] ) );
  NR2 U3277 ( .A(n520), .B(n73), .Z(\ab[24][67] ) );
  NR2 U3278 ( .A(n521), .B(n73), .Z(\ab[24][66] ) );
  NR2 U3279 ( .A(n522), .B(n73), .Z(\ab[24][65] ) );
  NR2 U3280 ( .A(n523), .B(n73), .Z(\ab[24][64] ) );
  NR2 U3281 ( .A(n524), .B(n73), .Z(\ab[24][63] ) );
  NR2 U3282 ( .A(n525), .B(n73), .Z(\ab[24][62] ) );
  NR2 U3283 ( .A(n526), .B(n73), .Z(\ab[24][61] ) );
  NR2 U3284 ( .A(n527), .B(n73), .Z(\ab[24][60] ) );
  NR2 U3285 ( .A(n528), .B(n74), .Z(\ab[24][59] ) );
  NR2 U3286 ( .A(n529), .B(n74), .Z(\ab[24][58] ) );
  NR2 U3287 ( .A(n530), .B(n74), .Z(\ab[24][57] ) );
  NR2 U3288 ( .A(n531), .B(n74), .Z(\ab[24][56] ) );
  NR2 U3289 ( .A(n532), .B(n74), .Z(\ab[24][55] ) );
  NR2 U3290 ( .A(n533), .B(n74), .Z(\ab[24][54] ) );
  NR2 U3291 ( .A(n534), .B(n74), .Z(\ab[24][53] ) );
  NR2 U3292 ( .A(n535), .B(n74), .Z(\ab[24][52] ) );
  NR2 U3293 ( .A(n536), .B(n74), .Z(\ab[24][51] ) );
  NR2 U3294 ( .A(n537), .B(n74), .Z(\ab[24][50] ) );
  NR2 U3295 ( .A(n538), .B(n74), .Z(\ab[24][49] ) );
  NR2 U3296 ( .A(n539), .B(n74), .Z(\ab[24][48] ) );
  NR2 U3297 ( .A(n540), .B(n75), .Z(\ab[24][47] ) );
  NR2 U3298 ( .A(n541), .B(n75), .Z(\ab[24][46] ) );
  NR2 U3299 ( .A(n542), .B(n75), .Z(\ab[24][45] ) );
  NR2 U3300 ( .A(n543), .B(n75), .Z(\ab[24][44] ) );
  NR2 U3301 ( .A(n544), .B(n75), .Z(\ab[24][43] ) );
  NR2 U3302 ( .A(n545), .B(n75), .Z(\ab[24][42] ) );
  NR2 U3303 ( .A(n546), .B(n75), .Z(\ab[24][41] ) );
  NR2 U3304 ( .A(n547), .B(n75), .Z(\ab[24][40] ) );
  NR2 U3305 ( .A(n548), .B(n75), .Z(\ab[24][39] ) );
  NR2 U3306 ( .A(n492), .B(n82), .Z(\ab[23][95] ) );
  NR2 U3307 ( .A(n493), .B(n82), .Z(\ab[23][94] ) );
  NR2 U3308 ( .A(n494), .B(n82), .Z(\ab[23][93] ) );
  NR2 U3309 ( .A(n495), .B(n82), .Z(\ab[23][92] ) );
  NR2 U3310 ( .A(n496), .B(n82), .Z(\ab[23][91] ) );
  NR2 U3311 ( .A(n497), .B(n82), .Z(\ab[23][90] ) );
  NR2 U3312 ( .A(n498), .B(n82), .Z(\ab[23][89] ) );
  NR2 U3313 ( .A(n499), .B(n82), .Z(\ab[23][88] ) );
  NR2 U3314 ( .A(n500), .B(n82), .Z(\ab[23][87] ) );
  NR2 U3315 ( .A(n501), .B(n82), .Z(\ab[23][86] ) );
  NR2 U3316 ( .A(n502), .B(n82), .Z(\ab[23][85] ) );
  NR2 U3317 ( .A(n503), .B(n82), .Z(\ab[23][84] ) );
  NR2 U3318 ( .A(n504), .B(n83), .Z(\ab[23][83] ) );
  NR2 U3319 ( .A(n505), .B(n83), .Z(\ab[23][82] ) );
  NR2 U3320 ( .A(n506), .B(n83), .Z(\ab[23][81] ) );
  NR2 U3321 ( .A(n507), .B(n83), .Z(\ab[23][80] ) );
  NR2 U3322 ( .A(n508), .B(n83), .Z(\ab[23][79] ) );
  NR2 U3323 ( .A(n509), .B(n83), .Z(\ab[23][78] ) );
  NR2 U3324 ( .A(n510), .B(n83), .Z(\ab[23][77] ) );
  NR2 U3325 ( .A(n511), .B(n83), .Z(\ab[23][76] ) );
  NR2 U3326 ( .A(n512), .B(n83), .Z(\ab[23][75] ) );
  NR2 U3327 ( .A(n513), .B(n83), .Z(\ab[23][74] ) );
  NR2 U3328 ( .A(n514), .B(n83), .Z(\ab[23][73] ) );
  NR2 U3329 ( .A(n515), .B(n83), .Z(\ab[23][72] ) );
  NR2 U3330 ( .A(n516), .B(n84), .Z(\ab[23][71] ) );
  NR2 U3331 ( .A(n517), .B(n84), .Z(\ab[23][70] ) );
  NR2 U3332 ( .A(n518), .B(n84), .Z(\ab[23][69] ) );
  NR2 U3333 ( .A(n519), .B(n84), .Z(\ab[23][68] ) );
  NR2 U3334 ( .A(n520), .B(n84), .Z(\ab[23][67] ) );
  NR2 U3335 ( .A(n521), .B(n84), .Z(\ab[23][66] ) );
  NR2 U3336 ( .A(n522), .B(n84), .Z(\ab[23][65] ) );
  NR2 U3337 ( .A(n523), .B(n84), .Z(\ab[23][64] ) );
  NR2 U3338 ( .A(n524), .B(n84), .Z(\ab[23][63] ) );
  NR2 U3339 ( .A(n525), .B(n84), .Z(\ab[23][62] ) );
  NR2 U3340 ( .A(n526), .B(n84), .Z(\ab[23][61] ) );
  NR2 U3341 ( .A(n527), .B(n84), .Z(\ab[23][60] ) );
  NR2 U3342 ( .A(n528), .B(n85), .Z(\ab[23][59] ) );
  NR2 U3343 ( .A(n529), .B(n85), .Z(\ab[23][58] ) );
  NR2 U3344 ( .A(n530), .B(n85), .Z(\ab[23][57] ) );
  NR2 U3345 ( .A(n531), .B(n85), .Z(\ab[23][56] ) );
  NR2 U3346 ( .A(n532), .B(n85), .Z(\ab[23][55] ) );
  NR2 U3347 ( .A(n533), .B(n85), .Z(\ab[23][54] ) );
  NR2 U3348 ( .A(n534), .B(n85), .Z(\ab[23][53] ) );
  NR2 U3349 ( .A(n535), .B(n85), .Z(\ab[23][52] ) );
  NR2 U3350 ( .A(n536), .B(n85), .Z(\ab[23][51] ) );
  NR2 U3351 ( .A(n537), .B(n85), .Z(\ab[23][50] ) );
  NR2 U3352 ( .A(n538), .B(n85), .Z(\ab[23][49] ) );
  NR2 U3353 ( .A(n539), .B(n85), .Z(\ab[23][48] ) );
  NR2 U3354 ( .A(n540), .B(n86), .Z(\ab[23][47] ) );
  NR2 U3355 ( .A(n541), .B(n86), .Z(\ab[23][46] ) );
  NR2 U3356 ( .A(n542), .B(n86), .Z(\ab[23][45] ) );
  NR2 U3357 ( .A(n543), .B(n86), .Z(\ab[23][44] ) );
  NR2 U3358 ( .A(n544), .B(n86), .Z(\ab[23][43] ) );
  NR2 U3359 ( .A(n545), .B(n86), .Z(\ab[23][42] ) );
  NR2 U3360 ( .A(n546), .B(n86), .Z(\ab[23][41] ) );
  NR2 U3361 ( .A(n547), .B(n86), .Z(\ab[23][40] ) );
  NR2 U3362 ( .A(n548), .B(n86), .Z(\ab[23][39] ) );
  NR2 U3363 ( .A(n492), .B(n4), .Z(\ab[22][95] ) );
  NR2 U3364 ( .A(n493), .B(n4), .Z(\ab[22][94] ) );
  NR2 U3365 ( .A(n494), .B(n4), .Z(\ab[22][93] ) );
  NR2 U3366 ( .A(n495), .B(n4), .Z(\ab[22][92] ) );
  NR2 U3367 ( .A(n496), .B(n4), .Z(\ab[22][91] ) );
  NR2 U3368 ( .A(n497), .B(n4), .Z(\ab[22][90] ) );
  NR2 U3369 ( .A(n498), .B(n4), .Z(\ab[22][89] ) );
  NR2 U3370 ( .A(n499), .B(n4), .Z(\ab[22][88] ) );
  NR2 U3371 ( .A(n500), .B(n4), .Z(\ab[22][87] ) );
  NR2 U3372 ( .A(n501), .B(n4), .Z(\ab[22][86] ) );
  NR2 U3373 ( .A(n502), .B(n4), .Z(\ab[22][85] ) );
  NR2 U3374 ( .A(n503), .B(n4), .Z(\ab[22][84] ) );
  NR2 U3375 ( .A(n504), .B(n557), .Z(\ab[22][83] ) );
  NR2 U3376 ( .A(n505), .B(n4), .Z(\ab[22][82] ) );
  NR2 U3377 ( .A(n506), .B(n557), .Z(\ab[22][81] ) );
  NR2 U3378 ( .A(n507), .B(n4), .Z(\ab[22][80] ) );
  NR2 U3379 ( .A(n508), .B(n4), .Z(\ab[22][79] ) );
  NR2 U3380 ( .A(n509), .B(n4), .Z(\ab[22][78] ) );
  NR2 U3381 ( .A(n510), .B(n4), .Z(\ab[22][77] ) );
  NR2 U3382 ( .A(n511), .B(n4), .Z(\ab[22][76] ) );
  NR2 U3383 ( .A(n512), .B(n4), .Z(\ab[22][75] ) );
  NR2 U3384 ( .A(n513), .B(n4), .Z(\ab[22][74] ) );
  NR2 U3385 ( .A(n514), .B(n4), .Z(\ab[22][73] ) );
  NR2 U3386 ( .A(n515), .B(n4), .Z(\ab[22][72] ) );
  NR2 U3387 ( .A(n516), .B(n557), .Z(\ab[22][71] ) );
  NR2 U3388 ( .A(n517), .B(n557), .Z(\ab[22][70] ) );
  NR2 U3389 ( .A(n518), .B(n557), .Z(\ab[22][69] ) );
  NR2 U3390 ( .A(n519), .B(n4), .Z(\ab[22][68] ) );
  NR2 U3391 ( .A(n520), .B(n557), .Z(\ab[22][67] ) );
  NR2 U3392 ( .A(n521), .B(n557), .Z(\ab[22][66] ) );
  NR2 U3393 ( .A(n522), .B(n557), .Z(\ab[22][65] ) );
  NR2 U3394 ( .A(n523), .B(n4), .Z(\ab[22][64] ) );
  NR2 U3395 ( .A(n524), .B(n557), .Z(\ab[22][63] ) );
  NR2 U3396 ( .A(n525), .B(n557), .Z(\ab[22][62] ) );
  NR2 U3397 ( .A(n526), .B(n557), .Z(\ab[22][61] ) );
  NR2 U3398 ( .A(n527), .B(n4), .Z(\ab[22][60] ) );
  NR2 U3399 ( .A(n528), .B(n557), .Z(\ab[22][59] ) );
  NR2 U3400 ( .A(n529), .B(n557), .Z(\ab[22][58] ) );
  NR2 U3401 ( .A(n530), .B(n557), .Z(\ab[22][57] ) );
  NR2 U3402 ( .A(n531), .B(n557), .Z(\ab[22][56] ) );
  NR2 U3403 ( .A(n532), .B(n557), .Z(\ab[22][55] ) );
  NR2 U3404 ( .A(n533), .B(n557), .Z(\ab[22][54] ) );
  NR2 U3405 ( .A(n534), .B(n557), .Z(\ab[22][53] ) );
  NR2 U3406 ( .A(n535), .B(n557), .Z(\ab[22][52] ) );
  NR2 U3407 ( .A(n536), .B(n557), .Z(\ab[22][51] ) );
  NR2 U3408 ( .A(n537), .B(n557), .Z(\ab[22][50] ) );
  NR2 U3409 ( .A(n538), .B(n557), .Z(\ab[22][49] ) );
  NR2 U3410 ( .A(n539), .B(n557), .Z(\ab[22][48] ) );
  NR2 U3411 ( .A(n540), .B(n557), .Z(\ab[22][47] ) );
  NR2 U3412 ( .A(n541), .B(n557), .Z(\ab[22][46] ) );
  NR2 U3413 ( .A(n542), .B(n557), .Z(\ab[22][45] ) );
  NR2 U3414 ( .A(n543), .B(n557), .Z(\ab[22][44] ) );
  NR2 U3415 ( .A(n544), .B(n557), .Z(\ab[22][43] ) );
  NR2 U3416 ( .A(n545), .B(n557), .Z(\ab[22][42] ) );
  NR2 U3417 ( .A(n546), .B(n557), .Z(\ab[22][41] ) );
  NR2 U3418 ( .A(n547), .B(n557), .Z(\ab[22][40] ) );
  NR2 U3419 ( .A(n548), .B(n557), .Z(\ab[22][39] ) );
  NR2 U3420 ( .A(n492), .B(n98), .Z(\ab[21][95] ) );
  NR2 U3421 ( .A(n493), .B(n98), .Z(\ab[21][94] ) );
  NR2 U3422 ( .A(n494), .B(n98), .Z(\ab[21][93] ) );
  NR2 U3423 ( .A(n495), .B(n98), .Z(\ab[21][92] ) );
  NR2 U3424 ( .A(n496), .B(n98), .Z(\ab[21][91] ) );
  NR2 U3425 ( .A(n497), .B(n98), .Z(\ab[21][90] ) );
  NR2 U3426 ( .A(n498), .B(n98), .Z(\ab[21][89] ) );
  NR2 U3427 ( .A(n499), .B(n98), .Z(\ab[21][88] ) );
  NR2 U3428 ( .A(n500), .B(n98), .Z(\ab[21][87] ) );
  NR2 U3429 ( .A(n501), .B(n98), .Z(\ab[21][86] ) );
  NR2 U3430 ( .A(n502), .B(n98), .Z(\ab[21][85] ) );
  NR2 U3431 ( .A(n503), .B(n98), .Z(\ab[21][84] ) );
  NR2 U3432 ( .A(n504), .B(n99), .Z(\ab[21][83] ) );
  NR2 U3433 ( .A(n505), .B(n99), .Z(\ab[21][82] ) );
  NR2 U3434 ( .A(n506), .B(n99), .Z(\ab[21][81] ) );
  NR2 U3435 ( .A(n507), .B(n99), .Z(\ab[21][80] ) );
  NR2 U3436 ( .A(n508), .B(n99), .Z(\ab[21][79] ) );
  NR2 U3437 ( .A(n509), .B(n99), .Z(\ab[21][78] ) );
  NR2 U3438 ( .A(n510), .B(n99), .Z(\ab[21][77] ) );
  NR2 U3439 ( .A(n511), .B(n99), .Z(\ab[21][76] ) );
  NR2 U3440 ( .A(n512), .B(n99), .Z(\ab[21][75] ) );
  NR2 U3441 ( .A(n513), .B(n99), .Z(\ab[21][74] ) );
  NR2 U3442 ( .A(n514), .B(n99), .Z(\ab[21][73] ) );
  NR2 U3443 ( .A(n515), .B(n99), .Z(\ab[21][72] ) );
  NR2 U3444 ( .A(n516), .B(n100), .Z(\ab[21][71] ) );
  NR2 U3445 ( .A(n517), .B(n100), .Z(\ab[21][70] ) );
  NR2 U3446 ( .A(n518), .B(n100), .Z(\ab[21][69] ) );
  NR2 U3447 ( .A(n519), .B(n100), .Z(\ab[21][68] ) );
  NR2 U3448 ( .A(n520), .B(n100), .Z(\ab[21][67] ) );
  NR2 U3449 ( .A(n521), .B(n100), .Z(\ab[21][66] ) );
  NR2 U3450 ( .A(n522), .B(n100), .Z(\ab[21][65] ) );
  NR2 U3451 ( .A(n523), .B(n100), .Z(\ab[21][64] ) );
  NR2 U3452 ( .A(n524), .B(n100), .Z(\ab[21][63] ) );
  NR2 U3453 ( .A(n525), .B(n100), .Z(\ab[21][62] ) );
  NR2 U3454 ( .A(n526), .B(n100), .Z(\ab[21][61] ) );
  NR2 U3455 ( .A(n527), .B(n100), .Z(\ab[21][60] ) );
  NR2 U3456 ( .A(n528), .B(n101), .Z(\ab[21][59] ) );
  NR2 U3457 ( .A(n529), .B(n101), .Z(\ab[21][58] ) );
  NR2 U3458 ( .A(n530), .B(n101), .Z(\ab[21][57] ) );
  NR2 U3459 ( .A(n531), .B(n101), .Z(\ab[21][56] ) );
  NR2 U3460 ( .A(n532), .B(n101), .Z(\ab[21][55] ) );
  NR2 U3461 ( .A(n533), .B(n101), .Z(\ab[21][54] ) );
  NR2 U3462 ( .A(n534), .B(n101), .Z(\ab[21][53] ) );
  NR2 U3463 ( .A(n535), .B(n101), .Z(\ab[21][52] ) );
  NR2 U3464 ( .A(n536), .B(n101), .Z(\ab[21][51] ) );
  NR2 U3465 ( .A(n537), .B(n101), .Z(\ab[21][50] ) );
  NR2 U3466 ( .A(n538), .B(n101), .Z(\ab[21][49] ) );
  NR2 U3467 ( .A(n539), .B(n101), .Z(\ab[21][48] ) );
  NR2 U3468 ( .A(n540), .B(n102), .Z(\ab[21][47] ) );
  NR2 U3469 ( .A(n541), .B(n102), .Z(\ab[21][46] ) );
  NR2 U3470 ( .A(n542), .B(n102), .Z(\ab[21][45] ) );
  NR2 U3471 ( .A(n543), .B(n102), .Z(\ab[21][44] ) );
  NR2 U3472 ( .A(n544), .B(n102), .Z(\ab[21][43] ) );
  NR2 U3473 ( .A(n545), .B(n102), .Z(\ab[21][42] ) );
  NR2 U3474 ( .A(n546), .B(n102), .Z(\ab[21][41] ) );
  NR2 U3475 ( .A(n547), .B(n102), .Z(\ab[21][40] ) );
  NR2 U3476 ( .A(n548), .B(n102), .Z(\ab[21][39] ) );
  NR2 U3477 ( .A(n492), .B(n109), .Z(\ab[20][95] ) );
  NR2 U3478 ( .A(n493), .B(n109), .Z(\ab[20][94] ) );
  NR2 U3479 ( .A(n494), .B(n109), .Z(\ab[20][93] ) );
  NR2 U3480 ( .A(n495), .B(n109), .Z(\ab[20][92] ) );
  NR2 U3481 ( .A(n496), .B(n109), .Z(\ab[20][91] ) );
  NR2 U3482 ( .A(n497), .B(n109), .Z(\ab[20][90] ) );
  NR2 U3483 ( .A(n498), .B(n109), .Z(\ab[20][89] ) );
  NR2 U3484 ( .A(n499), .B(n109), .Z(\ab[20][88] ) );
  NR2 U3485 ( .A(n500), .B(n109), .Z(\ab[20][87] ) );
  NR2 U3486 ( .A(n501), .B(n109), .Z(\ab[20][86] ) );
  NR2 U3487 ( .A(n502), .B(n109), .Z(\ab[20][85] ) );
  NR2 U3488 ( .A(n503), .B(n109), .Z(\ab[20][84] ) );
  NR2 U3489 ( .A(n504), .B(n110), .Z(\ab[20][83] ) );
  NR2 U3490 ( .A(n505), .B(n110), .Z(\ab[20][82] ) );
  NR2 U3491 ( .A(n506), .B(n110), .Z(\ab[20][81] ) );
  NR2 U3492 ( .A(n507), .B(n110), .Z(\ab[20][80] ) );
  NR2 U3493 ( .A(n508), .B(n110), .Z(\ab[20][79] ) );
  NR2 U3494 ( .A(n509), .B(n110), .Z(\ab[20][78] ) );
  NR2 U3495 ( .A(n510), .B(n110), .Z(\ab[20][77] ) );
  NR2 U3496 ( .A(n511), .B(n110), .Z(\ab[20][76] ) );
  NR2 U3497 ( .A(n512), .B(n110), .Z(\ab[20][75] ) );
  NR2 U3498 ( .A(n513), .B(n110), .Z(\ab[20][74] ) );
  NR2 U3499 ( .A(n514), .B(n110), .Z(\ab[20][73] ) );
  NR2 U3500 ( .A(n515), .B(n110), .Z(\ab[20][72] ) );
  NR2 U3501 ( .A(n516), .B(n111), .Z(\ab[20][71] ) );
  NR2 U3502 ( .A(n517), .B(n111), .Z(\ab[20][70] ) );
  NR2 U3503 ( .A(n518), .B(n111), .Z(\ab[20][69] ) );
  NR2 U3504 ( .A(n519), .B(n111), .Z(\ab[20][68] ) );
  NR2 U3505 ( .A(n520), .B(n111), .Z(\ab[20][67] ) );
  NR2 U3506 ( .A(n521), .B(n111), .Z(\ab[20][66] ) );
  NR2 U3507 ( .A(n522), .B(n111), .Z(\ab[20][65] ) );
  NR2 U3508 ( .A(n523), .B(n111), .Z(\ab[20][64] ) );
  NR2 U3509 ( .A(n524), .B(n111), .Z(\ab[20][63] ) );
  NR2 U3510 ( .A(n525), .B(n111), .Z(\ab[20][62] ) );
  NR2 U3511 ( .A(n526), .B(n111), .Z(\ab[20][61] ) );
  NR2 U3512 ( .A(n527), .B(n111), .Z(\ab[20][60] ) );
  NR2 U3513 ( .A(n528), .B(n112), .Z(\ab[20][59] ) );
  NR2 U3514 ( .A(n529), .B(n112), .Z(\ab[20][58] ) );
  NR2 U3515 ( .A(n530), .B(n112), .Z(\ab[20][57] ) );
  NR2 U3516 ( .A(n531), .B(n112), .Z(\ab[20][56] ) );
  NR2 U3517 ( .A(n532), .B(n112), .Z(\ab[20][55] ) );
  NR2 U3518 ( .A(n533), .B(n112), .Z(\ab[20][54] ) );
  NR2 U3519 ( .A(n534), .B(n112), .Z(\ab[20][53] ) );
  NR2 U3520 ( .A(n535), .B(n112), .Z(\ab[20][52] ) );
  NR2 U3521 ( .A(n536), .B(n112), .Z(\ab[20][51] ) );
  NR2 U3522 ( .A(n537), .B(n112), .Z(\ab[20][50] ) );
  NR2 U3523 ( .A(n538), .B(n112), .Z(\ab[20][49] ) );
  NR2 U3524 ( .A(n539), .B(n112), .Z(\ab[20][48] ) );
  NR2 U3525 ( .A(n540), .B(n113), .Z(\ab[20][47] ) );
  NR2 U3526 ( .A(n541), .B(n113), .Z(\ab[20][46] ) );
  NR2 U3527 ( .A(n542), .B(n113), .Z(\ab[20][45] ) );
  NR2 U3528 ( .A(n543), .B(n113), .Z(\ab[20][44] ) );
  NR2 U3529 ( .A(n544), .B(n113), .Z(\ab[20][43] ) );
  NR2 U3530 ( .A(n545), .B(n113), .Z(\ab[20][42] ) );
  NR2 U3531 ( .A(n546), .B(n113), .Z(\ab[20][41] ) );
  NR2 U3532 ( .A(n547), .B(n113), .Z(\ab[20][40] ) );
  NR2 U3533 ( .A(n548), .B(n113), .Z(\ab[20][39] ) );
  NR2 U3534 ( .A(n492), .B(n120), .Z(\ab[19][95] ) );
  NR2 U3535 ( .A(n493), .B(n120), .Z(\ab[19][94] ) );
  NR2 U3536 ( .A(n494), .B(n120), .Z(\ab[19][93] ) );
  NR2 U3537 ( .A(n495), .B(n120), .Z(\ab[19][92] ) );
  NR2 U3538 ( .A(n496), .B(n120), .Z(\ab[19][91] ) );
  NR2 U3539 ( .A(n497), .B(n120), .Z(\ab[19][90] ) );
  NR2 U3540 ( .A(n498), .B(n120), .Z(\ab[19][89] ) );
  NR2 U3541 ( .A(n499), .B(n120), .Z(\ab[19][88] ) );
  NR2 U3542 ( .A(n500), .B(n120), .Z(\ab[19][87] ) );
  NR2 U3543 ( .A(n501), .B(n120), .Z(\ab[19][86] ) );
  NR2 U3544 ( .A(n502), .B(n120), .Z(\ab[19][85] ) );
  NR2 U3545 ( .A(n503), .B(n120), .Z(\ab[19][84] ) );
  NR2 U3546 ( .A(n504), .B(n121), .Z(\ab[19][83] ) );
  NR2 U3547 ( .A(n505), .B(n121), .Z(\ab[19][82] ) );
  NR2 U3548 ( .A(n506), .B(n121), .Z(\ab[19][81] ) );
  NR2 U3549 ( .A(n507), .B(n121), .Z(\ab[19][80] ) );
  NR2 U3550 ( .A(n508), .B(n121), .Z(\ab[19][79] ) );
  NR2 U3551 ( .A(n509), .B(n121), .Z(\ab[19][78] ) );
  NR2 U3552 ( .A(n510), .B(n121), .Z(\ab[19][77] ) );
  NR2 U3553 ( .A(n511), .B(n121), .Z(\ab[19][76] ) );
  NR2 U3554 ( .A(n512), .B(n121), .Z(\ab[19][75] ) );
  NR2 U3555 ( .A(n513), .B(n121), .Z(\ab[19][74] ) );
  NR2 U3556 ( .A(n514), .B(n121), .Z(\ab[19][73] ) );
  NR2 U3557 ( .A(n515), .B(n121), .Z(\ab[19][72] ) );
  NR2 U3558 ( .A(n516), .B(n122), .Z(\ab[19][71] ) );
  NR2 U3559 ( .A(n517), .B(n122), .Z(\ab[19][70] ) );
  NR2 U3560 ( .A(n518), .B(n122), .Z(\ab[19][69] ) );
  NR2 U3561 ( .A(n519), .B(n122), .Z(\ab[19][68] ) );
  NR2 U3562 ( .A(n520), .B(n122), .Z(\ab[19][67] ) );
  NR2 U3563 ( .A(n521), .B(n122), .Z(\ab[19][66] ) );
  NR2 U3564 ( .A(n522), .B(n122), .Z(\ab[19][65] ) );
  NR2 U3565 ( .A(n523), .B(n122), .Z(\ab[19][64] ) );
  NR2 U3566 ( .A(n524), .B(n122), .Z(\ab[19][63] ) );
  NR2 U3567 ( .A(n525), .B(n122), .Z(\ab[19][62] ) );
  NR2 U3568 ( .A(n526), .B(n122), .Z(\ab[19][61] ) );
  NR2 U3569 ( .A(n527), .B(n122), .Z(\ab[19][60] ) );
  NR2 U3570 ( .A(n528), .B(n123), .Z(\ab[19][59] ) );
  NR2 U3571 ( .A(n529), .B(n123), .Z(\ab[19][58] ) );
  NR2 U3572 ( .A(n530), .B(n123), .Z(\ab[19][57] ) );
  NR2 U3573 ( .A(n531), .B(n123), .Z(\ab[19][56] ) );
  NR2 U3574 ( .A(n532), .B(n123), .Z(\ab[19][55] ) );
  NR2 U3575 ( .A(n533), .B(n123), .Z(\ab[19][54] ) );
  NR2 U3576 ( .A(n534), .B(n123), .Z(\ab[19][53] ) );
  NR2 U3577 ( .A(n535), .B(n123), .Z(\ab[19][52] ) );
  NR2 U3578 ( .A(n536), .B(n123), .Z(\ab[19][51] ) );
  NR2 U3579 ( .A(n537), .B(n123), .Z(\ab[19][50] ) );
  NR2 U3580 ( .A(n538), .B(n123), .Z(\ab[19][49] ) );
  NR2 U3581 ( .A(n539), .B(n123), .Z(\ab[19][48] ) );
  NR2 U3582 ( .A(n540), .B(n124), .Z(\ab[19][47] ) );
  NR2 U3583 ( .A(n541), .B(n124), .Z(\ab[19][46] ) );
  NR2 U3584 ( .A(n542), .B(n124), .Z(\ab[19][45] ) );
  NR2 U3585 ( .A(n543), .B(n124), .Z(\ab[19][44] ) );
  NR2 U3586 ( .A(n544), .B(n124), .Z(\ab[19][43] ) );
  NR2 U3587 ( .A(n545), .B(n124), .Z(\ab[19][42] ) );
  NR2 U3588 ( .A(n546), .B(n124), .Z(\ab[19][41] ) );
  NR2 U3589 ( .A(n547), .B(n124), .Z(\ab[19][40] ) );
  NR2 U3590 ( .A(n548), .B(n124), .Z(\ab[19][39] ) );
  NR2 U3591 ( .A(n492), .B(n131), .Z(\ab[18][95] ) );
  NR2 U3592 ( .A(n493), .B(n131), .Z(\ab[18][94] ) );
  NR2 U3593 ( .A(n494), .B(n131), .Z(\ab[18][93] ) );
  NR2 U3594 ( .A(n495), .B(n131), .Z(\ab[18][92] ) );
  NR2 U3595 ( .A(n496), .B(n131), .Z(\ab[18][91] ) );
  NR2 U3596 ( .A(n497), .B(n131), .Z(\ab[18][90] ) );
  NR2 U3597 ( .A(n498), .B(n131), .Z(\ab[18][89] ) );
  NR2 U3598 ( .A(n499), .B(n131), .Z(\ab[18][88] ) );
  NR2 U3599 ( .A(n500), .B(n131), .Z(\ab[18][87] ) );
  NR2 U3600 ( .A(n501), .B(n131), .Z(\ab[18][86] ) );
  NR2 U3601 ( .A(n502), .B(n131), .Z(\ab[18][85] ) );
  NR2 U3602 ( .A(n503), .B(n131), .Z(\ab[18][84] ) );
  NR2 U3603 ( .A(n504), .B(n132), .Z(\ab[18][83] ) );
  NR2 U3604 ( .A(n505), .B(n132), .Z(\ab[18][82] ) );
  NR2 U3605 ( .A(n506), .B(n132), .Z(\ab[18][81] ) );
  NR2 U3606 ( .A(n507), .B(n132), .Z(\ab[18][80] ) );
  NR2 U3607 ( .A(n508), .B(n132), .Z(\ab[18][79] ) );
  NR2 U3608 ( .A(n509), .B(n132), .Z(\ab[18][78] ) );
  NR2 U3609 ( .A(n510), .B(n132), .Z(\ab[18][77] ) );
  NR2 U3610 ( .A(n511), .B(n132), .Z(\ab[18][76] ) );
  NR2 U3611 ( .A(n512), .B(n132), .Z(\ab[18][75] ) );
  NR2 U3612 ( .A(n513), .B(n132), .Z(\ab[18][74] ) );
  NR2 U3613 ( .A(n514), .B(n132), .Z(\ab[18][73] ) );
  NR2 U3614 ( .A(n515), .B(n132), .Z(\ab[18][72] ) );
  NR2 U3615 ( .A(n516), .B(n133), .Z(\ab[18][71] ) );
  NR2 U3616 ( .A(n517), .B(n133), .Z(\ab[18][70] ) );
  NR2 U3617 ( .A(n518), .B(n133), .Z(\ab[18][69] ) );
  NR2 U3618 ( .A(n519), .B(n133), .Z(\ab[18][68] ) );
  NR2 U3619 ( .A(n520), .B(n133), .Z(\ab[18][67] ) );
  NR2 U3620 ( .A(n521), .B(n133), .Z(\ab[18][66] ) );
  NR2 U3621 ( .A(n522), .B(n133), .Z(\ab[18][65] ) );
  NR2 U3622 ( .A(n523), .B(n133), .Z(\ab[18][64] ) );
  NR2 U3623 ( .A(n524), .B(n133), .Z(\ab[18][63] ) );
  NR2 U3624 ( .A(n525), .B(n133), .Z(\ab[18][62] ) );
  NR2 U3625 ( .A(n526), .B(n133), .Z(\ab[18][61] ) );
  NR2 U3626 ( .A(n527), .B(n133), .Z(\ab[18][60] ) );
  NR2 U3627 ( .A(n528), .B(n134), .Z(\ab[18][59] ) );
  NR2 U3628 ( .A(n529), .B(n134), .Z(\ab[18][58] ) );
  NR2 U3629 ( .A(n530), .B(n134), .Z(\ab[18][57] ) );
  NR2 U3630 ( .A(n531), .B(n134), .Z(\ab[18][56] ) );
  NR2 U3631 ( .A(n532), .B(n134), .Z(\ab[18][55] ) );
  NR2 U3632 ( .A(n533), .B(n134), .Z(\ab[18][54] ) );
  NR2 U3633 ( .A(n534), .B(n134), .Z(\ab[18][53] ) );
  NR2 U3634 ( .A(n535), .B(n134), .Z(\ab[18][52] ) );
  NR2 U3635 ( .A(n536), .B(n134), .Z(\ab[18][51] ) );
  NR2 U3636 ( .A(n537), .B(n134), .Z(\ab[18][50] ) );
  NR2 U3637 ( .A(n538), .B(n134), .Z(\ab[18][49] ) );
  NR2 U3638 ( .A(n539), .B(n134), .Z(\ab[18][48] ) );
  NR2 U3639 ( .A(n540), .B(n135), .Z(\ab[18][47] ) );
  NR2 U3640 ( .A(n541), .B(n135), .Z(\ab[18][46] ) );
  NR2 U3641 ( .A(n542), .B(n135), .Z(\ab[18][45] ) );
  NR2 U3642 ( .A(n543), .B(n135), .Z(\ab[18][44] ) );
  NR2 U3643 ( .A(n544), .B(n135), .Z(\ab[18][43] ) );
  NR2 U3644 ( .A(n545), .B(n135), .Z(\ab[18][42] ) );
  NR2 U3645 ( .A(n546), .B(n135), .Z(\ab[18][41] ) );
  NR2 U3646 ( .A(n547), .B(n135), .Z(\ab[18][40] ) );
  NR2 U3647 ( .A(n548), .B(n135), .Z(\ab[18][39] ) );
  NR2 U3648 ( .A(n492), .B(n142), .Z(\ab[17][95] ) );
  NR2 U3649 ( .A(n493), .B(n142), .Z(\ab[17][94] ) );
  NR2 U3650 ( .A(n494), .B(n142), .Z(\ab[17][93] ) );
  NR2 U3651 ( .A(n495), .B(n142), .Z(\ab[17][92] ) );
  NR2 U3652 ( .A(n496), .B(n142), .Z(\ab[17][91] ) );
  NR2 U3653 ( .A(n497), .B(n142), .Z(\ab[17][90] ) );
  NR2 U3654 ( .A(n498), .B(n142), .Z(\ab[17][89] ) );
  NR2 U3655 ( .A(n499), .B(n142), .Z(\ab[17][88] ) );
  NR2 U3656 ( .A(n500), .B(n142), .Z(\ab[17][87] ) );
  NR2 U3657 ( .A(n501), .B(n142), .Z(\ab[17][86] ) );
  NR2 U3658 ( .A(n502), .B(n142), .Z(\ab[17][85] ) );
  NR2 U3659 ( .A(n503), .B(n142), .Z(\ab[17][84] ) );
  NR2 U3660 ( .A(n504), .B(n143), .Z(\ab[17][83] ) );
  NR2 U3661 ( .A(n505), .B(n143), .Z(\ab[17][82] ) );
  NR2 U3662 ( .A(n506), .B(n143), .Z(\ab[17][81] ) );
  NR2 U3663 ( .A(n507), .B(n143), .Z(\ab[17][80] ) );
  NR2 U3664 ( .A(n508), .B(n143), .Z(\ab[17][79] ) );
  NR2 U3665 ( .A(n509), .B(n143), .Z(\ab[17][78] ) );
  NR2 U3666 ( .A(n510), .B(n143), .Z(\ab[17][77] ) );
  NR2 U3667 ( .A(n511), .B(n143), .Z(\ab[17][76] ) );
  NR2 U3668 ( .A(n512), .B(n143), .Z(\ab[17][75] ) );
  NR2 U3669 ( .A(n513), .B(n143), .Z(\ab[17][74] ) );
  NR2 U3670 ( .A(n514), .B(n143), .Z(\ab[17][73] ) );
  NR2 U3671 ( .A(n515), .B(n143), .Z(\ab[17][72] ) );
  NR2 U3672 ( .A(n516), .B(n144), .Z(\ab[17][71] ) );
  NR2 U3673 ( .A(n517), .B(n144), .Z(\ab[17][70] ) );
  NR2 U3674 ( .A(n518), .B(n144), .Z(\ab[17][69] ) );
  NR2 U3675 ( .A(n519), .B(n144), .Z(\ab[17][68] ) );
  NR2 U3676 ( .A(n520), .B(n144), .Z(\ab[17][67] ) );
  NR2 U3677 ( .A(n521), .B(n144), .Z(\ab[17][66] ) );
  NR2 U3678 ( .A(n522), .B(n144), .Z(\ab[17][65] ) );
  NR2 U3679 ( .A(n523), .B(n144), .Z(\ab[17][64] ) );
  NR2 U3680 ( .A(n524), .B(n144), .Z(\ab[17][63] ) );
  NR2 U3681 ( .A(n525), .B(n144), .Z(\ab[17][62] ) );
  NR2 U3682 ( .A(n526), .B(n144), .Z(\ab[17][61] ) );
  NR2 U3683 ( .A(n527), .B(n144), .Z(\ab[17][60] ) );
  NR2 U3684 ( .A(n528), .B(n145), .Z(\ab[17][59] ) );
  NR2 U3685 ( .A(n529), .B(n145), .Z(\ab[17][58] ) );
  NR2 U3686 ( .A(n530), .B(n145), .Z(\ab[17][57] ) );
  NR2 U3687 ( .A(n531), .B(n145), .Z(\ab[17][56] ) );
  NR2 U3688 ( .A(n532), .B(n145), .Z(\ab[17][55] ) );
  NR2 U3689 ( .A(n533), .B(n145), .Z(\ab[17][54] ) );
  NR2 U3690 ( .A(n534), .B(n145), .Z(\ab[17][53] ) );
  NR2 U3691 ( .A(n535), .B(n145), .Z(\ab[17][52] ) );
  NR2 U3692 ( .A(n536), .B(n145), .Z(\ab[17][51] ) );
  NR2 U3693 ( .A(n537), .B(n145), .Z(\ab[17][50] ) );
  NR2 U3694 ( .A(n538), .B(n145), .Z(\ab[17][49] ) );
  NR2 U3695 ( .A(n539), .B(n145), .Z(\ab[17][48] ) );
  NR2 U3696 ( .A(n540), .B(n146), .Z(\ab[17][47] ) );
  NR2 U3697 ( .A(n541), .B(n146), .Z(\ab[17][46] ) );
  NR2 U3698 ( .A(n542), .B(n146), .Z(\ab[17][45] ) );
  NR2 U3699 ( .A(n543), .B(n146), .Z(\ab[17][44] ) );
  NR2 U3700 ( .A(n544), .B(n146), .Z(\ab[17][43] ) );
  NR2 U3701 ( .A(n545), .B(n146), .Z(\ab[17][42] ) );
  NR2 U3702 ( .A(n546), .B(n146), .Z(\ab[17][41] ) );
  NR2 U3703 ( .A(n547), .B(n146), .Z(\ab[17][40] ) );
  NR2 U3704 ( .A(n548), .B(n146), .Z(\ab[17][39] ) );
  NR2 U3705 ( .A(n492), .B(n153), .Z(\ab[16][95] ) );
  NR2 U3706 ( .A(n493), .B(n153), .Z(\ab[16][94] ) );
  NR2 U3707 ( .A(n494), .B(n153), .Z(\ab[16][93] ) );
  NR2 U3708 ( .A(n495), .B(n153), .Z(\ab[16][92] ) );
  NR2 U3709 ( .A(n496), .B(n153), .Z(\ab[16][91] ) );
  NR2 U3710 ( .A(n497), .B(n153), .Z(\ab[16][90] ) );
  NR2 U3711 ( .A(n498), .B(n153), .Z(\ab[16][89] ) );
  NR2 U3712 ( .A(n499), .B(n153), .Z(\ab[16][88] ) );
  NR2 U3713 ( .A(n500), .B(n153), .Z(\ab[16][87] ) );
  NR2 U3714 ( .A(n501), .B(n153), .Z(\ab[16][86] ) );
  NR2 U3715 ( .A(n502), .B(n153), .Z(\ab[16][85] ) );
  NR2 U3716 ( .A(n503), .B(n153), .Z(\ab[16][84] ) );
  NR2 U3717 ( .A(n504), .B(n154), .Z(\ab[16][83] ) );
  NR2 U3718 ( .A(n505), .B(n154), .Z(\ab[16][82] ) );
  NR2 U3719 ( .A(n506), .B(n154), .Z(\ab[16][81] ) );
  NR2 U3720 ( .A(n507), .B(n154), .Z(\ab[16][80] ) );
  NR2 U3721 ( .A(n508), .B(n154), .Z(\ab[16][79] ) );
  NR2 U3722 ( .A(n509), .B(n154), .Z(\ab[16][78] ) );
  NR2 U3723 ( .A(n510), .B(n154), .Z(\ab[16][77] ) );
  NR2 U3724 ( .A(n511), .B(n154), .Z(\ab[16][76] ) );
  NR2 U3725 ( .A(n512), .B(n154), .Z(\ab[16][75] ) );
  NR2 U3726 ( .A(n513), .B(n154), .Z(\ab[16][74] ) );
  NR2 U3727 ( .A(n514), .B(n154), .Z(\ab[16][73] ) );
  NR2 U3728 ( .A(n515), .B(n154), .Z(\ab[16][72] ) );
  NR2 U3729 ( .A(n516), .B(n155), .Z(\ab[16][71] ) );
  NR2 U3730 ( .A(n517), .B(n155), .Z(\ab[16][70] ) );
  NR2 U3731 ( .A(n518), .B(n155), .Z(\ab[16][69] ) );
  NR2 U3732 ( .A(n519), .B(n155), .Z(\ab[16][68] ) );
  NR2 U3733 ( .A(n520), .B(n155), .Z(\ab[16][67] ) );
  NR2 U3734 ( .A(n521), .B(n155), .Z(\ab[16][66] ) );
  NR2 U3735 ( .A(n522), .B(n155), .Z(\ab[16][65] ) );
  NR2 U3736 ( .A(n523), .B(n155), .Z(\ab[16][64] ) );
  NR2 U3737 ( .A(n524), .B(n155), .Z(\ab[16][63] ) );
  NR2 U3738 ( .A(n525), .B(n155), .Z(\ab[16][62] ) );
  NR2 U3739 ( .A(n526), .B(n155), .Z(\ab[16][61] ) );
  NR2 U3740 ( .A(n527), .B(n155), .Z(\ab[16][60] ) );
  NR2 U3741 ( .A(n528), .B(n156), .Z(\ab[16][59] ) );
  NR2 U3742 ( .A(n529), .B(n156), .Z(\ab[16][58] ) );
  NR2 U3743 ( .A(n530), .B(n156), .Z(\ab[16][57] ) );
  NR2 U3744 ( .A(n531), .B(n156), .Z(\ab[16][56] ) );
  NR2 U3745 ( .A(n532), .B(n156), .Z(\ab[16][55] ) );
  NR2 U3746 ( .A(n533), .B(n156), .Z(\ab[16][54] ) );
  NR2 U3747 ( .A(n534), .B(n156), .Z(\ab[16][53] ) );
  NR2 U3748 ( .A(n535), .B(n156), .Z(\ab[16][52] ) );
  NR2 U3749 ( .A(n536), .B(n156), .Z(\ab[16][51] ) );
  NR2 U3750 ( .A(n537), .B(n156), .Z(\ab[16][50] ) );
  NR2 U3751 ( .A(n538), .B(n156), .Z(\ab[16][49] ) );
  NR2 U3752 ( .A(n539), .B(n156), .Z(\ab[16][48] ) );
  NR2 U3753 ( .A(n540), .B(n157), .Z(\ab[16][47] ) );
  NR2 U3754 ( .A(n541), .B(n157), .Z(\ab[16][46] ) );
  NR2 U3755 ( .A(n542), .B(n157), .Z(\ab[16][45] ) );
  NR2 U3756 ( .A(n543), .B(n157), .Z(\ab[16][44] ) );
  NR2 U3757 ( .A(n544), .B(n157), .Z(\ab[16][43] ) );
  NR2 U3758 ( .A(n545), .B(n157), .Z(\ab[16][42] ) );
  NR2 U3759 ( .A(n546), .B(n157), .Z(\ab[16][41] ) );
  NR2 U3760 ( .A(n547), .B(n157), .Z(\ab[16][40] ) );
  NR2 U3761 ( .A(n548), .B(n157), .Z(\ab[16][39] ) );
  NR2 U3762 ( .A(n492), .B(n5), .Z(\ab[15][95] ) );
  NR2 U3763 ( .A(n493), .B(n5), .Z(\ab[15][94] ) );
  NR2 U3764 ( .A(n494), .B(n5), .Z(\ab[15][93] ) );
  NR2 U3765 ( .A(n495), .B(n5), .Z(\ab[15][92] ) );
  NR2 U3766 ( .A(n496), .B(n5), .Z(\ab[15][91] ) );
  NR2 U3767 ( .A(n497), .B(n5), .Z(\ab[15][90] ) );
  NR2 U3768 ( .A(n498), .B(n5), .Z(\ab[15][89] ) );
  NR2 U3769 ( .A(n499), .B(n5), .Z(\ab[15][88] ) );
  NR2 U3770 ( .A(n500), .B(n5), .Z(\ab[15][87] ) );
  NR2 U3771 ( .A(n501), .B(n5), .Z(\ab[15][86] ) );
  NR2 U3772 ( .A(n502), .B(n5), .Z(\ab[15][85] ) );
  NR2 U3773 ( .A(n503), .B(n5), .Z(\ab[15][84] ) );
  NR2 U3774 ( .A(n504), .B(n6), .Z(\ab[15][83] ) );
  NR2 U3775 ( .A(n505), .B(n6), .Z(\ab[15][82] ) );
  NR2 U3776 ( .A(n506), .B(n6), .Z(\ab[15][81] ) );
  NR2 U3777 ( .A(n507), .B(n6), .Z(\ab[15][80] ) );
  NR2 U3778 ( .A(n508), .B(n6), .Z(\ab[15][79] ) );
  NR2 U3779 ( .A(n509), .B(n6), .Z(\ab[15][78] ) );
  NR2 U3780 ( .A(n510), .B(n6), .Z(\ab[15][77] ) );
  NR2 U3781 ( .A(n511), .B(n6), .Z(\ab[15][76] ) );
  NR2 U3782 ( .A(n512), .B(n6), .Z(\ab[15][75] ) );
  NR2 U3783 ( .A(n513), .B(n6), .Z(\ab[15][74] ) );
  NR2 U3784 ( .A(n514), .B(n6), .Z(\ab[15][73] ) );
  NR2 U3785 ( .A(n515), .B(n6), .Z(\ab[15][72] ) );
  NR2 U3786 ( .A(n516), .B(n7), .Z(\ab[15][71] ) );
  NR2 U3787 ( .A(n517), .B(n7), .Z(\ab[15][70] ) );
  NR2 U3788 ( .A(n518), .B(n7), .Z(\ab[15][69] ) );
  NR2 U3789 ( .A(n519), .B(n7), .Z(\ab[15][68] ) );
  NR2 U3790 ( .A(n520), .B(n7), .Z(\ab[15][67] ) );
  NR2 U3791 ( .A(n521), .B(n7), .Z(\ab[15][66] ) );
  NR2 U3792 ( .A(n522), .B(n7), .Z(\ab[15][65] ) );
  NR2 U3793 ( .A(n523), .B(n7), .Z(\ab[15][64] ) );
  NR2 U3794 ( .A(n524), .B(n7), .Z(\ab[15][63] ) );
  NR2 U3795 ( .A(n525), .B(n7), .Z(\ab[15][62] ) );
  NR2 U3796 ( .A(n526), .B(n7), .Z(\ab[15][61] ) );
  NR2 U3797 ( .A(n527), .B(n7), .Z(\ab[15][60] ) );
  NR2 U3798 ( .A(n528), .B(n8), .Z(\ab[15][59] ) );
  NR2 U3799 ( .A(n529), .B(n8), .Z(\ab[15][58] ) );
  NR2 U3800 ( .A(n530), .B(n8), .Z(\ab[15][57] ) );
  NR2 U3801 ( .A(n531), .B(n8), .Z(\ab[15][56] ) );
  NR2 U3802 ( .A(n532), .B(n8), .Z(\ab[15][55] ) );
  NR2 U3803 ( .A(n533), .B(n8), .Z(\ab[15][54] ) );
  NR2 U3804 ( .A(n534), .B(n8), .Z(\ab[15][53] ) );
  NR2 U3805 ( .A(n535), .B(n8), .Z(\ab[15][52] ) );
  NR2 U3806 ( .A(n536), .B(n8), .Z(\ab[15][51] ) );
  NR2 U3807 ( .A(n537), .B(n8), .Z(\ab[15][50] ) );
  NR2 U3808 ( .A(n538), .B(n8), .Z(\ab[15][49] ) );
  NR2 U3809 ( .A(n539), .B(n8), .Z(\ab[15][48] ) );
  NR2 U3810 ( .A(n540), .B(n9), .Z(\ab[15][47] ) );
  NR2 U3811 ( .A(n541), .B(n9), .Z(\ab[15][46] ) );
  NR2 U3812 ( .A(n542), .B(n9), .Z(\ab[15][45] ) );
  NR2 U3813 ( .A(n543), .B(n9), .Z(\ab[15][44] ) );
  NR2 U3814 ( .A(n544), .B(n9), .Z(\ab[15][43] ) );
  NR2 U3815 ( .A(n545), .B(n9), .Z(\ab[15][42] ) );
  NR2 U3816 ( .A(n546), .B(n9), .Z(\ab[15][41] ) );
  NR2 U3817 ( .A(n547), .B(n9), .Z(\ab[15][40] ) );
  NR2 U3818 ( .A(n548), .B(n9), .Z(\ab[15][39] ) );
endmodule


module LOG_POLY_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:0] carry;

  EO3P U2_6 ( .A(A[6]), .B(n3), .C(carry[6]), .Z(DIFF[6]) );
  FA1A U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1A U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1A U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1A U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA1A U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  IVP U1 ( .A(A[0]), .Z(n1) );
  EN U2 ( .A(A[0]), .B(n9), .Z(DIFF[0]) );
  IVP U3 ( .A(B[1]), .Z(n8) );
  ND2 U4 ( .A(n1), .B(n2), .Z(carry[1]) );
  IVP U5 ( .A(n9), .Z(n2) );
  IVP U6 ( .A(B[2]), .Z(n7) );
  IVP U7 ( .A(B[3]), .Z(n6) );
  IVP U8 ( .A(B[4]), .Z(n5) );
  IVP U9 ( .A(B[5]), .Z(n4) );
  IVP U10 ( .A(B[6]), .Z(n3) );
  IVP U11 ( .A(B[0]), .Z(n9) );
endmodule


module LOG_POLY_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [24:0] carry;

  FA1A U2_22 ( .A(A[22]), .B(n3), .CI(carry[22]), .CO(carry[23]), .S(DIFF[22])
         );
  FA1A U2_21 ( .A(A[21]), .B(n4), .CI(carry[21]), .CO(carry[22]), .S(DIFF[21])
         );
  FA1A U2_20 ( .A(A[20]), .B(n5), .CI(carry[20]), .CO(carry[21]), .S(DIFF[20])
         );
  FA1A U2_19 ( .A(A[19]), .B(n6), .CI(carry[19]), .CO(carry[20]), .S(DIFF[19])
         );
  FA1A U2_18 ( .A(A[18]), .B(n7), .CI(carry[18]), .CO(carry[19]), .S(DIFF[18])
         );
  FA1A U2_17 ( .A(A[17]), .B(n8), .CI(carry[17]), .CO(carry[18]), .S(DIFF[17])
         );
  FA1A U2_16 ( .A(A[16]), .B(n9), .CI(carry[16]), .CO(carry[17]), .S(DIFF[16])
         );
  FA1A U2_15 ( .A(A[15]), .B(n10), .CI(carry[15]), .CO(carry[16]), .S(DIFF[15]) );
  FA1A U2_14 ( .A(A[14]), .B(n11), .CI(carry[14]), .CO(carry[15]), .S(DIFF[14]) );
  FA1A U2_13 ( .A(A[13]), .B(n12), .CI(carry[13]), .CO(carry[14]), .S(DIFF[13]) );
  FA1A U2_12 ( .A(A[12]), .B(n13), .CI(carry[12]), .CO(carry[13]), .S(DIFF[12]) );
  FA1A U2_11 ( .A(A[11]), .B(n14), .CI(carry[11]), .CO(carry[12]), .S(DIFF[11]) );
  FA1A U2_10 ( .A(A[10]), .B(n15), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  FA1A U2_9 ( .A(A[9]), .B(n16), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]) );
  FA1A U2_8 ( .A(A[8]), .B(n17), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA1A U2_7 ( .A(A[7]), .B(n18), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA1A U2_6 ( .A(A[6]), .B(n19), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1A U2_5 ( .A(A[5]), .B(n20), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1A U2_4 ( .A(A[4]), .B(n21), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1A U2_3 ( .A(A[3]), .B(n22), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1A U2_2 ( .A(A[2]), .B(n23), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA1A U2_1 ( .A(A[1]), .B(n24), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  EN U1 ( .A(A[23]), .B(carry[23]), .Z(DIFF[23]) );
  IVP U2 ( .A(n25), .Z(n2) );
  IVP U3 ( .A(B[0]), .Z(n25) );
  ND2 U4 ( .A(n1), .B(n2), .Z(carry[1]) );
  IVP U5 ( .A(B[1]), .Z(n24) );
  IVP U6 ( .A(A[0]), .Z(n1) );
  IVP U7 ( .A(B[2]), .Z(n23) );
  IVP U8 ( .A(B[3]), .Z(n22) );
  IVP U9 ( .A(B[4]), .Z(n21) );
  IVP U10 ( .A(B[5]), .Z(n20) );
  IVP U11 ( .A(B[6]), .Z(n19) );
  IVP U12 ( .A(B[7]), .Z(n18) );
  IVP U13 ( .A(B[8]), .Z(n17) );
  IVP U14 ( .A(B[9]), .Z(n16) );
  IVP U15 ( .A(B[10]), .Z(n15) );
  IVP U16 ( .A(B[11]), .Z(n14) );
  IVP U17 ( .A(B[12]), .Z(n13) );
  IVP U18 ( .A(B[13]), .Z(n12) );
  IVP U19 ( .A(B[14]), .Z(n11) );
  IVP U20 ( .A(B[15]), .Z(n10) );
  IVP U21 ( .A(B[16]), .Z(n9) );
  IVP U22 ( .A(B[17]), .Z(n8) );
  IVP U23 ( .A(B[18]), .Z(n7) );
  IVP U24 ( .A(B[19]), .Z(n6) );
  IVP U25 ( .A(B[20]), .Z(n5) );
  IVP U26 ( .A(B[21]), .Z(n4) );
  IVP U27 ( .A(B[22]), .Z(n3) );
  EN U28 ( .A(A[0]), .B(n25), .Z(DIFF[0]) );
endmodule


module LOG_POLY_DW01_add_5 ( A, B, CI, SUM, CO );
  input [93:0] A;
  input [93:0] B;
  output [93:0] SUM;
  input CI;
  output CO;
  wire   \A[46] , \A[45] , \A[44] , \A[43] , \A[42] , \A[41] , \A[40] ,
         \A[39] , \A[38] , \A[37] , \A[36] , \A[35] , \A[34] , \A[33] ,
         \A[32] , \A[31] , \A[30] , \A[29] , \A[28] , \A[27] , \A[26] ,
         \A[25] , \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] ,
         \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] ,
         \A[11] , \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] ,
         \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467;
  assign SUM[46] = \A[46] ;
  assign \A[46]  = A[46];
  assign SUM[45] = \A[45] ;
  assign \A[45]  = A[45];
  assign SUM[44] = \A[44] ;
  assign \A[44]  = A[44];
  assign SUM[43] = \A[43] ;
  assign \A[43]  = A[43];
  assign SUM[42] = \A[42] ;
  assign \A[42]  = A[42];
  assign SUM[41] = \A[41] ;
  assign \A[41]  = A[41];
  assign SUM[40] = \A[40] ;
  assign \A[40]  = A[40];
  assign SUM[39] = \A[39] ;
  assign \A[39]  = A[39];
  assign SUM[38] = \A[38] ;
  assign \A[38]  = A[38];
  assign SUM[37] = \A[37] ;
  assign \A[37]  = A[37];
  assign SUM[36] = \A[36] ;
  assign \A[36]  = A[36];
  assign SUM[35] = \A[35] ;
  assign \A[35]  = A[35];
  assign SUM[34] = \A[34] ;
  assign \A[34]  = A[34];
  assign SUM[33] = \A[33] ;
  assign \A[33]  = A[33];
  assign SUM[32] = \A[32] ;
  assign \A[32]  = A[32];
  assign SUM[31] = \A[31] ;
  assign \A[31]  = A[31];
  assign SUM[30] = \A[30] ;
  assign \A[30]  = A[30];
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AO4 U2 ( .A(A[55]), .B(B[55]), .C(A[54]), .D(B[54]), .Z(n338) );
  B5I U3 ( .A(n299), .Z(n177) );
  IVDA U4 ( .A(A[72]), .Z(n1) );
  IVP U5 ( .A(n259), .Z(n2) );
  IVP U6 ( .A(n316), .Z(n172) );
  ND4 U7 ( .A(n412), .B(n413), .C(n343), .D(n414), .Z(n325) );
  AO3P U8 ( .A(n208), .B(n209), .C(n210), .D(n211), .Z(n195) );
  IVA U9 ( .A(n193), .Z(n208) );
  AO3P U10 ( .A(n338), .B(n339), .C(n340), .D(n341), .Z(n337) );
  ND2 U11 ( .A(B[60]), .B(A[60]), .Z(n352) );
  ND2P U12 ( .A(n417), .B(n412), .Z(n340) );
  B5I U13 ( .A(n382), .Z(n362) );
  AN2P U14 ( .A(n50), .B(n57), .Z(n101) );
  ND2 U15 ( .A(n147), .B(n148), .Z(n142) );
  IVP U16 ( .A(n236), .Z(n235) );
  IVP U17 ( .A(n311), .Z(n309) );
  AN2 U18 ( .A(n108), .B(n109), .Z(n103) );
  AO3P U19 ( .A(n347), .B(n348), .C(n349), .D(n350), .Z(n346) );
  IVP U20 ( .A(n282), .Z(n281) );
  B5I U21 ( .A(n170), .Z(n114) );
  IV U22 ( .A(n223), .Z(n222) );
  AO7 U23 ( .A(n294), .B(n198), .C(n197), .Z(n268) );
  IV U24 ( .A(n245), .Z(n244) );
  ND2 U25 ( .A(n342), .B(n343), .Z(n339) );
  IVDAP U26 ( .A(n213), .Y(n4), .Z(n3) );
  ND2P U27 ( .A(n370), .B(n371), .Z(n364) );
  NR2P U28 ( .A(n65), .B(n66), .Z(n108) );
  ND4P U29 ( .A(n332), .B(n333), .C(n334), .D(n335), .Z(n331) );
  ND2P U30 ( .A(n308), .B(n180), .Z(n307) );
  B5I U31 ( .A(n466), .Z(n335) );
  AN2 U32 ( .A(n204), .B(n205), .Z(n6) );
  ENP U33 ( .A(n3), .B(n19), .Z(SUM[78]) );
  IV U34 ( .A(n268), .Z(n290) );
  B5I U35 ( .A(n322), .Z(n411) );
  IVDA U36 ( .A(A[84]), .Y(n139) );
  NR2 U37 ( .A(n324), .B(n325), .Z(n323) );
  IVAP U38 ( .A(A[87]), .Z(n100) );
  IVA U39 ( .A(B[87]), .Z(n99) );
  ND3P U40 ( .A(n301), .B(n361), .C(n302), .Z(n316) );
  B5I U41 ( .A(n128), .Z(n127) );
  ND2P U42 ( .A(n116), .B(n106), .Z(n50) );
  ND3P U43 ( .A(n131), .B(n132), .C(n133), .Z(n126) );
  NR2P U44 ( .A(A[64]), .B(B[64]), .Z(n8) );
  IV U45 ( .A(n88), .Z(n90) );
  ND2P U46 ( .A(n393), .B(n379), .Z(n406) );
  NR2P U47 ( .A(n325), .B(n331), .Z(n326) );
  ENP U48 ( .A(n279), .B(n278), .Z(SUM[70]) );
  AN2 U49 ( .A(n15), .B(n85), .Z(n17) );
  AO7P U50 ( .A(n94), .B(n95), .C(n96), .Z(n88) );
  IVA U51 ( .A(n93), .Z(n94) );
  IV U52 ( .A(n74), .Z(n76) );
  AO7P U53 ( .A(n79), .B(n13), .C(n80), .Z(n74) );
  ND3 U54 ( .A(n140), .B(n141), .C(n142), .Z(n133) );
  IV U55 ( .A(n197), .Z(n178) );
  ND2 U56 ( .A(n155), .B(n149), .Z(n147) );
  ND2 U57 ( .A(n156), .B(n157), .Z(n155) );
  IV U58 ( .A(B[82]), .Z(n152) );
  NR3 U59 ( .A(n196), .B(n178), .C(n66), .Z(n185) );
  ND4 U60 ( .A(n191), .B(n192), .C(n193), .D(n190), .Z(n176) );
  ND2 U61 ( .A(n391), .B(n392), .Z(n356) );
  NR2 U62 ( .A(A[50]), .B(B[50]), .Z(n444) );
  ND2 U63 ( .A(n55), .B(n56), .Z(n54) );
  NR2 U64 ( .A(n380), .B(n381), .Z(n378) );
  AO6 U65 ( .A(n249), .B(n238), .C(n250), .Z(n248) );
  IVP U66 ( .A(n8), .Z(n305) );
  ND2 U67 ( .A(B[56]), .B(A[56]), .Z(n359) );
  EN U68 ( .A(n117), .B(n42), .Z(SUM[86]) );
  EN U69 ( .A(n422), .B(n423), .Z(SUM[55]) );
  EO U70 ( .A(n43), .B(B[93]), .Z(SUM[93]) );
  AO3 U71 ( .A(n58), .B(n59), .C(n60), .D(n12), .Z(n44) );
  EN U72 ( .A(n70), .B(n18), .Z(SUM[87]) );
  EO U73 ( .A(n260), .B(n261), .Z(SUM[72]) );
  EN U74 ( .A(n255), .B(n256), .Z(SUM[73]) );
  EN U75 ( .A(n226), .B(n20), .Z(SUM[76]) );
  EN U76 ( .A(n221), .B(n21), .Z(SUM[77]) );
  EO U77 ( .A(n292), .B(n293), .Z(SUM[68]) );
  EO U78 ( .A(n383), .B(n384), .Z(SUM[60]) );
  NR2 U79 ( .A(n385), .B(n380), .Z(n384) );
  EO U80 ( .A(n449), .B(n450), .Z(SUM[51]) );
  EN U81 ( .A(n136), .B(n137), .Z(SUM[84]) );
  EN U82 ( .A(n145), .B(n35), .Z(SUM[83]) );
  EN U83 ( .A(n129), .B(n36), .Z(SUM[85]) );
  EN U84 ( .A(n158), .B(n40), .Z(SUM[81]) );
  EN U85 ( .A(n151), .B(n41), .Z(SUM[82]) );
  AN2P U86 ( .A(n375), .B(n352), .Z(n5) );
  ND3 U87 ( .A(n351), .B(n352), .C(n353), .Z(n169) );
  AN2P U88 ( .A(n420), .B(n421), .Z(n7) );
  IVAP U89 ( .A(A[62]), .Z(n373) );
  IVP U90 ( .A(n107), .Z(n105) );
  IV U91 ( .A(B[51]), .Z(n451) );
  AO6P U92 ( .A(n368), .B(n363), .C(n369), .Z(n367) );
  AO7P U93 ( .A(n243), .B(n244), .C(n233), .Z(n240) );
  IVAP U94 ( .A(n415), .Z(n409) );
  ND2 U95 ( .A(n315), .B(n287), .Z(n314) );
  ND2P U96 ( .A(n61), .B(n62), .Z(n104) );
  NR2P U97 ( .A(n441), .B(n442), .Z(n440) );
  NR3P U98 ( .A(n443), .B(n444), .C(n445), .Z(n442) );
  ND2P U99 ( .A(n127), .B(n124), .Z(n107) );
  IVDA U100 ( .A(n266), .Z(n9) );
  B3I U101 ( .A(n202), .Z1(n11), .Z2(n10) );
  IVP U102 ( .A(A[81]), .Z(n160) );
  OR2P U103 ( .A(n134), .B(n135), .Z(n128) );
  AO6 U104 ( .A(n188), .B(n176), .C(n189), .Z(n187) );
  ND2P U105 ( .A(n365), .B(n353), .Z(n301) );
  IV U106 ( .A(n252), .Z(n249) );
  ND2P U107 ( .A(B[71]), .B(A[71]), .Z(n263) );
  OR2P U108 ( .A(n329), .B(n24), .Z(n415) );
  AN2 U109 ( .A(n17), .B(n78), .Z(n16) );
  AO7P U110 ( .A(n208), .B(n4), .C(n211), .Z(n212) );
  ND2P U111 ( .A(n265), .B(n266), .Z(n262) );
  NR2 U112 ( .A(n328), .B(n329), .Z(n327) );
  AO3 U113 ( .A(A[50]), .B(B[50]), .C(n436), .D(n437), .Z(n329) );
  OR2P U114 ( .A(B[61]), .B(A[61]), .Z(n374) );
  IV U115 ( .A(n258), .Z(n257) );
  ND2P U116 ( .A(n217), .B(n192), .Z(n216) );
  IV U117 ( .A(n338), .Z(n419) );
  IV U118 ( .A(n198), .Z(n196) );
  OR2P U119 ( .A(n66), .B(n174), .Z(n225) );
  OR2P U120 ( .A(n259), .B(n66), .Z(n254) );
  ND4P U121 ( .A(n203), .B(n266), .C(n265), .D(n267), .Z(n66) );
  NR3P U122 ( .A(n174), .B(n234), .C(n235), .Z(n227) );
  IV U123 ( .A(n239), .Z(n259) );
  OR2P U124 ( .A(A[59]), .B(B[59]), .Z(n330) );
  AO7P U125 ( .A(n403), .B(n14), .C(n357), .Z(n400) );
  AN2P U126 ( .A(n359), .B(n405), .Z(n14) );
  ND2P U127 ( .A(n122), .B(n123), .Z(n116) );
  AO7P U128 ( .A(n431), .B(n432), .C(n420), .Z(n429) );
  IV U129 ( .A(n433), .Z(n432) );
  IVP U130 ( .A(n304), .Z(n361) );
  IVAP U131 ( .A(A[60]), .Z(n395) );
  IVP U132 ( .A(B[60]), .Z(n394) );
  ND2 U133 ( .A(n224), .B(n191), .Z(n220) );
  IVAP U134 ( .A(n374), .Z(n365) );
  AN2P U135 ( .A(n86), .B(n87), .Z(n13) );
  IV U136 ( .A(B[84]), .Z(n138) );
  AN2P U137 ( .A(n72), .B(n73), .Z(n25) );
  IVP U138 ( .A(A[56]), .Z(n408) );
  OR2 U139 ( .A(B[89]), .B(A[89]), .Z(n85) );
  AO7 U140 ( .A(n48), .B(n25), .C(n49), .Z(n47) );
  IVAP U141 ( .A(n163), .Z(n120) );
  AO7P U142 ( .A(n365), .B(n5), .C(n351), .Z(n368) );
  ND2P U143 ( .A(n263), .B(n264), .Z(n202) );
  AO7P U144 ( .A(n6), .B(n262), .C(n11), .Z(n236) );
  IV U145 ( .A(n251), .Z(n250) );
  ND3P U146 ( .A(n321), .B(n322), .C(n323), .Z(n113) );
  ND2P U147 ( .A(n110), .B(n113), .Z(n270) );
  AO7P U148 ( .A(n270), .B(n271), .C(n272), .Z(n269) );
  IV U149 ( .A(n335), .Z(n24) );
  IV U150 ( .A(n330), .Z(n328) );
  IVAP U151 ( .A(n461), .Z(n438) );
  OR2P U152 ( .A(B[76]), .B(A[76]), .Z(n191) );
  OR2P U153 ( .A(B[77]), .B(A[77]), .Z(n192) );
  NR3P U154 ( .A(n174), .B(n175), .C(n176), .Z(n173) );
  AO3P U155 ( .A(n228), .B(n229), .C(n230), .D(n231), .Z(n183) );
  OR2P U156 ( .A(B[78]), .B(A[78]), .Z(n193) );
  OR2P U157 ( .A(B[79]), .B(A[79]), .Z(n190) );
  ND3P U158 ( .A(n351), .B(n362), .C(n353), .Z(n302) );
  IV U159 ( .A(B[81]), .Z(n159) );
  IVP U160 ( .A(A[82]), .Z(n153) );
  OR2P U161 ( .A(B[66]), .B(A[66]), .Z(n180) );
  OR2P U162 ( .A(B[67]), .B(A[67]), .Z(n197) );
  OR2P U163 ( .A(B[83]), .B(A[83]), .Z(n140) );
  ND2P U164 ( .A(n394), .B(n395), .Z(n382) );
  OR2P U165 ( .A(B[68]), .B(A[68]), .Z(n267) );
  OR2P U166 ( .A(B[88]), .B(A[88]), .Z(n93) );
  IV U167 ( .A(B[56]), .Z(n407) );
  AN2 U168 ( .A(B[72]), .B(n1), .Z(n28) );
  ND2P U169 ( .A(n99), .B(n100), .Z(n92) );
  OR2P U170 ( .A(B[85]), .B(A[85]), .Z(n124) );
  ND2P U171 ( .A(n118), .B(n119), .Z(n106) );
  ND2P U172 ( .A(n372), .B(n373), .Z(n363) );
  IVP U173 ( .A(n57), .Z(n55) );
  OR2P U174 ( .A(B[91]), .B(A[91]), .Z(n71) );
  IVP U175 ( .A(B[63]), .Z(n370) );
  IVA U176 ( .A(n467), .Z(SUM[47]) );
  OR2P U177 ( .A(B[92]), .B(A[92]), .Z(n56) );
  ENP U178 ( .A(n212), .B(n38), .Z(SUM[79]) );
  ENP U179 ( .A(n240), .B(n37), .Z(SUM[75]) );
  ENP U180 ( .A(n306), .B(n39), .Z(SUM[67]) );
  EOP U181 ( .A(n367), .B(n366), .Z(SUM[63]) );
  ENP U182 ( .A(n274), .B(n34), .Z(SUM[71]) );
  ENP U183 ( .A(n81), .B(n31), .Z(SUM[90]) );
  ENP U184 ( .A(n75), .B(n32), .Z(SUM[91]) );
  ENP U185 ( .A(n67), .B(n33), .Z(SUM[92]) );
  ENP U186 ( .A(n97), .B(n29), .Z(SUM[88]) );
  ENP U187 ( .A(n89), .B(n30), .Z(SUM[89]) );
  AO7 U188 ( .A(n120), .B(n107), .C(n121), .Z(n117) );
  ND2 U189 ( .A(n13), .B(n84), .Z(n81) );
  ND2 U190 ( .A(n17), .B(n70), .Z(n84) );
  ND2 U191 ( .A(n76), .B(n77), .Z(n75) );
  ND2 U192 ( .A(n16), .B(n70), .Z(n77) );
  ND4 U193 ( .A(n349), .B(n358), .C(n359), .D(n357), .Z(n386) );
  ND2 U194 ( .A(n219), .B(n192), .Z(n215) );
  ND2 U195 ( .A(n166), .B(n64), .Z(n165) );
  IV U196 ( .A(n359), .Z(n354) );
  ND2 U197 ( .A(n357), .B(n358), .Z(n355) );
  AN2P U198 ( .A(n105), .B(n106), .Z(n12) );
  AO7 U199 ( .A(n161), .B(n120), .C(n162), .Z(n158) );
  AO7 U200 ( .A(n120), .B(n154), .C(n147), .Z(n151) );
  ND2 U201 ( .A(n376), .B(n377), .Z(n375) );
  IVP U202 ( .A(n346), .Z(n273) );
  IVA U203 ( .A(n169), .Z(n350) );
  ND2 U204 ( .A(n25), .B(n68), .Z(n67) );
  ND2 U205 ( .A(n69), .B(n70), .Z(n68) );
  ND3 U206 ( .A(n181), .B(n182), .C(n183), .Z(n61) );
  ND2 U207 ( .A(n236), .B(n203), .Z(n258) );
  AN2P U208 ( .A(n92), .B(n93), .Z(n15) );
  NR2 U209 ( .A(n288), .B(n289), .Z(n286) );
  ND2 U210 ( .A(n92), .B(n95), .Z(n18) );
  ND2 U211 ( .A(n264), .B(n9), .Z(n279) );
  EN U212 ( .A(n246), .B(n245), .Z(SUM[74]) );
  ND2 U213 ( .A(n233), .B(n237), .Z(n246) );
  ND2 U214 ( .A(n193), .B(n211), .Z(n19) );
  EO U215 ( .A(n400), .B(n401), .Z(SUM[58]) );
  NR2 U216 ( .A(n402), .B(n391), .Z(n401) );
  NR2 U217 ( .A(n259), .B(n28), .Z(n261) );
  ND2 U218 ( .A(n238), .B(n251), .Z(n256) );
  ND2 U219 ( .A(n191), .B(n194), .Z(n20) );
  ND2 U220 ( .A(n192), .B(n209), .Z(n21) );
  EN U221 ( .A(n164), .B(n163), .Z(SUM[80]) );
  EO U222 ( .A(n404), .B(n14), .Z(SUM[57]) );
  EO U223 ( .A(n5), .B(n22), .Z(SUM[61]) );
  ND2 U224 ( .A(n374), .B(n351), .Z(n22) );
  ND2 U225 ( .A(n267), .B(n204), .Z(n292) );
  EN U226 ( .A(n283), .B(n282), .Z(SUM[69]) );
  EN U227 ( .A(n406), .B(n23), .Z(SUM[56]) );
  ND2 U228 ( .A(n333), .B(n359), .Z(n23) );
  ND2 U229 ( .A(n455), .B(n456), .Z(n454) );
  EN U230 ( .A(n434), .B(n433), .Z(SUM[52]) );
  ND2 U231 ( .A(n420), .B(n414), .Z(n434) );
  EN U232 ( .A(n457), .B(n455), .Z(SUM[50]) );
  ND2 U233 ( .A(n453), .B(n456), .Z(n457) );
  IV U234 ( .A(B[75]), .Z(n241) );
  IVP U235 ( .A(B[90]), .Z(n82) );
  ND2 U236 ( .A(B[80]), .B(A[80]), .Z(n157) );
  ND2 U237 ( .A(n435), .B(n415), .Z(n433) );
  ND2 U238 ( .A(B[81]), .B(A[81]), .Z(n156) );
  IV U239 ( .A(B[71]), .Z(n275) );
  IV U240 ( .A(A[71]), .Z(n276) );
  ND2 U241 ( .A(B[72]), .B(n1), .Z(n229) );
  AO3 U242 ( .A(n7), .B(n416), .C(n341), .D(n340), .Z(n381) );
  ND2 U243 ( .A(B[74]), .B(A[74]), .Z(n233) );
  ND2 U244 ( .A(B[78]), .B(A[78]), .Z(n211) );
  ND4 U245 ( .A(n301), .B(n197), .C(n302), .D(n303), .Z(n289) );
  ND2 U246 ( .A(B[59]), .B(A[59]), .Z(n349) );
  ND2 U247 ( .A(B[58]), .B(A[58]), .Z(n358) );
  ND2 U248 ( .A(B[59]), .B(A[59]), .Z(n392) );
  ND2 U249 ( .A(B[82]), .B(A[82]), .Z(n148) );
  ND2 U250 ( .A(B[88]), .B(A[88]), .Z(n96) );
  ND2 U251 ( .A(B[90]), .B(A[90]), .Z(n80) );
  ND2 U252 ( .A(B[89]), .B(A[89]), .Z(n87) );
  ND2 U253 ( .A(B[51]), .B(A[51]), .Z(n446) );
  ND4 U254 ( .A(n387), .B(n388), .C(n389), .D(n390), .Z(n360) );
  IV U255 ( .A(B[57]), .Z(n390) );
  ND2 U256 ( .A(B[58]), .B(A[58]), .Z(n388) );
  AO7 U257 ( .A(n201), .B(n10), .C(n203), .Z(n200) );
  NR2 U258 ( .A(n48), .B(n53), .Z(n60) );
  ND2 U259 ( .A(B[75]), .B(A[75]), .Z(n232) );
  ND2 U260 ( .A(B[59]), .B(A[59]), .Z(n387) );
  EN U261 ( .A(n308), .B(n26), .Z(SUM[66]) );
  ND2 U262 ( .A(n180), .B(n296), .Z(n26) );
  EN U263 ( .A(n368), .B(n27), .Z(SUM[62]) );
  ND2 U264 ( .A(n363), .B(n353), .Z(n27) );
  EN U265 ( .A(n426), .B(n425), .Z(SUM[54]) );
  ND2 U266 ( .A(B[52]), .B(A[52]), .Z(n420) );
  ND2 U267 ( .A(B[77]), .B(A[77]), .Z(n209) );
  ND2 U268 ( .A(B[83]), .B(A[83]), .Z(n132) );
  ND2 U269 ( .A(B[66]), .B(A[66]), .Z(n296) );
  ND2 U270 ( .A(B[76]), .B(A[76]), .Z(n194) );
  ND2 U271 ( .A(B[86]), .B(A[86]), .Z(n57) );
  ND2 U272 ( .A(B[79]), .B(A[79]), .Z(n210) );
  ND2 U273 ( .A(B[84]), .B(A[84]), .Z(n131) );
  ND2 U274 ( .A(B[85]), .B(A[85]), .Z(n123) );
  ND2 U275 ( .A(B[67]), .B(A[67]), .Z(n295) );
  IVP U276 ( .A(A[86]), .Z(n119) );
  IVP U277 ( .A(B[86]), .Z(n118) );
  EN U278 ( .A(n430), .B(n429), .Z(SUM[53]) );
  ND2 U279 ( .A(B[49]), .B(A[49]), .Z(n459) );
  ND2 U280 ( .A(B[58]), .B(A[58]), .Z(n399) );
  EN U281 ( .A(n462), .B(n460), .Z(SUM[49]) );
  ND2 U282 ( .A(B[80]), .B(A[80]), .Z(n162) );
  ND2 U283 ( .A(B[50]), .B(A[50]), .Z(n453) );
  ND2 U284 ( .A(B[50]), .B(A[50]), .Z(n447) );
  ND2 U285 ( .A(n344), .B(n345), .Z(n342) );
  ND2 U286 ( .A(B[52]), .B(A[52]), .Z(n344) );
  ND2 U287 ( .A(B[53]), .B(A[53]), .Z(n345) );
  NR2 U288 ( .A(n300), .B(n168), .Z(n294) );
  ND2 U289 ( .A(B[53]), .B(A[53]), .Z(n421) );
  ND2 U290 ( .A(n350), .B(n168), .Z(n115) );
  ND2 U291 ( .A(B[91]), .B(A[91]), .Z(n73) );
  IVP U292 ( .A(n56), .Z(n48) );
  EO U293 ( .A(n319), .B(n320), .Z(SUM[64]) );
  EN U294 ( .A(n312), .B(n311), .Z(SUM[65]) );
  ND2 U295 ( .A(n463), .B(n464), .Z(n460) );
  ND2 U296 ( .A(n436), .B(n335), .Z(n464) );
  EN U297 ( .A(n465), .B(n335), .Z(SUM[48]) );
  ND2 U298 ( .A(n436), .B(n463), .Z(n465) );
  ND2 U299 ( .A(B[48]), .B(A[48]), .Z(n443) );
  ND4 U300 ( .A(n295), .B(n296), .C(n297), .D(n298), .Z(n198) );
  ND2 U301 ( .A(B[63]), .B(A[63]), .Z(n168) );
  ND2 U302 ( .A(B[92]), .B(A[92]), .Z(n49) );
  ND2 U303 ( .A(B[48]), .B(A[48]), .Z(n463) );
  ND2 U304 ( .A(B[65]), .B(A[65]), .Z(n310) );
  ND2 U305 ( .A(n93), .B(n96), .Z(n29) );
  ND2 U306 ( .A(n85), .B(n87), .Z(n30) );
  ND2 U307 ( .A(n78), .B(n80), .Z(n31) );
  ND2 U308 ( .A(n71), .B(n73), .Z(n32) );
  ND2 U309 ( .A(n49), .B(n56), .Z(n33) );
  ND2 U310 ( .A(n263), .B(n203), .Z(n34) );
  ND2 U311 ( .A(n132), .B(n140), .Z(n35) );
  ND2 U312 ( .A(n124), .B(n123), .Z(n36) );
  ND2 U313 ( .A(n232), .B(n181), .Z(n37) );
  ND2 U314 ( .A(n364), .B(n168), .Z(n366) );
  ND2 U315 ( .A(n210), .B(n190), .Z(n38) );
  ND2 U316 ( .A(n295), .B(n197), .Z(n39) );
  ND2 U317 ( .A(n156), .B(n149), .Z(n40) );
  ND2 U318 ( .A(n148), .B(n141), .Z(n41) );
  ND2 U319 ( .A(n106), .B(n57), .Z(n42) );
  ND2 U320 ( .A(B[57]), .B(A[57]), .Z(n357) );
  IV U321 ( .A(A[57]), .Z(n389) );
  NR2 U322 ( .A(n300), .B(n304), .Z(n303) );
  ND2 U323 ( .A(n425), .B(n413), .Z(n424) );
  IV U324 ( .A(n176), .Z(n182) );
  NR2 U325 ( .A(n8), .B(n316), .Z(n315) );
  ND2 U326 ( .A(B[64]), .B(A[64]), .Z(n318) );
  ND2 U327 ( .A(n61), .B(n62), .Z(n59) );
  IVDA U328 ( .A(n334), .Y(n403) );
  ND2 U329 ( .A(n357), .B(n334), .Z(n404) );
  ND2 U330 ( .A(B[55]), .B(A[55]), .Z(n341) );
  ND2 U331 ( .A(n150), .B(n149), .Z(n154) );
  IVDA U332 ( .A(n150), .Y(n161) );
  ND2 U333 ( .A(n162), .B(n150), .Z(n164) );
  ND2 U334 ( .A(n412), .B(n341), .Z(n423) );
  ND2 U335 ( .A(B[73]), .B(A[73]), .Z(n251) );
  AO4 U336 ( .A(A[74]), .B(B[74]), .C(A[73]), .D(B[73]), .Z(n228) );
  AO3 U337 ( .A(A[74]), .B(B[74]), .C(A[73]), .D(B[73]), .Z(n230) );
  ND2 U338 ( .A(n273), .B(n170), .Z(n271) );
  ND3 U339 ( .A(A[65]), .B(B[65]), .C(n180), .Z(n298) );
  AO6 U340 ( .A(n171), .B(n305), .C(n317), .Z(n313) );
  ND2 U341 ( .A(n305), .B(n318), .Z(n319) );
  AO7 U342 ( .A(n214), .B(n220), .C(n218), .Z(n221) );
  AO7 U343 ( .A(n214), .B(n225), .C(n223), .Z(n226) );
  AO7 U344 ( .A(n214), .B(n254), .C(n252), .Z(n255) );
  AO7 U345 ( .A(n214), .B(n66), .C(n258), .Z(n260) );
  ND2 U346 ( .A(n382), .B(n352), .Z(n383) );
  ND2 U347 ( .A(n398), .B(n399), .Z(n396) );
  ND2 U348 ( .A(n400), .B(n332), .Z(n398) );
  ND2P U349 ( .A(n284), .B(n285), .Z(n282) );
  ND2 U350 ( .A(B[87]), .B(A[87]), .Z(n95) );
  ND2 U351 ( .A(n90), .B(n91), .Z(n89) );
  ND2 U352 ( .A(n15), .B(n70), .Z(n91) );
  ND2 U353 ( .A(n88), .B(n85), .Z(n86) );
  IV U354 ( .A(n324), .Z(n336) );
  AO7 U355 ( .A(A[47]), .B(B[47]), .C(n466), .Z(n467) );
  ND2 U356 ( .A(n378), .B(n379), .Z(n377) );
  ND2P U357 ( .A(n143), .B(n140), .Z(n135) );
  ND2 U358 ( .A(n205), .B(n265), .Z(n283) );
  AO6 U359 ( .A(n204), .B(n205), .C(n206), .Z(n201) );
  AO4 U360 ( .A(A[69]), .B(B[69]), .C(A[70]), .D(B[70]), .Z(n206) );
  OR2P U361 ( .A(A[69]), .B(B[69]), .Z(n265) );
  IV U362 ( .A(n418), .Z(n417) );
  NR2 U363 ( .A(n207), .B(n195), .Z(n199) );
  IVP U364 ( .A(n195), .Z(n188) );
  IV U365 ( .A(n180), .Z(n179) );
  AO7 U366 ( .A(n438), .B(n458), .C(n459), .Z(n455) );
  AO3 U367 ( .A(A[50]), .B(B[50]), .C(A[49]), .D(B[49]), .Z(n448) );
  NR2 U368 ( .A(A[49]), .B(B[49]), .Z(n445) );
  OR2P U369 ( .A(A[52]), .B(B[52]), .Z(n414) );
  ND2 U370 ( .A(n98), .B(n95), .Z(n97) );
  ND2 U371 ( .A(n92), .B(n70), .Z(n98) );
  AO7 U372 ( .A(n257), .B(n28), .C(n2), .Z(n252) );
  ND2 U373 ( .A(n459), .B(n461), .Z(n462) );
  OR2 U374 ( .A(n48), .B(n53), .Z(n51) );
  ND2 U375 ( .A(n321), .B(n322), .Z(n435) );
  OR2P U376 ( .A(A[54]), .B(B[54]), .Z(n413) );
  NR2 U377 ( .A(n114), .B(n115), .Z(n167) );
  OR2P U378 ( .A(A[53]), .B(B[53]), .Z(n343) );
  OR2P U379 ( .A(A[49]), .B(B[49]), .Z(n461) );
  ND2 U380 ( .A(n74), .B(n71), .Z(n72) );
  AO7 U381 ( .A(n50), .B(n51), .C(n52), .Z(n46) );
  ND2 U382 ( .A(n406), .B(n333), .Z(n405) );
  NR2P U383 ( .A(n411), .B(n438), .Z(n437) );
  IVA U384 ( .A(A[63]), .Z(n371) );
  ND2 U385 ( .A(n418), .B(n424), .Z(n422) );
  ND2 U386 ( .A(n413), .B(n418), .Z(n426) );
  NR2 U387 ( .A(n46), .B(n47), .Z(n45) );
  IV U388 ( .A(n78), .Z(n79) );
  IV U389 ( .A(A[90]), .Z(n83) );
  OR2P U390 ( .A(A[72]), .B(B[72]), .Z(n239) );
  AO7 U391 ( .A(n120), .B(n128), .C(n130), .Z(n129) );
  AO7 U392 ( .A(n120), .B(n144), .C(n146), .Z(n145) );
  ND2 U393 ( .A(n142), .B(n141), .Z(n146) );
  IVP U394 ( .A(n144), .Z(n143) );
  OR2P U395 ( .A(A[70]), .B(B[70]), .Z(n266) );
  IV U396 ( .A(n125), .Z(n134) );
  ND2 U397 ( .A(n131), .B(n125), .Z(n137) );
  ND2 U398 ( .A(n126), .B(n125), .Z(n130) );
  AO3 U399 ( .A(n120), .B(n135), .C(n133), .D(n132), .Z(n136) );
  IV U400 ( .A(A[75]), .Z(n242) );
  IVA U401 ( .A(B[62]), .Z(n372) );
  ND3 U402 ( .A(n194), .B(n174), .C(n188), .Z(n186) );
  OR2P U403 ( .A(A[73]), .B(B[73]), .Z(n238) );
  OR2P U404 ( .A(A[74]), .B(B[74]), .Z(n237) );
  OR2P U405 ( .A(A[55]), .B(B[55]), .Z(n412) );
  OR2P U406 ( .A(A[48]), .B(B[48]), .Z(n436) );
  ND3 U407 ( .A(n124), .B(n125), .C(n126), .Z(n122) );
  IV U408 ( .A(A[51]), .Z(n452) );
  ND2 U409 ( .A(n421), .B(n343), .Z(n430) );
  ND4 U410 ( .A(n110), .B(n111), .C(n167), .D(n113), .Z(n64) );
  ND4 U411 ( .A(n110), .B(n111), .C(n112), .D(n113), .Z(n109) );
  NR2 U412 ( .A(n411), .B(n325), .Z(n410) );
  ND2 U413 ( .A(n343), .B(n419), .Z(n416) );
  ND4P U414 ( .A(n330), .B(n332), .C(n334), .D(n333), .Z(n324) );
  OR2P U415 ( .A(A[57]), .B(B[57]), .Z(n334) );
  OR2P U416 ( .A(A[58]), .B(B[58]), .Z(n332) );
  ND2 U417 ( .A(n310), .B(n299), .Z(n312) );
  NR2 U418 ( .A(n65), .B(n66), .Z(n63) );
  NR2 U419 ( .A(n65), .B(n66), .Z(n166) );
  ND3 U420 ( .A(n299), .B(n305), .C(n180), .Z(n300) );
  ND4 U421 ( .A(B[64]), .B(A[64]), .C(n299), .D(n180), .Z(n297) );
  OR2P U422 ( .A(A[65]), .B(B[65]), .Z(n299) );
  ND2 U423 ( .A(n392), .B(n330), .Z(n397) );
  ND2 U424 ( .A(n278), .B(n9), .Z(n277) );
  AO6 U425 ( .A(n272), .B(n287), .C(n290), .Z(n293) );
  AO6 U426 ( .A(n172), .B(n287), .C(n171), .Z(n320) );
  AO6 U427 ( .A(n393), .B(n379), .C(n324), .Z(n385) );
  ND2 U428 ( .A(n286), .B(n287), .Z(n285) );
  AO6 U429 ( .A(n324), .B(n111), .C(n362), .Z(n376) );
  ND4 U430 ( .A(n356), .B(n360), .C(n330), .D(n386), .Z(n111) );
  ND2 U431 ( .A(n360), .B(n330), .Z(n347) );
  OR2P U432 ( .A(A[80]), .B(B[80]), .Z(n150) );
  ND2 U433 ( .A(n44), .B(n45), .Z(n43) );
  OR2 U434 ( .A(n53), .B(n54), .Z(n52) );
  AN2P U435 ( .A(n63), .B(n64), .Z(n58) );
  IVA U436 ( .A(n53), .Z(n69) );
  ND2P U437 ( .A(n16), .B(n71), .Z(n53) );
  ND2P U438 ( .A(n82), .B(n83), .Z(n78) );
  ND2P U439 ( .A(n101), .B(n102), .Z(n70) );
  AO7P U440 ( .A(n103), .B(n104), .C(n12), .Z(n102) );
  NR2P U441 ( .A(n114), .B(n115), .Z(n112) );
  IVA U442 ( .A(n116), .Z(n121) );
  ND2P U443 ( .A(n138), .B(n139), .Z(n125) );
  ND3P U444 ( .A(n149), .B(n141), .C(n150), .Z(n144) );
  ND2P U445 ( .A(n152), .B(n153), .Z(n141) );
  ND2P U446 ( .A(n159), .B(n160), .Z(n149) );
  ND3P U447 ( .A(n62), .B(n61), .C(n165), .Z(n163) );
  AO7P U448 ( .A(n171), .B(n172), .C(n173), .Z(n65) );
  OR4 U449 ( .A(n177), .B(n8), .C(n178), .D(n179), .Z(n175) );
  AO3P U450 ( .A(n184), .B(n185), .C(n186), .D(n187), .Z(n62) );
  IVA U451 ( .A(n190), .Z(n189) );
  ND2 U452 ( .A(n199), .B(n200), .Z(n184) );
  AO3P U453 ( .A(n214), .B(n215), .C(n216), .D(n209), .Z(n213) );
  IVA U454 ( .A(n218), .Z(n217) );
  IVA U455 ( .A(n220), .Z(n219) );
  AO7P U456 ( .A(n207), .B(n222), .C(n191), .Z(n218) );
  IVA U457 ( .A(n194), .Z(n207) );
  IVA U458 ( .A(n225), .Z(n224) );
  AO7P U459 ( .A(n227), .B(n183), .C(n181), .Z(n223) );
  AN2P U460 ( .A(n232), .B(n233), .Z(n231) );
  IVA U461 ( .A(n203), .Z(n234) );
  ND4P U462 ( .A(n181), .B(n237), .C(n238), .D(n239), .Z(n174) );
  ND2P U463 ( .A(n241), .B(n242), .Z(n181) );
  IVA U464 ( .A(n237), .Z(n243) );
  AO7P U465 ( .A(n214), .B(n247), .C(n248), .Z(n245) );
  ND2 U466 ( .A(n253), .B(n238), .Z(n247) );
  IVA U467 ( .A(n254), .Z(n253) );
  AN2P U468 ( .A(n268), .B(n269), .Z(n214) );
  ND2P U469 ( .A(n275), .B(n276), .Z(n203) );
  ND2 U470 ( .A(n277), .B(n264), .Z(n274) );
  AO7P U471 ( .A(n280), .B(n281), .C(n205), .Z(n278) );
  IVA U472 ( .A(n265), .Z(n280) );
  ND2P U473 ( .A(B[70]), .B(A[70]), .Z(n264) );
  IVA U474 ( .A(n267), .Z(n288) );
  AO6P U475 ( .A(n290), .B(n267), .C(n291), .Z(n284) );
  IVA U476 ( .A(n204), .Z(n291) );
  ND2P U477 ( .A(B[69]), .B(A[69]), .Z(n205) );
  IVA U478 ( .A(n289), .Z(n272) );
  ND2P U479 ( .A(B[68]), .B(A[68]), .Z(n204) );
  ND2 U480 ( .A(n296), .B(n307), .Z(n306) );
  AO7P U481 ( .A(n177), .B(n309), .C(n310), .Z(n308) );
  ND2P U482 ( .A(n313), .B(n314), .Z(n311) );
  IVA U483 ( .A(n318), .Z(n317) );
  IVA U484 ( .A(n168), .Z(n171) );
  ND4P U485 ( .A(n273), .B(n170), .C(n110), .D(n113), .Z(n287) );
  ND2P U486 ( .A(n326), .B(n327), .Z(n110) );
  ND2P U487 ( .A(n336), .B(n337), .Z(n170) );
  AO7P U488 ( .A(n354), .B(n355), .C(n356), .Z(n348) );
  ND2P U489 ( .A(n363), .B(n364), .Z(n304) );
  IVA U490 ( .A(n353), .Z(n369) );
  ND2P U491 ( .A(B[62]), .B(A[62]), .Z(n353) );
  ND2P U492 ( .A(B[61]), .B(A[61]), .Z(n351) );
  IVA U493 ( .A(n111), .Z(n380) );
  ENP U494 ( .A(n396), .B(n397), .Z(SUM[59]) );
  IVA U495 ( .A(n332), .Z(n391) );
  IVA U496 ( .A(n399), .Z(n402) );
  ND2P U497 ( .A(n407), .B(n408), .Z(n333) );
  AO7P U498 ( .A(n409), .B(n321), .C(n410), .Z(n379) );
  IVA U499 ( .A(n381), .Z(n393) );
  AO7P U500 ( .A(n427), .B(n428), .C(n421), .Z(n425) );
  IVA U501 ( .A(n429), .Z(n428) );
  IVA U502 ( .A(n343), .Z(n427) );
  ND2P U503 ( .A(B[54]), .B(A[54]), .Z(n418) );
  IVA U504 ( .A(n414), .Z(n431) );
  ND2P U505 ( .A(n439), .B(n440), .Z(n321) );
  IVA U506 ( .A(n446), .Z(n441) );
  AN2P U507 ( .A(n447), .B(n448), .Z(n439) );
  AN2P U508 ( .A(n446), .B(n322), .Z(n450) );
  ND2P U509 ( .A(n451), .B(n452), .Z(n322) );
  ND2 U510 ( .A(n453), .B(n454), .Z(n449) );
  IVA U511 ( .A(n460), .Z(n458) );
  OR2 U512 ( .A(A[50]), .B(B[50]), .Z(n456) );
  ND2P U513 ( .A(B[47]), .B(A[47]), .Z(n466) );
endmodule


module LOG_POLY_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [47:0] A;
  input [47:0] B;
  output [95:0] PRODUCT;
  input TC;
  wire   \B[0] , \ab[47][47] , \ab[47][45] , \ab[47][44] , \ab[47][43] ,
         \ab[47][42] , \ab[47][41] , \ab[47][40] , \ab[47][39] , \ab[47][38] ,
         \ab[47][37] , \ab[47][36] , \ab[47][35] , \ab[47][34] , \ab[47][33] ,
         \ab[47][32] , \ab[47][31] , \ab[47][30] , \ab[47][29] , \ab[47][28] ,
         \ab[47][27] , \ab[47][26] , \ab[47][25] , \ab[47][24] , \ab[47][23] ,
         \ab[47][22] , \ab[47][21] , \ab[47][20] , \ab[47][19] , \ab[47][18] ,
         \ab[47][17] , \ab[47][16] , \ab[47][15] , \ab[47][14] , \ab[47][13] ,
         \ab[47][12] , \ab[47][11] , \ab[47][10] , \ab[46][46] , \ab[46][45] ,
         \ab[46][44] , \ab[46][43] , \ab[46][42] , \ab[46][41] , \ab[46][40] ,
         \ab[46][39] , \ab[46][38] , \ab[46][37] , \ab[46][36] , \ab[46][35] ,
         \ab[46][34] , \ab[46][33] , \ab[46][32] , \ab[46][31] , \ab[46][30] ,
         \ab[46][29] , \ab[46][28] , \ab[46][27] , \ab[46][26] , \ab[46][25] ,
         \ab[46][24] , \ab[46][23] , \ab[46][22] , \ab[46][21] , \ab[46][20] ,
         \ab[46][19] , \ab[46][18] , \ab[46][17] , \ab[46][16] , \ab[46][15] ,
         \ab[46][14] , \ab[46][13] , \ab[46][12] , \ab[46][11] , \ab[46][10] ,
         \ab[45][45] , \ab[45][44] , \ab[45][43] , \ab[45][42] , \ab[45][41] ,
         \ab[45][40] , \ab[45][39] , \ab[45][38] , \ab[45][37] , \ab[45][36] ,
         \ab[45][35] , \ab[45][34] , \ab[45][33] , \ab[45][32] , \ab[45][31] ,
         \ab[45][30] , \ab[45][29] , \ab[45][28] , \ab[45][27] , \ab[45][26] ,
         \ab[45][25] , \ab[45][24] , \ab[45][23] , \ab[45][22] , \ab[45][21] ,
         \ab[45][20] , \ab[45][19] , \ab[45][18] , \ab[45][17] , \ab[45][16] ,
         \ab[45][15] , \ab[45][14] , \ab[45][13] , \ab[45][12] , \ab[45][11] ,
         \ab[45][10] , \ab[44][44] , \ab[44][43] , \ab[44][42] , \ab[44][41] ,
         \ab[44][40] , \ab[44][39] , \ab[44][38] , \ab[44][37] , \ab[44][36] ,
         \ab[44][35] , \ab[44][34] , \ab[44][33] , \ab[44][32] , \ab[44][31] ,
         \ab[44][30] , \ab[44][29] , \ab[44][28] , \ab[44][27] , \ab[44][26] ,
         \ab[44][25] , \ab[44][24] , \ab[44][23] , \ab[44][22] , \ab[44][21] ,
         \ab[44][20] , \ab[44][19] , \ab[44][18] , \ab[44][17] , \ab[44][16] ,
         \ab[44][15] , \ab[44][14] , \ab[44][13] , \ab[44][12] , \ab[44][11] ,
         \ab[44][10] , \ab[43][43] , \ab[43][42] , \ab[43][41] , \ab[43][40] ,
         \ab[43][39] , \ab[43][38] , \ab[43][37] , \ab[43][36] , \ab[43][35] ,
         \ab[43][34] , \ab[43][33] , \ab[43][32] , \ab[43][31] , \ab[43][30] ,
         \ab[43][29] , \ab[43][28] , \ab[43][27] , \ab[43][26] , \ab[43][25] ,
         \ab[43][24] , \ab[43][23] , \ab[43][22] , \ab[43][21] , \ab[43][20] ,
         \ab[43][19] , \ab[43][18] , \ab[43][17] , \ab[43][16] , \ab[43][15] ,
         \ab[43][14] , \ab[43][13] , \ab[43][12] , \ab[43][11] , \ab[43][10] ,
         \ab[42][42] , \ab[42][41] , \ab[42][40] , \ab[42][39] , \ab[42][38] ,
         \ab[42][37] , \ab[42][36] , \ab[42][35] , \ab[42][34] , \ab[42][33] ,
         \ab[42][32] , \ab[42][31] , \ab[42][30] , \ab[42][29] , \ab[42][28] ,
         \ab[42][27] , \ab[42][26] , \ab[42][25] , \ab[42][24] , \ab[42][23] ,
         \ab[42][22] , \ab[42][21] , \ab[42][20] , \ab[42][19] , \ab[42][18] ,
         \ab[42][17] , \ab[42][16] , \ab[42][15] , \ab[42][14] , \ab[42][13] ,
         \ab[42][12] , \ab[42][11] , \ab[42][10] , \ab[41][41] , \ab[41][40] ,
         \ab[41][39] , \ab[41][38] , \ab[41][37] , \ab[41][36] , \ab[41][35] ,
         \ab[41][34] , \ab[41][33] , \ab[41][32] , \ab[41][31] , \ab[41][30] ,
         \ab[41][29] , \ab[41][28] , \ab[41][27] , \ab[41][26] , \ab[41][25] ,
         \ab[41][24] , \ab[41][23] , \ab[41][22] , \ab[41][21] , \ab[41][20] ,
         \ab[41][19] , \ab[41][18] , \ab[41][17] , \ab[41][16] , \ab[41][15] ,
         \ab[41][14] , \ab[41][13] , \ab[41][12] , \ab[41][11] , \ab[41][10] ,
         \ab[40][40] , \ab[40][39] , \ab[40][38] , \ab[40][37] , \ab[40][36] ,
         \ab[40][35] , \ab[40][34] , \ab[40][33] , \ab[40][32] , \ab[40][31] ,
         \ab[40][30] , \ab[40][29] , \ab[40][28] , \ab[40][27] , \ab[40][26] ,
         \ab[40][25] , \ab[40][24] , \ab[40][23] , \ab[40][22] , \ab[40][21] ,
         \ab[40][20] , \ab[40][19] , \ab[40][18] , \ab[40][17] , \ab[40][16] ,
         \ab[40][15] , \ab[40][14] , \ab[40][13] , \ab[40][12] , \ab[40][11] ,
         \ab[40][10] , \ab[39][39] , \ab[39][38] , \ab[39][37] , \ab[39][36] ,
         \ab[39][35] , \ab[39][34] , \ab[39][33] , \ab[39][32] , \ab[39][31] ,
         \ab[39][30] , \ab[39][29] , \ab[39][28] , \ab[39][27] , \ab[39][26] ,
         \ab[39][25] , \ab[39][24] , \ab[39][23] , \ab[39][22] , \ab[39][21] ,
         \ab[39][20] , \ab[39][19] , \ab[39][18] , \ab[39][17] , \ab[39][16] ,
         \ab[39][15] , \ab[39][14] , \ab[39][13] , \ab[39][12] , \ab[39][11] ,
         \ab[39][10] , \ab[38][38] , \ab[38][37] , \ab[38][36] , \ab[38][35] ,
         \ab[38][34] , \ab[38][33] , \ab[38][32] , \ab[38][31] , \ab[38][30] ,
         \ab[38][29] , \ab[38][28] , \ab[38][27] , \ab[38][26] , \ab[38][25] ,
         \ab[38][24] , \ab[38][23] , \ab[38][22] , \ab[38][21] , \ab[38][20] ,
         \ab[38][19] , \ab[38][18] , \ab[38][17] , \ab[38][16] , \ab[38][15] ,
         \ab[38][14] , \ab[38][13] , \ab[38][12] , \ab[38][11] , \ab[38][10] ,
         \ab[37][37] , \ab[37][36] , \ab[37][35] , \ab[37][34] , \ab[37][33] ,
         \ab[37][32] , \ab[37][31] , \ab[37][30] , \ab[37][29] , \ab[37][28] ,
         \ab[37][27] , \ab[37][26] , \ab[37][25] , \ab[37][24] , \ab[37][23] ,
         \ab[37][22] , \ab[37][21] , \ab[37][20] , \ab[37][19] , \ab[37][18] ,
         \ab[37][17] , \ab[37][16] , \ab[37][15] , \ab[37][14] , \ab[37][13] ,
         \ab[37][12] , \ab[37][11] , \ab[36][36] , \ab[36][35] , \ab[36][34] ,
         \ab[36][33] , \ab[36][32] , \ab[36][31] , \ab[36][30] , \ab[36][29] ,
         \ab[36][28] , \ab[36][27] , \ab[36][26] , \ab[36][25] , \ab[36][24] ,
         \ab[36][23] , \ab[36][22] , \ab[36][21] , \ab[36][20] , \ab[36][19] ,
         \ab[36][18] , \ab[36][17] , \ab[36][16] , \ab[36][15] , \ab[36][14] ,
         \ab[36][13] , \ab[36][12] , \ab[36][11] , \ab[35][35] , \ab[35][34] ,
         \ab[35][33] , \ab[35][32] , \ab[35][31] , \ab[35][30] , \ab[35][29] ,
         \ab[35][28] , \ab[35][27] , \ab[35][26] , \ab[35][25] , \ab[35][24] ,
         \ab[35][23] , \ab[35][22] , \ab[35][21] , \ab[35][20] , \ab[35][19] ,
         \ab[35][18] , \ab[35][17] , \ab[35][16] , \ab[35][15] , \ab[35][14] ,
         \ab[35][13] , \ab[35][12] , \ab[35][11] , \ab[34][34] , \ab[34][33] ,
         \ab[34][32] , \ab[34][31] , \ab[34][30] , \ab[34][29] , \ab[34][28] ,
         \ab[34][27] , \ab[34][26] , \ab[34][25] , \ab[34][24] , \ab[34][23] ,
         \ab[34][22] , \ab[34][21] , \ab[34][20] , \ab[34][19] , \ab[34][18] ,
         \ab[34][17] , \ab[34][16] , \ab[34][15] , \ab[34][14] , \ab[34][13] ,
         \ab[34][12] , \ab[33][33] , \ab[33][32] , \ab[33][31] , \ab[33][30] ,
         \ab[33][29] , \ab[33][28] , \ab[33][27] , \ab[33][26] , \ab[33][25] ,
         \ab[33][24] , \ab[33][23] , \ab[33][22] , \ab[33][21] , \ab[33][20] ,
         \ab[33][19] , \ab[33][18] , \ab[33][17] , \ab[33][16] , \ab[33][15] ,
         \ab[33][14] , \ab[33][13] , \ab[33][12] , \ab[32][32] , \ab[32][31] ,
         \ab[32][30] , \ab[32][29] , \ab[32][28] , \ab[32][27] , \ab[32][26] ,
         \ab[32][25] , \ab[32][24] , \ab[32][23] , \ab[32][22] , \ab[32][21] ,
         \ab[32][20] , \ab[32][19] , \ab[32][18] , \ab[32][17] , \ab[32][16] ,
         \ab[32][15] , \ab[32][14] , \ab[32][13] , \ab[31][31] , \ab[31][30] ,
         \ab[31][29] , \ab[31][28] , \ab[31][27] , \ab[31][26] , \ab[31][25] ,
         \ab[31][24] , \ab[31][23] , \ab[31][22] , \ab[31][21] , \ab[31][20] ,
         \ab[31][19] , \ab[31][18] , \ab[31][17] , \ab[31][16] , \ab[31][15] ,
         \ab[31][14] , \ab[31][13] , \ab[30][30] , \ab[30][29] , \ab[30][28] ,
         \ab[30][27] , \ab[30][26] , \ab[30][25] , \ab[30][24] , \ab[30][23] ,
         \ab[30][22] , \ab[30][21] , \ab[30][20] , \ab[30][19] , \ab[30][18] ,
         \ab[30][17] , \ab[30][16] , \ab[30][15] , \ab[30][14] , \ab[29][29] ,
         \ab[29][28] , \ab[29][27] , \ab[29][26] , \ab[29][25] , \ab[29][24] ,
         \ab[29][23] , \ab[29][22] , \ab[29][21] , \ab[29][20] , \ab[29][19] ,
         \ab[29][18] , \ab[29][17] , \ab[29][16] , \ab[29][15] , \ab[29][14] ,
         \ab[28][28] , \ab[28][27] , \ab[28][26] , \ab[28][25] , \ab[28][24] ,
         \ab[28][23] , \ab[28][22] , \ab[28][21] , \ab[28][20] , \ab[28][19] ,
         \ab[28][18] , \ab[28][17] , \ab[28][16] , \ab[28][15] , \ab[28][14] ,
         \ab[27][27] , \ab[27][26] , \ab[27][25] , \ab[27][24] , \ab[27][23] ,
         \ab[27][22] , \ab[27][21] , \ab[27][20] , \ab[27][19] , \ab[27][18] ,
         \ab[27][17] , \ab[27][16] , \ab[27][15] , \ab[27][14] , \ab[26][26] ,
         \ab[26][25] , \ab[26][24] , \ab[26][23] , \ab[26][22] , \ab[26][21] ,
         \ab[26][20] , \ab[26][19] , \ab[26][18] , \ab[26][17] , \ab[26][16] ,
         \ab[26][15] , \ab[25][25] , \ab[25][24] , \ab[25][23] , \ab[25][22] ,
         \ab[25][21] , \ab[25][20] , \ab[25][19] , \ab[25][18] , \ab[25][17] ,
         \ab[25][16] , \ab[25][15] , \ab[24][24] , \ab[24][23] , \ab[24][22] ,
         \ab[24][21] , \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] ,
         \ab[24][16] , \ab[24][15] , \ab[23][23] , \ab[23][22] , \ab[23][21] ,
         \ab[23][20] , \ab[23][19] , \ab[23][18] , \ab[23][17] , \ab[23][16] ,
         \ab[23][15] , \ab[22][22] , \ab[22][21] , \ab[22][20] , \ab[22][19] ,
         \ab[22][18] , \ab[22][17] , \ab[22][16] , \ab[22][15] , \ab[21][21] ,
         \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] , \ab[21][16] ,
         \ab[21][15] , \ab[20][20] , \ab[20][19] , \ab[20][18] , \ab[20][17] ,
         \ab[20][16] , \ab[20][15] , \ab[19][19] , \ab[19][18] , \ab[19][17] ,
         \ab[19][16] , \ab[19][15] , \ab[18][18] , \ab[18][17] , \ab[18][16] ,
         \ab[18][15] , \ab[17][17] , \ab[17][16] , \ab[17][15] , \ab[16][16] ,
         \ab[16][15] , \ab[15][15] , \ab[14][14] , \ab[13][13] , \ab[12][12] ,
         \ab[11][11] , \ab[10][10] , \ab[9][47] , \ab[9][46] , \ab[9][45] ,
         \ab[9][44] , \ab[9][43] , \ab[9][42] , \ab[9][41] , \ab[9][40] ,
         \ab[9][9] , \ab[8][47] , \ab[8][46] , \ab[8][45] , \ab[8][44] ,
         \ab[8][8] , \ab[7][47] , \ab[7][46] , \ab[7][7] , \ab[6][47] ,
         \ab[6][6] , \ab[5][5] , \ab[4][4] , \ab[3][3] , \ab[2][2] ,
         \ab[1][1] , \ab[1][0] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][46] , \CARRYB[4][45] ,
         \CARRYB[4][44] , \CARRYB[4][43] , \CARRYB[4][42] , \CARRYB[4][41] ,
         \CARRYB[4][40] , \CARRYB[4][39] , \CARRYB[4][38] , \CARRYB[4][37] ,
         \CARRYB[4][36] , \CARRYB[4][35] , \CARRYB[4][34] , \CARRYB[4][33] ,
         \CARRYB[4][32] , \CARRYB[4][31] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][46] , \CARRYB[3][45] , \CARRYB[3][44] ,
         \CARRYB[3][43] , \CARRYB[3][42] , \CARRYB[3][41] , \CARRYB[3][40] ,
         \CARRYB[3][39] , \CARRYB[3][38] , \CARRYB[3][37] , \CARRYB[3][36] ,
         \CARRYB[3][35] , \CARRYB[3][34] , \CARRYB[3][33] , \CARRYB[3][32] ,
         \CARRYB[3][31] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][46] , \CARRYB[2][45] , \CARRYB[2][44] , \CARRYB[2][43] ,
         \CARRYB[2][42] , \CARRYB[2][41] , \CARRYB[2][40] , \CARRYB[2][39] ,
         \CARRYB[2][38] , \CARRYB[2][37] , \CARRYB[2][36] , \CARRYB[2][35] ,
         \CARRYB[2][34] , \CARRYB[2][33] , \CARRYB[2][32] , \CARRYB[2][31] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][46] ,
         \CARRYB[1][45] , \CARRYB[1][44] , \CARRYB[1][43] , \CARRYB[1][42] ,
         \CARRYB[1][41] , \CARRYB[1][40] , \CARRYB[1][39] , \CARRYB[1][38] ,
         \CARRYB[1][37] , \CARRYB[1][36] , \CARRYB[1][35] , \CARRYB[1][34] ,
         \CARRYB[1][33] , \CARRYB[1][32] , \CARRYB[1][31] , \CARRYB[1][30] ,
         \CARRYB[1][29] , \CARRYB[1][28] , \CARRYB[1][27] , \CARRYB[1][26] ,
         \CARRYB[1][25] , \CARRYB[1][23] , \CARRYB[1][22] , \CARRYB[1][21] ,
         \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] , \CARRYB[1][17] ,
         \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][46] , \SUMB[4][45] ,
         \SUMB[4][44] , \SUMB[4][43] , \SUMB[4][42] , \SUMB[4][41] ,
         \SUMB[4][40] , \SUMB[4][39] , \SUMB[4][38] , \SUMB[4][37] ,
         \SUMB[4][36] , \SUMB[4][35] , \SUMB[4][34] , \SUMB[4][33] ,
         \SUMB[4][32] , \SUMB[4][31] , \SUMB[4][30] , \SUMB[4][29] ,
         \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] , \SUMB[4][25] ,
         \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] , \SUMB[4][21] ,
         \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] , \SUMB[4][17] ,
         \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] ,
         \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] ,
         \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][46] ,
         \SUMB[3][45] , \SUMB[3][44] , \SUMB[3][43] , \SUMB[3][42] ,
         \SUMB[3][41] , \SUMB[3][40] , \SUMB[3][39] , \SUMB[3][38] ,
         \SUMB[3][37] , \SUMB[3][36] , \SUMB[3][35] , \SUMB[3][34] ,
         \SUMB[3][33] , \SUMB[3][32] , \SUMB[3][31] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][46] ,
         \SUMB[2][45] , \SUMB[2][44] , \SUMB[2][43] , \SUMB[2][42] ,
         \SUMB[2][41] , \SUMB[2][40] , \SUMB[2][39] , \SUMB[2][38] ,
         \SUMB[2][37] , \SUMB[2][36] , \SUMB[2][35] , \SUMB[2][34] ,
         \SUMB[2][33] , \SUMB[2][32] , \SUMB[2][31] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][46] ,
         \SUMB[1][45] , \SUMB[1][44] , \SUMB[1][43] , \SUMB[1][42] ,
         \SUMB[1][41] , \SUMB[1][40] , \SUMB[1][39] , \SUMB[1][38] ,
         \SUMB[1][37] , \SUMB[1][36] , \SUMB[1][35] , \SUMB[1][34] ,
         \SUMB[1][33] , \SUMB[1][32] , \SUMB[1][31] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[15][46] , \CARRYB[15][45] , \CARRYB[15][44] ,
         \CARRYB[15][43] , \CARRYB[15][42] , \CARRYB[15][41] ,
         \CARRYB[15][40] , \CARRYB[15][39] , \CARRYB[15][38] ,
         \CARRYB[15][37] , \CARRYB[15][36] , \CARRYB[15][35] ,
         \CARRYB[15][34] , \CARRYB[15][33] , \CARRYB[15][32] ,
         \CARRYB[15][31] , \CARRYB[15][30] , \CARRYB[15][29] ,
         \CARRYB[15][28] , \CARRYB[15][27] , \CARRYB[15][26] ,
         \CARRYB[15][25] , \CARRYB[15][24] , \CARRYB[15][23] ,
         \CARRYB[15][22] , \CARRYB[15][21] , \CARRYB[15][20] ,
         \CARRYB[15][19] , \CARRYB[15][18] , \CARRYB[15][17] ,
         \CARRYB[15][16] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][46] ,
         \CARRYB[14][45] , \CARRYB[14][44] , \CARRYB[14][43] ,
         \CARRYB[14][42] , \CARRYB[14][41] , \CARRYB[14][40] ,
         \CARRYB[14][39] , \CARRYB[14][38] , \CARRYB[14][37] ,
         \CARRYB[14][36] , \CARRYB[14][35] , \CARRYB[14][34] ,
         \CARRYB[14][33] , \CARRYB[14][32] , \CARRYB[14][31] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][46] , \CARRYB[13][45] , \CARRYB[13][44] ,
         \CARRYB[13][43] , \CARRYB[13][42] , \CARRYB[13][41] ,
         \CARRYB[13][40] , \CARRYB[13][39] , \CARRYB[13][38] ,
         \CARRYB[13][37] , \CARRYB[13][36] , \CARRYB[13][35] ,
         \CARRYB[13][34] , \CARRYB[13][33] , \CARRYB[13][32] ,
         \CARRYB[13][31] , \CARRYB[13][30] , \CARRYB[13][29] ,
         \CARRYB[13][28] , \CARRYB[13][27] , \CARRYB[13][26] ,
         \CARRYB[13][25] , \CARRYB[13][24] , \CARRYB[13][23] ,
         \CARRYB[13][22] , \CARRYB[13][21] , \CARRYB[13][20] ,
         \CARRYB[13][19] , \CARRYB[13][18] , \CARRYB[13][17] ,
         \CARRYB[13][16] , \CARRYB[13][15] , \CARRYB[13][14] ,
         \CARRYB[13][13] , \CARRYB[13][12] , \CARRYB[13][11] ,
         \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] , \CARRYB[13][7] ,
         \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] , \CARRYB[13][3] ,
         \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] , \CARRYB[12][46] ,
         \CARRYB[12][45] , \CARRYB[12][44] , \CARRYB[12][43] ,
         \CARRYB[12][42] , \CARRYB[12][41] , \CARRYB[12][40] ,
         \CARRYB[12][39] , \CARRYB[12][38] , \CARRYB[12][37] ,
         \CARRYB[12][36] , \CARRYB[12][35] , \CARRYB[12][34] ,
         \CARRYB[12][33] , \CARRYB[12][32] , \CARRYB[12][31] ,
         \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][46] , \CARRYB[11][45] , \CARRYB[11][44] ,
         \CARRYB[11][43] , \CARRYB[11][42] , \CARRYB[11][41] ,
         \CARRYB[11][40] , \CARRYB[11][39] , \CARRYB[11][38] ,
         \CARRYB[11][37] , \CARRYB[11][36] , \CARRYB[11][35] ,
         \CARRYB[11][34] , \CARRYB[11][33] , \CARRYB[11][32] ,
         \CARRYB[11][31] , \CARRYB[11][30] , \CARRYB[11][29] ,
         \CARRYB[11][28] , \CARRYB[11][27] , \CARRYB[11][26] ,
         \CARRYB[11][25] , \CARRYB[11][24] , \CARRYB[11][23] ,
         \CARRYB[11][22] , \CARRYB[11][21] , \CARRYB[11][20] ,
         \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \CARRYB[11][15] , \CARRYB[11][14] ,
         \CARRYB[11][13] , \CARRYB[11][12] , \CARRYB[11][11] ,
         \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] , \CARRYB[11][7] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][46] ,
         \CARRYB[10][45] , \CARRYB[10][44] , \CARRYB[10][43] ,
         \CARRYB[10][42] , \CARRYB[10][41] , \CARRYB[10][40] ,
         \CARRYB[10][39] , \CARRYB[10][38] , \CARRYB[10][37] ,
         \CARRYB[10][36] , \CARRYB[10][35] , \CARRYB[10][34] ,
         \CARRYB[10][33] , \CARRYB[10][32] , \CARRYB[10][31] ,
         \CARRYB[10][30] , \CARRYB[10][29] , \CARRYB[10][28] ,
         \CARRYB[10][27] , \CARRYB[10][26] , \CARRYB[10][25] ,
         \CARRYB[10][24] , \CARRYB[10][23] , \CARRYB[10][22] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][46] , \CARRYB[9][45] , \CARRYB[9][44] ,
         \CARRYB[9][43] , \CARRYB[9][42] , \CARRYB[9][41] , \CARRYB[9][40] ,
         \CARRYB[9][39] , \CARRYB[9][38] , \CARRYB[9][37] , \CARRYB[9][36] ,
         \CARRYB[9][35] , \CARRYB[9][34] , \CARRYB[9][33] , \CARRYB[9][32] ,
         \CARRYB[9][31] , \CARRYB[9][30] , \CARRYB[9][29] , \CARRYB[9][28] ,
         \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][25] , \CARRYB[9][24] ,
         \CARRYB[9][23] , \CARRYB[9][22] , \CARRYB[9][21] , \CARRYB[9][20] ,
         \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] , \CARRYB[9][16] ,
         \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] ,
         \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] ,
         \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] ,
         \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] ,
         \CARRYB[8][46] , \CARRYB[8][45] , \CARRYB[8][44] , \CARRYB[8][43] ,
         \CARRYB[8][42] , \CARRYB[8][41] , \CARRYB[8][40] , \CARRYB[8][39] ,
         \CARRYB[8][38] , \CARRYB[8][37] , \CARRYB[8][36] , \CARRYB[8][35] ,
         \CARRYB[8][34] , \CARRYB[8][33] , \CARRYB[8][32] , \CARRYB[8][31] ,
         \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] , \CARRYB[8][27] ,
         \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] , \CARRYB[8][23] ,
         \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] , \CARRYB[8][19] ,
         \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] ,
         \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] ,
         \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] ,
         \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][46] ,
         \CARRYB[7][45] , \CARRYB[7][44] , \CARRYB[7][43] , \CARRYB[7][42] ,
         \CARRYB[7][41] , \CARRYB[7][40] , \CARRYB[7][39] , \CARRYB[7][38] ,
         \CARRYB[7][37] , \CARRYB[7][36] , \CARRYB[7][35] , \CARRYB[7][34] ,
         \CARRYB[7][33] , \CARRYB[7][32] , \CARRYB[7][31] , \CARRYB[7][30] ,
         \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] ,
         \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] ,
         \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] ,
         \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][46] , \CARRYB[6][45] ,
         \CARRYB[6][44] , \CARRYB[6][43] , \CARRYB[6][42] , \CARRYB[6][41] ,
         \CARRYB[6][40] , \CARRYB[6][39] , \CARRYB[6][38] , \CARRYB[6][37] ,
         \CARRYB[6][36] , \CARRYB[6][35] , \CARRYB[6][34] , \CARRYB[6][33] ,
         \CARRYB[6][32] , \CARRYB[6][31] , \CARRYB[6][30] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][46] , \CARRYB[5][45] , \CARRYB[5][44] ,
         \CARRYB[5][43] , \CARRYB[5][42] , \CARRYB[5][41] , \CARRYB[5][40] ,
         \CARRYB[5][39] , \CARRYB[5][38] , \CARRYB[5][37] , \CARRYB[5][36] ,
         \CARRYB[5][35] , \CARRYB[5][34] , \CARRYB[5][33] , \CARRYB[5][32] ,
         \CARRYB[5][31] , \CARRYB[5][30] , \CARRYB[5][29] , \CARRYB[5][28] ,
         \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] , \CARRYB[5][24] ,
         \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] , \CARRYB[5][20] ,
         \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] , \CARRYB[5][16] ,
         \SUMB[15][46] , \SUMB[15][45] , \SUMB[15][44] , \SUMB[15][43] ,
         \SUMB[15][42] , \SUMB[15][41] , \SUMB[15][40] , \SUMB[15][39] ,
         \SUMB[15][38] , \SUMB[15][37] , \SUMB[15][36] , \SUMB[15][35] ,
         \SUMB[15][34] , \SUMB[15][33] , \SUMB[15][32] , \SUMB[15][31] ,
         \SUMB[15][30] , \SUMB[15][29] , \SUMB[15][28] , \SUMB[15][27] ,
         \SUMB[15][26] , \SUMB[15][25] , \SUMB[15][24] , \SUMB[15][23] ,
         \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] , \SUMB[15][19] ,
         \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] , \SUMB[15][15] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][46] , \SUMB[14][45] ,
         \SUMB[14][44] , \SUMB[14][43] , \SUMB[14][42] , \SUMB[14][41] ,
         \SUMB[14][40] , \SUMB[14][39] , \SUMB[14][38] , \SUMB[14][37] ,
         \SUMB[14][36] , \SUMB[14][35] , \SUMB[14][34] , \SUMB[14][33] ,
         \SUMB[14][32] , \SUMB[14][31] , \SUMB[14][30] , \SUMB[14][29] ,
         \SUMB[14][28] , \SUMB[14][27] , \SUMB[14][26] , \SUMB[14][25] ,
         \SUMB[14][24] , \SUMB[14][23] , \SUMB[14][22] , \SUMB[14][21] ,
         \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] , \SUMB[14][17] ,
         \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][46] , \SUMB[13][45] , \SUMB[13][44] , \SUMB[13][43] ,
         \SUMB[13][42] , \SUMB[13][41] , \SUMB[13][40] , \SUMB[13][39] ,
         \SUMB[13][38] , \SUMB[13][37] , \SUMB[13][36] , \SUMB[13][35] ,
         \SUMB[13][34] , \SUMB[13][33] , \SUMB[13][32] , \SUMB[13][31] ,
         \SUMB[13][30] , \SUMB[13][29] , \SUMB[13][28] , \SUMB[13][27] ,
         \SUMB[13][26] , \SUMB[13][25] , \SUMB[13][24] , \SUMB[13][23] ,
         \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] , \SUMB[13][19] ,
         \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] , \SUMB[13][15] ,
         \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] ,
         \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][46] , \SUMB[12][45] ,
         \SUMB[12][44] , \SUMB[12][43] , \SUMB[12][42] , \SUMB[12][41] ,
         \SUMB[12][40] , \SUMB[12][39] , \SUMB[12][38] , \SUMB[12][37] ,
         \SUMB[12][36] , \SUMB[12][35] , \SUMB[12][34] , \SUMB[12][33] ,
         \SUMB[12][32] , \SUMB[12][31] , \SUMB[12][30] , \SUMB[12][29] ,
         \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] , \SUMB[12][25] ,
         \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] , \SUMB[12][21] ,
         \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] , \SUMB[12][17] ,
         \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] ,
         \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] ,
         \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][46] , \SUMB[11][45] , \SUMB[11][44] , \SUMB[11][43] ,
         \SUMB[11][42] , \SUMB[11][41] , \SUMB[11][40] , \SUMB[11][39] ,
         \SUMB[11][38] , \SUMB[11][37] , \SUMB[11][36] , \SUMB[11][35] ,
         \SUMB[11][34] , \SUMB[11][33] , \SUMB[11][32] , \SUMB[11][31] ,
         \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] , \SUMB[11][27] ,
         \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] , \SUMB[11][23] ,
         \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] , \SUMB[11][19] ,
         \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][46] , \SUMB[10][45] ,
         \SUMB[10][44] , \SUMB[10][43] , \SUMB[10][42] , \SUMB[10][41] ,
         \SUMB[10][40] , \SUMB[10][39] , \SUMB[10][38] , \SUMB[10][37] ,
         \SUMB[10][36] , \SUMB[10][35] , \SUMB[10][34] , \SUMB[10][33] ,
         \SUMB[10][32] , \SUMB[10][31] , \SUMB[10][30] , \SUMB[10][29] ,
         \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] , \SUMB[10][25] ,
         \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] , \SUMB[10][21] ,
         \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] ,
         \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][46] , \SUMB[9][45] , \SUMB[9][44] , \SUMB[9][43] ,
         \SUMB[9][42] , \SUMB[9][41] , \SUMB[9][40] , \SUMB[9][39] ,
         \SUMB[9][38] , \SUMB[9][37] , \SUMB[9][36] , \SUMB[9][35] ,
         \SUMB[9][34] , \SUMB[9][33] , \SUMB[9][32] , \SUMB[9][31] ,
         \SUMB[9][30] , \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] ,
         \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] ,
         \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] ,
         \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] ,
         \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] ,
         \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][46] , \SUMB[8][45] , \SUMB[8][44] , \SUMB[8][43] ,
         \SUMB[8][42] , \SUMB[8][41] , \SUMB[8][40] , \SUMB[8][39] ,
         \SUMB[8][38] , \SUMB[8][37] , \SUMB[8][36] , \SUMB[8][35] ,
         \SUMB[8][34] , \SUMB[8][33] , \SUMB[8][32] , \SUMB[8][31] ,
         \SUMB[8][30] , \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] ,
         \SUMB[8][26] , \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] ,
         \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][46] , \SUMB[7][45] , \SUMB[7][44] , \SUMB[7][43] ,
         \SUMB[7][42] , \SUMB[7][41] , \SUMB[7][40] , \SUMB[7][39] ,
         \SUMB[7][38] , \SUMB[7][37] , \SUMB[7][36] , \SUMB[7][35] ,
         \SUMB[7][34] , \SUMB[7][33] , \SUMB[7][32] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][46] , \SUMB[6][45] , \SUMB[6][44] , \SUMB[6][43] ,
         \SUMB[6][42] , \SUMB[6][41] , \SUMB[6][40] , \SUMB[6][39] ,
         \SUMB[6][38] , \SUMB[6][37] , \SUMB[6][36] , \SUMB[6][35] ,
         \SUMB[6][34] , \SUMB[6][33] , \SUMB[6][32] , \SUMB[6][31] ,
         \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] ,
         \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] ,
         \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] ,
         \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][46] , \SUMB[5][45] , \SUMB[5][44] , \SUMB[5][43] ,
         \SUMB[5][42] , \SUMB[5][41] , \SUMB[5][40] , \SUMB[5][39] ,
         \SUMB[5][38] , \SUMB[5][37] , \SUMB[5][36] , \SUMB[5][35] ,
         \SUMB[5][34] , \SUMB[5][33] , \SUMB[5][32] , \SUMB[5][31] ,
         \SUMB[5][30] , \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] ,
         \SUMB[5][26] , \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] ,
         \SUMB[5][22] , \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] ,
         \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] , \CARRYB[26][31] ,
         \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][46] , \CARRYB[25][45] , \CARRYB[25][44] ,
         \CARRYB[25][43] , \CARRYB[25][42] , \CARRYB[25][41] ,
         \CARRYB[25][40] , \CARRYB[25][39] , \CARRYB[25][38] ,
         \CARRYB[25][37] , \CARRYB[25][36] , \CARRYB[25][35] ,
         \CARRYB[25][34] , \CARRYB[25][33] , \CARRYB[25][32] ,
         \CARRYB[25][31] , \CARRYB[25][30] , \CARRYB[25][29] ,
         \CARRYB[25][28] , \CARRYB[25][27] , \CARRYB[25][26] ,
         \CARRYB[25][25] , \CARRYB[25][24] , \CARRYB[25][23] ,
         \CARRYB[25][22] , \CARRYB[25][21] , \CARRYB[25][20] ,
         \CARRYB[25][19] , \CARRYB[25][18] , \CARRYB[25][17] ,
         \CARRYB[25][16] , \CARRYB[25][15] , \CARRYB[25][14] ,
         \CARRYB[25][13] , \CARRYB[25][12] , \CARRYB[25][11] ,
         \CARRYB[25][10] , \CARRYB[25][9] , \CARRYB[25][8] , \CARRYB[25][7] ,
         \CARRYB[25][6] , \CARRYB[25][5] , \CARRYB[25][4] , \CARRYB[25][3] ,
         \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] , \CARRYB[24][46] ,
         \CARRYB[24][45] , \CARRYB[24][44] , \CARRYB[24][43] ,
         \CARRYB[24][42] , \CARRYB[24][41] , \CARRYB[24][40] ,
         \CARRYB[24][39] , \CARRYB[24][38] , \CARRYB[24][37] ,
         \CARRYB[24][36] , \CARRYB[24][35] , \CARRYB[24][34] ,
         \CARRYB[24][33] , \CARRYB[24][32] , \CARRYB[24][31] ,
         \CARRYB[24][30] , \CARRYB[24][29] , \CARRYB[24][28] ,
         \CARRYB[24][27] , \CARRYB[24][26] , \CARRYB[24][25] ,
         \CARRYB[24][24] , \CARRYB[24][23] , \CARRYB[24][22] ,
         \CARRYB[24][21] , \CARRYB[24][20] , \CARRYB[24][19] ,
         \CARRYB[24][18] , \CARRYB[24][17] , \CARRYB[24][16] ,
         \CARRYB[24][15] , \CARRYB[24][14] , \CARRYB[24][13] ,
         \CARRYB[24][12] , \CARRYB[24][11] , \CARRYB[24][10] , \CARRYB[24][9] ,
         \CARRYB[24][8] , \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] ,
         \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] ,
         \CARRYB[24][0] , \CARRYB[23][46] , \CARRYB[23][45] , \CARRYB[23][44] ,
         \CARRYB[23][43] , \CARRYB[23][42] , \CARRYB[23][41] ,
         \CARRYB[23][40] , \CARRYB[23][39] , \CARRYB[23][38] ,
         \CARRYB[23][37] , \CARRYB[23][36] , \CARRYB[23][35] ,
         \CARRYB[23][34] , \CARRYB[23][33] , \CARRYB[23][32] ,
         \CARRYB[23][31] , \CARRYB[23][30] , \CARRYB[23][29] ,
         \CARRYB[23][28] , \CARRYB[23][27] , \CARRYB[23][26] ,
         \CARRYB[23][25] , \CARRYB[23][24] , \CARRYB[23][23] ,
         \CARRYB[23][22] , \CARRYB[23][21] , \CARRYB[23][20] ,
         \CARRYB[23][19] , \CARRYB[23][18] , \CARRYB[23][17] ,
         \CARRYB[23][16] , \CARRYB[23][15] , \CARRYB[23][14] ,
         \CARRYB[23][13] , \CARRYB[23][12] , \CARRYB[23][11] ,
         \CARRYB[23][10] , \CARRYB[23][9] , \CARRYB[23][8] , \CARRYB[23][7] ,
         \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] ,
         \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][46] ,
         \CARRYB[22][45] , \CARRYB[22][44] , \CARRYB[22][43] ,
         \CARRYB[22][42] , \CARRYB[22][41] , \CARRYB[22][40] ,
         \CARRYB[22][39] , \CARRYB[22][38] , \CARRYB[22][37] ,
         \CARRYB[22][36] , \CARRYB[22][35] , \CARRYB[22][34] ,
         \CARRYB[22][33] , \CARRYB[22][32] , \CARRYB[22][31] ,
         \CARRYB[22][30] , \CARRYB[22][29] , \CARRYB[22][28] ,
         \CARRYB[22][27] , \CARRYB[22][26] , \CARRYB[22][25] ,
         \CARRYB[22][24] , \CARRYB[22][23] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][12] , \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] ,
         \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][46] , \CARRYB[21][45] , \CARRYB[21][44] ,
         \CARRYB[21][43] , \CARRYB[21][42] , \CARRYB[21][41] ,
         \CARRYB[21][40] , \CARRYB[21][39] , \CARRYB[21][38] ,
         \CARRYB[21][37] , \CARRYB[21][36] , \CARRYB[21][35] ,
         \CARRYB[21][34] , \CARRYB[21][33] , \CARRYB[21][32] ,
         \CARRYB[21][31] , \CARRYB[21][30] , \CARRYB[21][29] ,
         \CARRYB[21][28] , \CARRYB[21][27] , \CARRYB[21][26] ,
         \CARRYB[21][25] , \CARRYB[21][24] , \CARRYB[21][23] ,
         \CARRYB[21][22] , \CARRYB[21][21] , \CARRYB[21][20] ,
         \CARRYB[21][19] , \CARRYB[21][18] , \CARRYB[21][17] ,
         \CARRYB[21][16] , \CARRYB[21][15] , \CARRYB[21][14] ,
         \CARRYB[21][13] , \CARRYB[21][12] , \CARRYB[21][11] ,
         \CARRYB[21][10] , \CARRYB[21][9] , \CARRYB[21][8] , \CARRYB[21][7] ,
         \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] , \CARRYB[21][3] ,
         \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] , \CARRYB[20][46] ,
         \CARRYB[20][45] , \CARRYB[20][44] , \CARRYB[20][43] ,
         \CARRYB[20][42] , \CARRYB[20][41] , \CARRYB[20][40] ,
         \CARRYB[20][39] , \CARRYB[20][38] , \CARRYB[20][37] ,
         \CARRYB[20][36] , \CARRYB[20][35] , \CARRYB[20][34] ,
         \CARRYB[20][33] , \CARRYB[20][32] , \CARRYB[20][31] ,
         \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][46] , \CARRYB[19][45] , \CARRYB[19][44] ,
         \CARRYB[19][43] , \CARRYB[19][42] , \CARRYB[19][41] ,
         \CARRYB[19][40] , \CARRYB[19][39] , \CARRYB[19][38] ,
         \CARRYB[19][37] , \CARRYB[19][36] , \CARRYB[19][35] ,
         \CARRYB[19][34] , \CARRYB[19][33] , \CARRYB[19][32] ,
         \CARRYB[19][31] , \CARRYB[19][30] , \CARRYB[19][29] ,
         \CARRYB[19][28] , \CARRYB[19][27] , \CARRYB[19][26] ,
         \CARRYB[19][25] , \CARRYB[19][24] , \CARRYB[19][23] ,
         \CARRYB[19][22] , \CARRYB[19][21] , \CARRYB[19][20] ,
         \CARRYB[19][19] , \CARRYB[19][18] , \CARRYB[19][17] ,
         \CARRYB[19][16] , \CARRYB[19][15] , \CARRYB[19][14] ,
         \CARRYB[19][13] , \CARRYB[19][12] , \CARRYB[19][11] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][46] ,
         \CARRYB[18][45] , \CARRYB[18][44] , \CARRYB[18][43] ,
         \CARRYB[18][42] , \CARRYB[18][41] , \CARRYB[18][40] ,
         \CARRYB[18][39] , \CARRYB[18][38] , \CARRYB[18][37] ,
         \CARRYB[18][36] , \CARRYB[18][35] , \CARRYB[18][34] ,
         \CARRYB[18][33] , \CARRYB[18][32] , \CARRYB[18][31] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][46] , \CARRYB[17][45] , \CARRYB[17][44] ,
         \CARRYB[17][43] , \CARRYB[17][42] , \CARRYB[17][41] ,
         \CARRYB[17][40] , \CARRYB[17][39] , \CARRYB[17][38] ,
         \CARRYB[17][37] , \CARRYB[17][36] , \CARRYB[17][35] ,
         \CARRYB[17][34] , \CARRYB[17][33] , \CARRYB[17][32] ,
         \CARRYB[17][31] , \CARRYB[17][30] , \CARRYB[17][29] ,
         \CARRYB[17][28] , \CARRYB[17][27] , \CARRYB[17][26] ,
         \CARRYB[17][25] , \CARRYB[17][24] , \CARRYB[17][23] ,
         \CARRYB[17][22] , \CARRYB[17][21] , \CARRYB[17][20] ,
         \CARRYB[17][19] , \CARRYB[17][18] , \CARRYB[17][17] ,
         \CARRYB[17][16] , \CARRYB[17][15] , \CARRYB[17][14] ,
         \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][46] ,
         \CARRYB[16][45] , \CARRYB[16][44] , \CARRYB[16][43] ,
         \CARRYB[16][42] , \CARRYB[16][41] , \CARRYB[16][40] ,
         \CARRYB[16][39] , \CARRYB[16][38] , \CARRYB[16][37] ,
         \CARRYB[16][36] , \CARRYB[16][35] , \CARRYB[16][34] ,
         \CARRYB[16][33] , \CARRYB[16][32] , \CARRYB[16][31] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \SUMB[26][31] , \SUMB[26][30] , \SUMB[26][29] ,
         \SUMB[26][28] , \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] ,
         \SUMB[26][24] , \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] ,
         \SUMB[26][20] , \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] ,
         \SUMB[26][16] , \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] ,
         \SUMB[26][12] , \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] ,
         \SUMB[26][8] , \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] ,
         \SUMB[26][4] , \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] ,
         \SUMB[25][46] , \SUMB[25][45] , \SUMB[25][44] , \SUMB[25][43] ,
         \SUMB[25][42] , \SUMB[25][41] , \SUMB[25][40] , \SUMB[25][39] ,
         \SUMB[25][38] , \SUMB[25][37] , \SUMB[25][36] , \SUMB[25][35] ,
         \SUMB[25][34] , \SUMB[25][33] , \SUMB[25][32] , \SUMB[25][31] ,
         \SUMB[25][30] , \SUMB[25][29] , \SUMB[25][28] , \SUMB[25][27] ,
         \SUMB[25][26] , \SUMB[25][25] , \SUMB[25][24] , \SUMB[25][23] ,
         \SUMB[25][22] , \SUMB[25][21] , \SUMB[25][20] , \SUMB[25][19] ,
         \SUMB[25][18] , \SUMB[25][17] , \SUMB[25][16] , \SUMB[25][15] ,
         \SUMB[25][14] , \SUMB[25][13] , \SUMB[25][12] , \SUMB[25][11] ,
         \SUMB[25][10] , \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] ,
         \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] ,
         \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][46] , \SUMB[24][45] ,
         \SUMB[24][44] , \SUMB[24][43] , \SUMB[24][42] , \SUMB[24][41] ,
         \SUMB[24][40] , \SUMB[24][39] , \SUMB[24][38] , \SUMB[24][37] ,
         \SUMB[24][36] , \SUMB[24][35] , \SUMB[24][34] , \SUMB[24][33] ,
         \SUMB[24][32] , \SUMB[24][31] , \SUMB[24][30] , \SUMB[24][29] ,
         \SUMB[24][28] , \SUMB[24][27] , \SUMB[24][26] , \SUMB[24][25] ,
         \SUMB[24][24] , \SUMB[24][23] , \SUMB[24][22] , \SUMB[24][21] ,
         \SUMB[24][20] , \SUMB[24][19] , \SUMB[24][18] , \SUMB[24][17] ,
         \SUMB[24][16] , \SUMB[24][15] , \SUMB[24][14] , \SUMB[24][13] ,
         \SUMB[24][12] , \SUMB[24][11] , \SUMB[24][10] , \SUMB[24][9] ,
         \SUMB[24][8] , \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] ,
         \SUMB[24][4] , \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] ,
         \SUMB[23][46] , \SUMB[23][45] , \SUMB[23][44] , \SUMB[23][43] ,
         \SUMB[23][42] , \SUMB[23][41] , \SUMB[23][40] , \SUMB[23][39] ,
         \SUMB[23][38] , \SUMB[23][37] , \SUMB[23][36] , \SUMB[23][35] ,
         \SUMB[23][34] , \SUMB[23][33] , \SUMB[23][32] , \SUMB[23][31] ,
         \SUMB[23][30] , \SUMB[23][29] , \SUMB[23][28] , \SUMB[23][27] ,
         \SUMB[23][26] , \SUMB[23][25] , \SUMB[23][24] , \SUMB[23][23] ,
         \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] ,
         \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] ,
         \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] ,
         \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] ,
         \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] ,
         \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][46] , \SUMB[22][45] ,
         \SUMB[22][44] , \SUMB[22][43] , \SUMB[22][42] , \SUMB[22][41] ,
         \SUMB[22][40] , \SUMB[22][39] , \SUMB[22][38] , \SUMB[22][37] ,
         \SUMB[22][36] , \SUMB[22][35] , \SUMB[22][34] , \SUMB[22][33] ,
         \SUMB[22][32] , \SUMB[22][31] , \SUMB[22][30] , \SUMB[22][29] ,
         \SUMB[22][28] , \SUMB[22][27] , \SUMB[22][26] , \SUMB[22][25] ,
         \SUMB[22][24] , \SUMB[22][23] , \SUMB[22][22] , \SUMB[22][21] ,
         \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] ,
         \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][13] ,
         \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] , \SUMB[22][9] ,
         \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] ,
         \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] ,
         \SUMB[21][46] , \SUMB[21][45] , \SUMB[21][44] , \SUMB[21][43] ,
         \SUMB[21][42] , \SUMB[21][41] , \SUMB[21][40] , \SUMB[21][39] ,
         \SUMB[21][38] , \SUMB[21][37] , \SUMB[21][36] , \SUMB[21][35] ,
         \SUMB[21][34] , \SUMB[21][33] , \SUMB[21][32] , \SUMB[21][31] ,
         \SUMB[21][30] , \SUMB[21][29] , \SUMB[21][28] , \SUMB[21][27] ,
         \SUMB[21][26] , \SUMB[21][25] , \SUMB[21][24] , \SUMB[21][23] ,
         \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] , \SUMB[21][19] ,
         \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] , \SUMB[21][15] ,
         \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] , \SUMB[21][11] ,
         \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] ,
         \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] ,
         \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][46] , \SUMB[20][45] ,
         \SUMB[20][44] , \SUMB[20][43] , \SUMB[20][42] , \SUMB[20][41] ,
         \SUMB[20][40] , \SUMB[20][39] , \SUMB[20][38] , \SUMB[20][37] ,
         \SUMB[20][36] , \SUMB[20][35] , \SUMB[20][34] , \SUMB[20][33] ,
         \SUMB[20][32] , \SUMB[20][31] , \SUMB[20][30] , \SUMB[20][29] ,
         \SUMB[20][28] , \SUMB[20][27] , \SUMB[20][26] , \SUMB[20][25] ,
         \SUMB[20][24] , \SUMB[20][23] , \SUMB[20][22] , \SUMB[20][21] ,
         \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] ,
         \SUMB[20][16] , \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] ,
         \SUMB[20][12] , \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] ,
         \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] ,
         \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] ,
         \SUMB[19][46] , \SUMB[19][45] , \SUMB[19][44] , \SUMB[19][43] ,
         \SUMB[19][42] , \SUMB[19][41] , \SUMB[19][40] , \SUMB[19][39] ,
         \SUMB[19][38] , \SUMB[19][37] , \SUMB[19][36] , \SUMB[19][35] ,
         \SUMB[19][34] , \SUMB[19][33] , \SUMB[19][32] , \SUMB[19][31] ,
         \SUMB[19][30] , \SUMB[19][29] , \SUMB[19][28] , \SUMB[19][27] ,
         \SUMB[19][26] , \SUMB[19][25] , \SUMB[19][24] , \SUMB[19][23] ,
         \SUMB[19][22] , \SUMB[19][21] , \SUMB[19][20] , \SUMB[19][19] ,
         \SUMB[19][18] , \SUMB[19][17] , \SUMB[19][16] , \SUMB[19][15] ,
         \SUMB[19][14] , \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] ,
         \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][46] , \SUMB[18][45] ,
         \SUMB[18][44] , \SUMB[18][43] , \SUMB[18][42] , \SUMB[18][41] ,
         \SUMB[18][40] , \SUMB[18][39] , \SUMB[18][38] , \SUMB[18][37] ,
         \SUMB[18][36] , \SUMB[18][35] , \SUMB[18][34] , \SUMB[18][33] ,
         \SUMB[18][32] , \SUMB[18][31] , \SUMB[18][30] , \SUMB[18][29] ,
         \SUMB[18][28] , \SUMB[18][27] , \SUMB[18][26] , \SUMB[18][25] ,
         \SUMB[18][24] , \SUMB[18][23] , \SUMB[18][22] , \SUMB[18][21] ,
         \SUMB[18][20] , \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][17] ,
         \SUMB[18][16] , \SUMB[18][15] , \SUMB[18][14] , \SUMB[18][13] ,
         \SUMB[18][12] , \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] ,
         \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] ,
         \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] ,
         \SUMB[17][46] , \SUMB[17][45] , \SUMB[17][44] , \SUMB[17][43] ,
         \SUMB[17][42] , \SUMB[17][41] , \SUMB[17][40] , \SUMB[17][39] ,
         \SUMB[17][38] , \SUMB[17][37] , \SUMB[17][36] , \SUMB[17][35] ,
         \SUMB[17][34] , \SUMB[17][33] , \SUMB[17][32] , \SUMB[17][31] ,
         \SUMB[17][30] , \SUMB[17][29] , \SUMB[17][28] , \SUMB[17][27] ,
         \SUMB[17][26] , \SUMB[17][25] , \SUMB[17][24] , \SUMB[17][23] ,
         \SUMB[17][22] , \SUMB[17][21] , \SUMB[17][20] , \SUMB[17][19] ,
         \SUMB[17][18] , \SUMB[17][17] , \SUMB[17][16] , \SUMB[17][15] ,
         \SUMB[17][14] , \SUMB[17][13] , \SUMB[17][12] , \SUMB[17][11] ,
         \SUMB[17][10] , \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] ,
         \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] ,
         \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][46] , \SUMB[16][45] ,
         \SUMB[16][44] , \SUMB[16][43] , \SUMB[16][42] , \SUMB[16][41] ,
         \SUMB[16][40] , \SUMB[16][39] , \SUMB[16][38] , \SUMB[16][37] ,
         \SUMB[16][36] , \SUMB[16][35] , \SUMB[16][34] , \SUMB[16][33] ,
         \SUMB[16][32] , \SUMB[16][31] , \SUMB[16][30] , \SUMB[16][29] ,
         \SUMB[16][28] , \SUMB[16][27] , \SUMB[16][26] , \SUMB[16][25] ,
         \SUMB[16][24] , \SUMB[16][23] , \SUMB[16][22] , \SUMB[16][21] ,
         \SUMB[16][20] , \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] ,
         \SUMB[16][16] , \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] ,
         \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] ,
         \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] ,
         \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] ,
         \CARRYB[37][15] , \CARRYB[37][14] , \CARRYB[37][13] ,
         \CARRYB[37][12] , \CARRYB[37][11] , \CARRYB[37][10] , \CARRYB[37][9] ,
         \CARRYB[37][8] , \CARRYB[37][7] , \CARRYB[37][6] , \CARRYB[37][5] ,
         \CARRYB[37][4] , \CARRYB[37][3] , \CARRYB[37][2] , \CARRYB[37][1] ,
         \CARRYB[37][0] , \CARRYB[36][46] , \CARRYB[36][45] , \CARRYB[36][44] ,
         \CARRYB[36][43] , \CARRYB[36][42] , \CARRYB[36][41] ,
         \CARRYB[36][40] , \CARRYB[36][39] , \CARRYB[36][38] ,
         \CARRYB[36][37] , \CARRYB[36][36] , \CARRYB[36][35] ,
         \CARRYB[36][34] , \CARRYB[36][33] , \CARRYB[36][32] ,
         \CARRYB[36][31] , \CARRYB[36][30] , \CARRYB[36][29] ,
         \CARRYB[36][28] , \CARRYB[36][27] , \CARRYB[36][26] ,
         \CARRYB[36][25] , \CARRYB[36][24] , \CARRYB[36][23] ,
         \CARRYB[36][22] , \CARRYB[36][21] , \CARRYB[36][20] ,
         \CARRYB[36][19] , \CARRYB[36][18] , \CARRYB[36][17] ,
         \CARRYB[36][16] , \CARRYB[36][15] , \CARRYB[36][14] ,
         \CARRYB[36][13] , \CARRYB[36][12] , \CARRYB[36][11] ,
         \CARRYB[36][10] , \CARRYB[36][9] , \CARRYB[36][8] , \CARRYB[36][7] ,
         \CARRYB[36][6] , \CARRYB[36][5] , \CARRYB[36][4] , \CARRYB[36][3] ,
         \CARRYB[36][2] , \CARRYB[36][1] , \CARRYB[36][0] , \CARRYB[35][46] ,
         \CARRYB[35][45] , \CARRYB[35][44] , \CARRYB[35][43] ,
         \CARRYB[35][42] , \CARRYB[35][41] , \CARRYB[35][40] ,
         \CARRYB[35][39] , \CARRYB[35][38] , \CARRYB[35][37] ,
         \CARRYB[35][36] , \CARRYB[35][35] , \CARRYB[35][34] ,
         \CARRYB[35][33] , \CARRYB[35][32] , \CARRYB[35][31] ,
         \CARRYB[35][30] , \CARRYB[35][29] , \CARRYB[35][28] ,
         \CARRYB[35][27] , \CARRYB[35][26] , \CARRYB[35][25] ,
         \CARRYB[35][24] , \CARRYB[35][23] , \CARRYB[35][22] ,
         \CARRYB[35][21] , \CARRYB[35][20] , \CARRYB[35][19] ,
         \CARRYB[35][18] , \CARRYB[35][17] , \CARRYB[35][16] ,
         \CARRYB[35][15] , \CARRYB[35][14] , \CARRYB[35][13] ,
         \CARRYB[35][12] , \CARRYB[35][11] , \CARRYB[35][10] , \CARRYB[35][9] ,
         \CARRYB[35][8] , \CARRYB[35][7] , \CARRYB[35][6] , \CARRYB[35][5] ,
         \CARRYB[35][4] , \CARRYB[35][3] , \CARRYB[35][2] , \CARRYB[35][1] ,
         \CARRYB[35][0] , \CARRYB[34][46] , \CARRYB[34][45] , \CARRYB[34][44] ,
         \CARRYB[34][43] , \CARRYB[34][42] , \CARRYB[34][41] ,
         \CARRYB[34][40] , \CARRYB[34][39] , \CARRYB[34][38] ,
         \CARRYB[34][37] , \CARRYB[34][36] , \CARRYB[34][35] ,
         \CARRYB[34][34] , \CARRYB[34][33] , \CARRYB[34][32] ,
         \CARRYB[34][31] , \CARRYB[34][30] , \CARRYB[34][29] ,
         \CARRYB[34][28] , \CARRYB[34][27] , \CARRYB[34][26] ,
         \CARRYB[34][25] , \CARRYB[34][24] , \CARRYB[34][23] ,
         \CARRYB[34][22] , \CARRYB[34][21] , \CARRYB[34][20] ,
         \CARRYB[34][19] , \CARRYB[34][18] , \CARRYB[34][17] ,
         \CARRYB[34][16] , \CARRYB[34][15] , \CARRYB[34][14] ,
         \CARRYB[34][13] , \CARRYB[34][12] , \CARRYB[34][11] ,
         \CARRYB[34][10] , \CARRYB[34][9] , \CARRYB[34][8] , \CARRYB[34][7] ,
         \CARRYB[34][6] , \CARRYB[34][5] , \CARRYB[34][4] , \CARRYB[34][3] ,
         \CARRYB[34][2] , \CARRYB[34][1] , \CARRYB[34][0] , \CARRYB[33][46] ,
         \CARRYB[33][45] , \CARRYB[33][44] , \CARRYB[33][43] ,
         \CARRYB[33][42] , \CARRYB[33][41] , \CARRYB[33][40] ,
         \CARRYB[33][39] , \CARRYB[33][38] , \CARRYB[33][37] ,
         \CARRYB[33][36] , \CARRYB[33][35] , \CARRYB[33][34] ,
         \CARRYB[33][33] , \CARRYB[33][32] , \CARRYB[33][31] ,
         \CARRYB[33][30] , \CARRYB[33][29] , \CARRYB[33][28] ,
         \CARRYB[33][27] , \CARRYB[33][26] , \CARRYB[33][25] ,
         \CARRYB[33][24] , \CARRYB[33][23] , \CARRYB[33][22] ,
         \CARRYB[33][21] , \CARRYB[33][20] , \CARRYB[33][19] ,
         \CARRYB[33][18] , \CARRYB[33][17] , \CARRYB[33][16] ,
         \CARRYB[33][15] , \CARRYB[33][14] , \CARRYB[33][13] ,
         \CARRYB[33][12] , \CARRYB[33][11] , \CARRYB[33][10] , \CARRYB[33][9] ,
         \CARRYB[33][8] , \CARRYB[33][7] , \CARRYB[33][6] , \CARRYB[33][5] ,
         \CARRYB[33][4] , \CARRYB[33][3] , \CARRYB[33][2] , \CARRYB[33][1] ,
         \CARRYB[33][0] , \CARRYB[32][46] , \CARRYB[32][45] , \CARRYB[32][44] ,
         \CARRYB[32][43] , \CARRYB[32][42] , \CARRYB[32][41] ,
         \CARRYB[32][40] , \CARRYB[32][39] , \CARRYB[32][38] ,
         \CARRYB[32][37] , \CARRYB[32][36] , \CARRYB[32][35] ,
         \CARRYB[32][34] , \CARRYB[32][33] , \CARRYB[32][32] ,
         \CARRYB[32][31] , \CARRYB[32][30] , \CARRYB[32][29] ,
         \CARRYB[32][28] , \CARRYB[32][27] , \CARRYB[32][26] ,
         \CARRYB[32][25] , \CARRYB[32][24] , \CARRYB[32][23] ,
         \CARRYB[32][22] , \CARRYB[32][21] , \CARRYB[32][20] ,
         \CARRYB[32][19] , \CARRYB[32][18] , \CARRYB[32][17] ,
         \CARRYB[32][16] , \CARRYB[32][15] , \CARRYB[32][14] ,
         \CARRYB[32][13] , \CARRYB[32][12] , \CARRYB[32][11] ,
         \CARRYB[32][10] , \CARRYB[32][9] , \CARRYB[32][8] , \CARRYB[32][7] ,
         \CARRYB[32][6] , \CARRYB[32][5] , \CARRYB[32][4] , \CARRYB[32][3] ,
         \CARRYB[32][2] , \CARRYB[32][1] , \CARRYB[32][0] , \CARRYB[31][46] ,
         \CARRYB[31][45] , \CARRYB[31][44] , \CARRYB[31][43] ,
         \CARRYB[31][42] , \CARRYB[31][41] , \CARRYB[31][40] ,
         \CARRYB[31][39] , \CARRYB[31][38] , \CARRYB[31][37] ,
         \CARRYB[31][36] , \CARRYB[31][35] , \CARRYB[31][34] ,
         \CARRYB[31][33] , \CARRYB[31][32] , \CARRYB[31][31] ,
         \CARRYB[31][30] , \CARRYB[31][29] , \CARRYB[31][28] ,
         \CARRYB[31][27] , \CARRYB[31][26] , \CARRYB[31][25] ,
         \CARRYB[31][24] , \CARRYB[31][23] , \CARRYB[31][22] ,
         \CARRYB[31][21] , \CARRYB[31][20] , \CARRYB[31][19] ,
         \CARRYB[31][18] , \CARRYB[31][17] , \CARRYB[31][16] ,
         \CARRYB[31][15] , \CARRYB[31][14] , \CARRYB[31][13] ,
         \CARRYB[31][12] , \CARRYB[31][11] , \CARRYB[31][10] , \CARRYB[31][9] ,
         \CARRYB[31][8] , \CARRYB[31][7] , \CARRYB[31][6] , \CARRYB[31][5] ,
         \CARRYB[31][4] , \CARRYB[31][3] , \CARRYB[31][2] , \CARRYB[31][1] ,
         \CARRYB[31][0] , \CARRYB[30][46] , \CARRYB[30][45] , \CARRYB[30][44] ,
         \CARRYB[30][43] , \CARRYB[30][42] , \CARRYB[30][41] ,
         \CARRYB[30][40] , \CARRYB[30][39] , \CARRYB[30][38] ,
         \CARRYB[30][37] , \CARRYB[30][36] , \CARRYB[30][35] ,
         \CARRYB[30][34] , \CARRYB[30][33] , \CARRYB[30][32] ,
         \CARRYB[30][31] , \CARRYB[30][30] , \CARRYB[30][29] ,
         \CARRYB[30][28] , \CARRYB[30][27] , \CARRYB[30][26] ,
         \CARRYB[30][25] , \CARRYB[30][24] , \CARRYB[30][23] ,
         \CARRYB[30][22] , \CARRYB[30][21] , \CARRYB[30][20] ,
         \CARRYB[30][19] , \CARRYB[30][18] , \CARRYB[30][17] ,
         \CARRYB[30][16] , \CARRYB[30][15] , \CARRYB[30][14] ,
         \CARRYB[30][13] , \CARRYB[30][12] , \CARRYB[30][11] ,
         \CARRYB[30][10] , \CARRYB[30][9] , \CARRYB[30][8] , \CARRYB[30][7] ,
         \CARRYB[30][6] , \CARRYB[30][5] , \CARRYB[30][4] , \CARRYB[30][3] ,
         \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] , \CARRYB[29][46] ,
         \CARRYB[29][45] , \CARRYB[29][44] , \CARRYB[29][43] ,
         \CARRYB[29][42] , \CARRYB[29][41] , \CARRYB[29][40] ,
         \CARRYB[29][39] , \CARRYB[29][38] , \CARRYB[29][37] ,
         \CARRYB[29][36] , \CARRYB[29][35] , \CARRYB[29][34] ,
         \CARRYB[29][33] , \CARRYB[29][32] , \CARRYB[29][31] ,
         \CARRYB[29][30] , \CARRYB[29][29] , \CARRYB[29][28] ,
         \CARRYB[29][27] , \CARRYB[29][26] , \CARRYB[29][25] ,
         \CARRYB[29][24] , \CARRYB[29][23] , \CARRYB[29][22] ,
         \CARRYB[29][21] , \CARRYB[29][20] , \CARRYB[29][19] ,
         \CARRYB[29][18] , \CARRYB[29][17] , \CARRYB[29][16] ,
         \CARRYB[29][15] , \CARRYB[29][14] , \CARRYB[29][13] ,
         \CARRYB[29][12] , \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] ,
         \CARRYB[29][4] , \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][46] , \CARRYB[28][45] , \CARRYB[28][44] ,
         \CARRYB[28][43] , \CARRYB[28][42] , \CARRYB[28][41] ,
         \CARRYB[28][40] , \CARRYB[28][39] , \CARRYB[28][38] ,
         \CARRYB[28][37] , \CARRYB[28][36] , \CARRYB[28][35] ,
         \CARRYB[28][34] , \CARRYB[28][33] , \CARRYB[28][32] ,
         \CARRYB[28][31] , \CARRYB[28][30] , \CARRYB[28][29] ,
         \CARRYB[28][28] , \CARRYB[28][27] , \CARRYB[28][26] ,
         \CARRYB[28][25] , \CARRYB[28][24] , \CARRYB[28][23] ,
         \CARRYB[28][22] , \CARRYB[28][21] , \CARRYB[28][20] ,
         \CARRYB[28][19] , \CARRYB[28][18] , \CARRYB[28][17] ,
         \CARRYB[28][16] , \CARRYB[28][15] , \CARRYB[28][14] ,
         \CARRYB[28][13] , \CARRYB[28][12] , \CARRYB[28][11] ,
         \CARRYB[28][10] , \CARRYB[28][9] , \CARRYB[28][8] , \CARRYB[28][7] ,
         \CARRYB[28][6] , \CARRYB[28][5] , \CARRYB[28][4] , \CARRYB[28][3] ,
         \CARRYB[28][2] , \CARRYB[28][1] , \CARRYB[28][0] , \CARRYB[27][46] ,
         \CARRYB[27][45] , \CARRYB[27][44] , \CARRYB[27][43] ,
         \CARRYB[27][42] , \CARRYB[27][41] , \CARRYB[27][40] ,
         \CARRYB[27][39] , \CARRYB[27][38] , \CARRYB[27][37] ,
         \CARRYB[27][36] , \CARRYB[27][35] , \CARRYB[27][34] ,
         \CARRYB[27][33] , \CARRYB[27][32] , \CARRYB[27][31] ,
         \CARRYB[27][30] , \CARRYB[27][29] , \CARRYB[27][28] ,
         \CARRYB[27][27] , \CARRYB[27][26] , \CARRYB[27][25] ,
         \CARRYB[27][24] , \CARRYB[27][23] , \CARRYB[27][22] ,
         \CARRYB[27][21] , \CARRYB[27][20] , \CARRYB[27][19] ,
         \CARRYB[27][18] , \CARRYB[27][17] , \CARRYB[27][16] ,
         \CARRYB[27][15] , \CARRYB[27][14] , \CARRYB[27][13] ,
         \CARRYB[27][12] , \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] ,
         \CARRYB[27][8] , \CARRYB[27][7] , \CARRYB[27][6] , \CARRYB[27][5] ,
         \CARRYB[27][4] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][46] , \CARRYB[26][45] , \CARRYB[26][44] ,
         \CARRYB[26][43] , \CARRYB[26][42] , \CARRYB[26][41] ,
         \CARRYB[26][40] , \CARRYB[26][39] , \CARRYB[26][38] ,
         \CARRYB[26][37] , \CARRYB[26][36] , \CARRYB[26][35] ,
         \CARRYB[26][34] , \CARRYB[26][33] , \CARRYB[26][32] , \SUMB[37][15] ,
         \SUMB[37][14] , \SUMB[37][13] , \SUMB[37][12] , \SUMB[37][11] ,
         \SUMB[37][10] , \SUMB[37][9] , \SUMB[37][8] , \SUMB[37][7] ,
         \SUMB[37][6] , \SUMB[37][5] , \SUMB[37][4] , \SUMB[37][3] ,
         \SUMB[37][2] , \SUMB[37][1] , \SUMB[36][46] , \SUMB[36][45] ,
         \SUMB[36][44] , \SUMB[36][43] , \SUMB[36][42] , \SUMB[36][41] ,
         \SUMB[36][40] , \SUMB[36][39] , \SUMB[36][38] , \SUMB[36][37] ,
         \SUMB[36][36] , \SUMB[36][35] , \SUMB[36][34] , \SUMB[36][33] ,
         \SUMB[36][32] , \SUMB[36][31] , \SUMB[36][30] , \SUMB[36][29] ,
         \SUMB[36][28] , \SUMB[36][27] , \SUMB[36][26] , \SUMB[36][25] ,
         \SUMB[36][24] , \SUMB[36][23] , \SUMB[36][22] , \SUMB[36][21] ,
         \SUMB[36][20] , \SUMB[36][19] , \SUMB[36][18] , \SUMB[36][17] ,
         \SUMB[36][16] , \SUMB[36][15] , \SUMB[36][14] , \SUMB[36][13] ,
         \SUMB[36][12] , \SUMB[36][11] , \SUMB[36][10] , \SUMB[36][9] ,
         \SUMB[36][8] , \SUMB[36][7] , \SUMB[36][6] , \SUMB[36][5] ,
         \SUMB[36][4] , \SUMB[36][3] , \SUMB[36][2] , \SUMB[36][1] ,
         \SUMB[35][46] , \SUMB[35][45] , \SUMB[35][44] , \SUMB[35][43] ,
         \SUMB[35][42] , \SUMB[35][41] , \SUMB[35][40] , \SUMB[35][39] ,
         \SUMB[35][38] , \SUMB[35][37] , \SUMB[35][36] , \SUMB[35][35] ,
         \SUMB[35][34] , \SUMB[35][33] , \SUMB[35][32] , \SUMB[35][31] ,
         \SUMB[35][30] , \SUMB[35][29] , \SUMB[35][28] , \SUMB[35][27] ,
         \SUMB[35][26] , \SUMB[35][25] , \SUMB[35][24] , \SUMB[35][23] ,
         \SUMB[35][22] , \SUMB[35][21] , \SUMB[35][20] , \SUMB[35][19] ,
         \SUMB[35][18] , \SUMB[35][17] , \SUMB[35][16] , \SUMB[35][15] ,
         \SUMB[35][14] , \SUMB[35][13] , \SUMB[35][12] , \SUMB[35][11] ,
         \SUMB[35][10] , \SUMB[35][9] , \SUMB[35][8] , \SUMB[35][7] ,
         \SUMB[35][6] , \SUMB[35][5] , \SUMB[35][4] , \SUMB[35][3] ,
         \SUMB[35][2] , \SUMB[35][1] , \SUMB[34][46] , \SUMB[34][45] ,
         \SUMB[34][44] , \SUMB[34][43] , \SUMB[34][42] , \SUMB[34][41] ,
         \SUMB[34][40] , \SUMB[34][39] , \SUMB[34][38] , \SUMB[34][37] ,
         \SUMB[34][36] , \SUMB[34][35] , \SUMB[34][34] , \SUMB[34][33] ,
         \SUMB[34][32] , \SUMB[34][31] , \SUMB[34][30] , \SUMB[34][29] ,
         \SUMB[34][28] , \SUMB[34][27] , \SUMB[34][26] , \SUMB[34][25] ,
         \SUMB[34][24] , \SUMB[34][23] , \SUMB[34][22] , \SUMB[34][21] ,
         \SUMB[34][20] , \SUMB[34][19] , \SUMB[34][18] , \SUMB[34][17] ,
         \SUMB[34][16] , \SUMB[34][15] , \SUMB[34][14] , \SUMB[34][13] ,
         \SUMB[34][12] , \SUMB[34][11] , \SUMB[34][10] , \SUMB[34][9] ,
         \SUMB[34][8] , \SUMB[34][7] , \SUMB[34][6] , \SUMB[34][5] ,
         \SUMB[34][4] , \SUMB[34][3] , \SUMB[34][2] , \SUMB[34][1] ,
         \SUMB[33][46] , \SUMB[33][45] , \SUMB[33][44] , \SUMB[33][43] ,
         \SUMB[33][42] , \SUMB[33][41] , \SUMB[33][40] , \SUMB[33][39] ,
         \SUMB[33][38] , \SUMB[33][37] , \SUMB[33][36] , \SUMB[33][35] ,
         \SUMB[33][34] , \SUMB[33][33] , \SUMB[33][32] , \SUMB[33][31] ,
         \SUMB[33][30] , \SUMB[33][29] , \SUMB[33][28] , \SUMB[33][27] ,
         \SUMB[33][26] , \SUMB[33][25] , \SUMB[33][24] , \SUMB[33][23] ,
         \SUMB[33][22] , \SUMB[33][21] , \SUMB[33][20] , \SUMB[33][19] ,
         \SUMB[33][18] , \SUMB[33][17] , \SUMB[33][16] , \SUMB[33][15] ,
         \SUMB[33][14] , \SUMB[33][13] , \SUMB[33][12] , \SUMB[33][11] ,
         \SUMB[33][10] , \SUMB[33][9] , \SUMB[33][8] , \SUMB[33][7] ,
         \SUMB[33][6] , \SUMB[33][5] , \SUMB[33][4] , \SUMB[33][3] ,
         \SUMB[33][2] , \SUMB[33][1] , \SUMB[32][46] , \SUMB[32][45] ,
         \SUMB[32][44] , \SUMB[32][43] , \SUMB[32][42] , \SUMB[32][41] ,
         \SUMB[32][40] , \SUMB[32][39] , \SUMB[32][38] , \SUMB[32][37] ,
         \SUMB[32][36] , \SUMB[32][35] , \SUMB[32][34] , \SUMB[32][33] ,
         \SUMB[32][32] , \SUMB[32][31] , \SUMB[32][30] , \SUMB[32][29] ,
         \SUMB[32][28] , \SUMB[32][27] , \SUMB[32][26] , \SUMB[32][25] ,
         \SUMB[32][24] , \SUMB[32][23] , \SUMB[32][22] , \SUMB[32][21] ,
         \SUMB[32][20] , \SUMB[32][19] , \SUMB[32][18] , \SUMB[32][17] ,
         \SUMB[32][16] , \SUMB[32][15] , \SUMB[32][14] , \SUMB[32][13] ,
         \SUMB[32][12] , \SUMB[32][11] , \SUMB[32][10] , \SUMB[32][9] ,
         \SUMB[32][8] , \SUMB[32][7] , \SUMB[32][6] , \SUMB[32][5] ,
         \SUMB[32][4] , \SUMB[32][3] , \SUMB[32][2] , \SUMB[32][1] ,
         \SUMB[31][46] , \SUMB[31][45] , \SUMB[31][44] , \SUMB[31][43] ,
         \SUMB[31][42] , \SUMB[31][41] , \SUMB[31][40] , \SUMB[31][39] ,
         \SUMB[31][38] , \SUMB[31][37] , \SUMB[31][36] , \SUMB[31][35] ,
         \SUMB[31][34] , \SUMB[31][33] , \SUMB[31][32] , \SUMB[31][31] ,
         \SUMB[31][30] , \SUMB[31][29] , \SUMB[31][28] , \SUMB[31][27] ,
         \SUMB[31][26] , \SUMB[31][25] , \SUMB[31][24] , \SUMB[31][23] ,
         \SUMB[31][22] , \SUMB[31][21] , \SUMB[31][20] , \SUMB[31][19] ,
         \SUMB[31][18] , \SUMB[31][17] , \SUMB[31][16] , \SUMB[31][15] ,
         \SUMB[31][14] , \SUMB[31][13] , \SUMB[31][12] , \SUMB[31][11] ,
         \SUMB[31][10] , \SUMB[31][9] , \SUMB[31][8] , \SUMB[31][7] ,
         \SUMB[31][6] , \SUMB[31][5] , \SUMB[31][4] , \SUMB[31][3] ,
         \SUMB[31][2] , \SUMB[31][1] , \SUMB[30][46] , \SUMB[30][45] ,
         \SUMB[30][44] , \SUMB[30][43] , \SUMB[30][42] , \SUMB[30][41] ,
         \SUMB[30][40] , \SUMB[30][39] , \SUMB[30][38] , \SUMB[30][37] ,
         \SUMB[30][36] , \SUMB[30][35] , \SUMB[30][34] , \SUMB[30][33] ,
         \SUMB[30][32] , \SUMB[30][31] , \SUMB[30][30] , \SUMB[30][29] ,
         \SUMB[30][28] , \SUMB[30][27] , \SUMB[30][26] , \SUMB[30][25] ,
         \SUMB[30][24] , \SUMB[30][23] , \SUMB[30][22] , \SUMB[30][21] ,
         \SUMB[30][20] , \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] ,
         \SUMB[30][16] , \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] ,
         \SUMB[30][12] , \SUMB[30][11] , \SUMB[30][10] , \SUMB[30][9] ,
         \SUMB[30][8] , \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] ,
         \SUMB[30][4] , \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] ,
         \SUMB[29][46] , \SUMB[29][45] , \SUMB[29][44] , \SUMB[29][43] ,
         \SUMB[29][42] , \SUMB[29][41] , \SUMB[29][40] , \SUMB[29][39] ,
         \SUMB[29][38] , \SUMB[29][37] , \SUMB[29][36] , \SUMB[29][35] ,
         \SUMB[29][34] , \SUMB[29][33] , \SUMB[29][32] , \SUMB[29][31] ,
         \SUMB[29][30] , \SUMB[29][29] , \SUMB[29][28] , \SUMB[29][27] ,
         \SUMB[29][26] , \SUMB[29][25] , \SUMB[29][24] , \SUMB[29][23] ,
         \SUMB[29][22] , \SUMB[29][21] , \SUMB[29][20] , \SUMB[29][19] ,
         \SUMB[29][18] , \SUMB[29][17] , \SUMB[29][16] , \SUMB[29][15] ,
         \SUMB[29][14] , \SUMB[29][13] , \SUMB[29][12] , \SUMB[29][11] ,
         \SUMB[29][10] , \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] ,
         \SUMB[29][6] , \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] ,
         \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][46] , \SUMB[28][45] ,
         \SUMB[28][44] , \SUMB[28][43] , \SUMB[28][42] , \SUMB[28][41] ,
         \SUMB[28][40] , \SUMB[28][39] , \SUMB[28][38] , \SUMB[28][37] ,
         \SUMB[28][36] , \SUMB[28][35] , \SUMB[28][34] , \SUMB[28][33] ,
         \SUMB[28][32] , \SUMB[28][31] , \SUMB[28][30] , \SUMB[28][29] ,
         \SUMB[28][28] , \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] ,
         \SUMB[28][24] , \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] ,
         \SUMB[28][20] , \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] ,
         \SUMB[28][16] , \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] ,
         \SUMB[28][12] , \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] ,
         \SUMB[28][8] , \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] ,
         \SUMB[28][4] , \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] ,
         \SUMB[27][46] , \SUMB[27][45] , \SUMB[27][44] , \SUMB[27][43] ,
         \SUMB[27][42] , \SUMB[27][41] , \SUMB[27][40] , \SUMB[27][39] ,
         \SUMB[27][38] , \SUMB[27][37] , \SUMB[27][36] , \SUMB[27][35] ,
         \SUMB[27][34] , \SUMB[27][33] , \SUMB[27][32] , \SUMB[27][31] ,
         \SUMB[27][30] , \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] ,
         \SUMB[27][26] , \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] ,
         \SUMB[27][22] , \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] ,
         \SUMB[27][18] , \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] ,
         \SUMB[27][14] , \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] ,
         \SUMB[27][10] , \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] ,
         \SUMB[27][6] , \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][46] , \SUMB[26][45] ,
         \SUMB[26][44] , \SUMB[26][43] , \SUMB[26][42] , \SUMB[26][41] ,
         \SUMB[26][40] , \SUMB[26][39] , \SUMB[26][38] , \SUMB[26][37] ,
         \SUMB[26][36] , \SUMB[26][35] , \SUMB[26][34] , \SUMB[26][33] ,
         \SUMB[26][32] , \CARRYB[47][46] , \CARRYB[47][45] , \CARRYB[47][44] ,
         \CARRYB[47][43] , \CARRYB[47][42] , \CARRYB[47][41] ,
         \CARRYB[47][40] , \CARRYB[47][39] , \CARRYB[47][38] ,
         \CARRYB[47][37] , \CARRYB[47][36] , \CARRYB[47][35] ,
         \CARRYB[47][34] , \CARRYB[47][33] , \CARRYB[47][32] ,
         \CARRYB[47][31] , \CARRYB[47][30] , \CARRYB[47][29] ,
         \CARRYB[47][28] , \CARRYB[47][27] , \CARRYB[47][26] ,
         \CARRYB[47][25] , \CARRYB[47][24] , \CARRYB[47][23] ,
         \CARRYB[47][22] , \CARRYB[47][21] , \CARRYB[47][20] ,
         \CARRYB[47][19] , \CARRYB[47][18] , \CARRYB[47][17] ,
         \CARRYB[47][16] , \CARRYB[47][15] , \CARRYB[47][14] ,
         \CARRYB[47][13] , \CARRYB[47][12] , \CARRYB[47][11] ,
         \CARRYB[47][10] , \CARRYB[47][9] , \CARRYB[47][8] , \CARRYB[47][7] ,
         \CARRYB[47][6] , \CARRYB[47][5] , \CARRYB[47][4] , \CARRYB[47][3] ,
         \CARRYB[47][2] , \CARRYB[47][1] , \CARRYB[47][0] , \CARRYB[46][46] ,
         \CARRYB[46][45] , \CARRYB[46][44] , \CARRYB[46][43] ,
         \CARRYB[46][42] , \CARRYB[46][41] , \CARRYB[46][40] ,
         \CARRYB[46][39] , \CARRYB[46][38] , \CARRYB[46][37] ,
         \CARRYB[46][36] , \CARRYB[46][35] , \CARRYB[46][34] ,
         \CARRYB[46][33] , \CARRYB[46][32] , \CARRYB[46][31] ,
         \CARRYB[46][30] , \CARRYB[46][29] , \CARRYB[46][28] ,
         \CARRYB[46][27] , \CARRYB[46][26] , \CARRYB[46][25] ,
         \CARRYB[46][24] , \CARRYB[46][23] , \CARRYB[46][22] ,
         \CARRYB[46][21] , \CARRYB[46][20] , \CARRYB[46][19] ,
         \CARRYB[46][18] , \CARRYB[46][17] , \CARRYB[46][16] ,
         \CARRYB[46][15] , \CARRYB[46][14] , \CARRYB[46][13] ,
         \CARRYB[46][12] , \CARRYB[46][11] , \CARRYB[46][10] , \CARRYB[46][9] ,
         \CARRYB[46][8] , \CARRYB[46][7] , \CARRYB[46][6] , \CARRYB[46][5] ,
         \CARRYB[46][4] , \CARRYB[46][3] , \CARRYB[46][2] , \CARRYB[46][1] ,
         \CARRYB[46][0] , \CARRYB[45][46] , \CARRYB[45][45] , \CARRYB[45][44] ,
         \CARRYB[45][43] , \CARRYB[45][42] , \CARRYB[45][41] ,
         \CARRYB[45][40] , \CARRYB[45][39] , \CARRYB[45][38] ,
         \CARRYB[45][37] , \CARRYB[45][36] , \CARRYB[45][35] ,
         \CARRYB[45][34] , \CARRYB[45][33] , \CARRYB[45][32] ,
         \CARRYB[45][31] , \CARRYB[45][30] , \CARRYB[45][29] ,
         \CARRYB[45][28] , \CARRYB[45][27] , \CARRYB[45][26] ,
         \CARRYB[45][25] , \CARRYB[45][24] , \CARRYB[45][23] ,
         \CARRYB[45][22] , \CARRYB[45][21] , \CARRYB[45][20] ,
         \CARRYB[45][19] , \CARRYB[45][18] , \CARRYB[45][17] ,
         \CARRYB[45][16] , \CARRYB[45][15] , \CARRYB[45][14] ,
         \CARRYB[45][13] , \CARRYB[45][12] , \CARRYB[45][11] ,
         \CARRYB[45][10] , \CARRYB[45][9] , \CARRYB[45][8] , \CARRYB[45][7] ,
         \CARRYB[45][6] , \CARRYB[45][5] , \CARRYB[45][4] , \CARRYB[45][3] ,
         \CARRYB[45][2] , \CARRYB[45][1] , \CARRYB[45][0] , \CARRYB[44][46] ,
         \CARRYB[44][45] , \CARRYB[44][44] , \CARRYB[44][43] ,
         \CARRYB[44][42] , \CARRYB[44][41] , \CARRYB[44][40] ,
         \CARRYB[44][39] , \CARRYB[44][38] , \CARRYB[44][37] ,
         \CARRYB[44][36] , \CARRYB[44][35] , \CARRYB[44][34] ,
         \CARRYB[44][33] , \CARRYB[44][32] , \CARRYB[44][31] ,
         \CARRYB[44][30] , \CARRYB[44][29] , \CARRYB[44][28] ,
         \CARRYB[44][27] , \CARRYB[44][26] , \CARRYB[44][25] ,
         \CARRYB[44][24] , \CARRYB[44][23] , \CARRYB[44][22] ,
         \CARRYB[44][21] , \CARRYB[44][20] , \CARRYB[44][19] ,
         \CARRYB[44][18] , \CARRYB[44][17] , \CARRYB[44][16] ,
         \CARRYB[44][15] , \CARRYB[44][14] , \CARRYB[44][13] ,
         \CARRYB[44][12] , \CARRYB[44][11] , \CARRYB[44][10] , \CARRYB[44][9] ,
         \CARRYB[44][8] , \CARRYB[44][7] , \CARRYB[44][6] , \CARRYB[44][5] ,
         \CARRYB[44][4] , \CARRYB[44][3] , \CARRYB[44][2] , \CARRYB[44][1] ,
         \CARRYB[44][0] , \CARRYB[43][46] , \CARRYB[43][45] , \CARRYB[43][44] ,
         \CARRYB[43][43] , \CARRYB[43][42] , \CARRYB[43][41] ,
         \CARRYB[43][40] , \CARRYB[43][39] , \CARRYB[43][38] ,
         \CARRYB[43][37] , \CARRYB[43][36] , \CARRYB[43][35] ,
         \CARRYB[43][34] , \CARRYB[43][33] , \CARRYB[43][32] ,
         \CARRYB[43][31] , \CARRYB[43][30] , \CARRYB[43][29] ,
         \CARRYB[43][28] , \CARRYB[43][27] , \CARRYB[43][26] ,
         \CARRYB[43][25] , \CARRYB[43][24] , \CARRYB[43][23] ,
         \CARRYB[43][22] , \CARRYB[43][21] , \CARRYB[43][20] ,
         \CARRYB[43][19] , \CARRYB[43][18] , \CARRYB[43][17] ,
         \CARRYB[43][16] , \CARRYB[43][15] , \CARRYB[43][14] ,
         \CARRYB[43][13] , \CARRYB[43][12] , \CARRYB[43][11] ,
         \CARRYB[43][10] , \CARRYB[43][9] , \CARRYB[43][8] , \CARRYB[43][7] ,
         \CARRYB[43][6] , \CARRYB[43][5] , \CARRYB[43][4] , \CARRYB[43][3] ,
         \CARRYB[43][2] , \CARRYB[43][1] , \CARRYB[43][0] , \CARRYB[42][46] ,
         \CARRYB[42][45] , \CARRYB[42][44] , \CARRYB[42][43] ,
         \CARRYB[42][42] , \CARRYB[42][41] , \CARRYB[42][40] ,
         \CARRYB[42][39] , \CARRYB[42][38] , \CARRYB[42][37] ,
         \CARRYB[42][36] , \CARRYB[42][35] , \CARRYB[42][34] ,
         \CARRYB[42][33] , \CARRYB[42][32] , \CARRYB[42][31] ,
         \CARRYB[42][30] , \CARRYB[42][29] , \CARRYB[42][28] ,
         \CARRYB[42][27] , \CARRYB[42][26] , \CARRYB[42][25] ,
         \CARRYB[42][24] , \CARRYB[42][23] , \CARRYB[42][22] ,
         \CARRYB[42][21] , \CARRYB[42][20] , \CARRYB[42][19] ,
         \CARRYB[42][18] , \CARRYB[42][17] , \CARRYB[42][16] ,
         \CARRYB[42][15] , \CARRYB[42][14] , \CARRYB[42][13] ,
         \CARRYB[42][12] , \CARRYB[42][11] , \CARRYB[42][10] , \CARRYB[42][9] ,
         \CARRYB[42][8] , \CARRYB[42][7] , \CARRYB[42][6] , \CARRYB[42][5] ,
         \CARRYB[42][4] , \CARRYB[42][3] , \CARRYB[42][2] , \CARRYB[42][1] ,
         \CARRYB[42][0] , \CARRYB[41][46] , \CARRYB[41][45] , \CARRYB[41][44] ,
         \CARRYB[41][43] , \CARRYB[41][42] , \CARRYB[41][41] ,
         \CARRYB[41][40] , \CARRYB[41][39] , \CARRYB[41][38] ,
         \CARRYB[41][37] , \CARRYB[41][36] , \CARRYB[41][35] ,
         \CARRYB[41][34] , \CARRYB[41][33] , \CARRYB[41][32] ,
         \CARRYB[41][31] , \CARRYB[41][30] , \CARRYB[41][29] ,
         \CARRYB[41][28] , \CARRYB[41][27] , \CARRYB[41][26] ,
         \CARRYB[41][25] , \CARRYB[41][24] , \CARRYB[41][23] ,
         \CARRYB[41][22] , \CARRYB[41][21] , \CARRYB[41][20] ,
         \CARRYB[41][19] , \CARRYB[41][18] , \CARRYB[41][17] ,
         \CARRYB[41][16] , \CARRYB[41][15] , \CARRYB[41][14] ,
         \CARRYB[41][13] , \CARRYB[41][12] , \CARRYB[41][11] ,
         \CARRYB[41][10] , \CARRYB[41][9] , \CARRYB[41][8] , \CARRYB[41][7] ,
         \CARRYB[41][6] , \CARRYB[41][5] , \CARRYB[41][4] , \CARRYB[41][3] ,
         \CARRYB[41][2] , \CARRYB[41][1] , \CARRYB[41][0] , \CARRYB[40][46] ,
         \CARRYB[40][45] , \CARRYB[40][44] , \CARRYB[40][43] ,
         \CARRYB[40][42] , \CARRYB[40][41] , \CARRYB[40][40] ,
         \CARRYB[40][39] , \CARRYB[40][38] , \CARRYB[40][37] ,
         \CARRYB[40][36] , \CARRYB[40][35] , \CARRYB[40][34] ,
         \CARRYB[40][33] , \CARRYB[40][32] , \CARRYB[40][31] ,
         \CARRYB[40][30] , \CARRYB[40][29] , \CARRYB[40][28] ,
         \CARRYB[40][27] , \CARRYB[40][26] , \CARRYB[40][25] ,
         \CARRYB[40][24] , \CARRYB[40][23] , \CARRYB[40][22] ,
         \CARRYB[40][21] , \CARRYB[40][20] , \CARRYB[40][19] ,
         \CARRYB[40][18] , \CARRYB[40][17] , \CARRYB[40][16] ,
         \CARRYB[40][15] , \CARRYB[40][14] , \CARRYB[40][13] ,
         \CARRYB[40][12] , \CARRYB[40][11] , \CARRYB[40][10] , \CARRYB[40][9] ,
         \CARRYB[40][8] , \CARRYB[40][7] , \CARRYB[40][6] , \CARRYB[40][5] ,
         \CARRYB[40][4] , \CARRYB[40][3] , \CARRYB[40][2] , \CARRYB[40][1] ,
         \CARRYB[40][0] , \CARRYB[39][46] , \CARRYB[39][45] , \CARRYB[39][44] ,
         \CARRYB[39][43] , \CARRYB[39][42] , \CARRYB[39][41] ,
         \CARRYB[39][40] , \CARRYB[39][39] , \CARRYB[39][38] ,
         \CARRYB[39][37] , \CARRYB[39][36] , \CARRYB[39][35] ,
         \CARRYB[39][34] , \CARRYB[39][33] , \CARRYB[39][32] ,
         \CARRYB[39][31] , \CARRYB[39][30] , \CARRYB[39][29] ,
         \CARRYB[39][28] , \CARRYB[39][27] , \CARRYB[39][26] ,
         \CARRYB[39][25] , \CARRYB[39][24] , \CARRYB[39][23] ,
         \CARRYB[39][22] , \CARRYB[39][21] , \CARRYB[39][20] ,
         \CARRYB[39][19] , \CARRYB[39][18] , \CARRYB[39][17] ,
         \CARRYB[39][16] , \CARRYB[39][15] , \CARRYB[39][14] ,
         \CARRYB[39][13] , \CARRYB[39][12] , \CARRYB[39][11] ,
         \CARRYB[39][10] , \CARRYB[39][9] , \CARRYB[39][8] , \CARRYB[39][7] ,
         \CARRYB[39][6] , \CARRYB[39][5] , \CARRYB[39][4] , \CARRYB[39][3] ,
         \CARRYB[39][2] , \CARRYB[39][1] , \CARRYB[39][0] , \CARRYB[38][46] ,
         \CARRYB[38][45] , \CARRYB[38][44] , \CARRYB[38][43] ,
         \CARRYB[38][42] , \CARRYB[38][41] , \CARRYB[38][40] ,
         \CARRYB[38][39] , \CARRYB[38][38] , \CARRYB[38][37] ,
         \CARRYB[38][36] , \CARRYB[38][35] , \CARRYB[38][34] ,
         \CARRYB[38][33] , \CARRYB[38][32] , \CARRYB[38][31] ,
         \CARRYB[38][30] , \CARRYB[38][29] , \CARRYB[38][28] ,
         \CARRYB[38][27] , \CARRYB[38][26] , \CARRYB[38][25] ,
         \CARRYB[38][24] , \CARRYB[38][23] , \CARRYB[38][22] ,
         \CARRYB[38][21] , \CARRYB[38][20] , \CARRYB[38][19] ,
         \CARRYB[38][18] , \CARRYB[38][17] , \CARRYB[38][16] ,
         \CARRYB[38][15] , \CARRYB[38][14] , \CARRYB[38][13] ,
         \CARRYB[38][12] , \CARRYB[38][11] , \CARRYB[38][10] , \CARRYB[38][9] ,
         \CARRYB[38][8] , \CARRYB[38][7] , \CARRYB[38][6] , \CARRYB[38][5] ,
         \CARRYB[38][4] , \CARRYB[38][3] , \CARRYB[38][2] , \CARRYB[38][1] ,
         \CARRYB[38][0] , \CARRYB[37][46] , \CARRYB[37][45] , \CARRYB[37][44] ,
         \CARRYB[37][43] , \CARRYB[37][42] , \CARRYB[37][41] ,
         \CARRYB[37][40] , \CARRYB[37][39] , \CARRYB[37][38] ,
         \CARRYB[37][37] , \CARRYB[37][36] , \CARRYB[37][35] ,
         \CARRYB[37][34] , \CARRYB[37][33] , \CARRYB[37][32] ,
         \CARRYB[37][31] , \CARRYB[37][30] , \CARRYB[37][29] ,
         \CARRYB[37][28] , \CARRYB[37][27] , \CARRYB[37][26] ,
         \CARRYB[37][25] , \CARRYB[37][24] , \CARRYB[37][23] ,
         \CARRYB[37][22] , \CARRYB[37][21] , \CARRYB[37][20] ,
         \CARRYB[37][19] , \CARRYB[37][18] , \CARRYB[37][17] ,
         \CARRYB[37][16] , \SUMB[47][45] , \SUMB[47][44] , \SUMB[47][43] ,
         \SUMB[47][42] , \SUMB[47][41] , \SUMB[47][40] , \SUMB[47][39] ,
         \SUMB[47][38] , \SUMB[47][37] , \SUMB[47][36] , \SUMB[47][35] ,
         \SUMB[47][34] , \SUMB[47][33] , \SUMB[47][32] , \SUMB[47][31] ,
         \SUMB[47][30] , \SUMB[47][29] , \SUMB[47][28] , \SUMB[47][27] ,
         \SUMB[47][26] , \SUMB[47][25] , \SUMB[47][24] , \SUMB[47][23] ,
         \SUMB[47][22] , \SUMB[47][21] , \SUMB[47][20] , \SUMB[47][19] ,
         \SUMB[47][18] , \SUMB[47][17] , \SUMB[47][16] , \SUMB[47][15] ,
         \SUMB[47][14] , \SUMB[47][13] , \SUMB[47][12] , \SUMB[47][11] ,
         \SUMB[47][10] , \SUMB[47][9] , \SUMB[47][8] , \SUMB[47][7] ,
         \SUMB[47][6] , \SUMB[47][5] , \SUMB[47][4] , \SUMB[47][3] ,
         \SUMB[47][2] , \SUMB[47][1] , \SUMB[47][0] , \SUMB[46][46] ,
         \SUMB[46][45] , \SUMB[46][44] , \SUMB[46][43] , \SUMB[46][42] ,
         \SUMB[46][41] , \SUMB[46][40] , \SUMB[46][39] , \SUMB[46][38] ,
         \SUMB[46][37] , \SUMB[46][36] , \SUMB[46][35] , \SUMB[46][34] ,
         \SUMB[46][33] , \SUMB[46][32] , \SUMB[46][31] , \SUMB[46][30] ,
         \SUMB[46][29] , \SUMB[46][28] , \SUMB[46][27] , \SUMB[46][26] ,
         \SUMB[46][25] , \SUMB[46][24] , \SUMB[46][23] , \SUMB[46][22] ,
         \SUMB[46][21] , \SUMB[46][20] , \SUMB[46][19] , \SUMB[46][18] ,
         \SUMB[46][17] , \SUMB[46][16] , \SUMB[46][15] , \SUMB[46][14] ,
         \SUMB[46][13] , \SUMB[46][12] , \SUMB[46][11] , \SUMB[46][10] ,
         \SUMB[46][9] , \SUMB[46][8] , \SUMB[46][7] , \SUMB[46][6] ,
         \SUMB[46][5] , \SUMB[46][4] , \SUMB[46][3] , \SUMB[46][2] ,
         \SUMB[46][1] , \SUMB[45][46] , \SUMB[45][45] , \SUMB[45][44] ,
         \SUMB[45][43] , \SUMB[45][42] , \SUMB[45][41] , \SUMB[45][40] ,
         \SUMB[45][39] , \SUMB[45][38] , \SUMB[45][37] , \SUMB[45][36] ,
         \SUMB[45][35] , \SUMB[45][34] , \SUMB[45][33] , \SUMB[45][32] ,
         \SUMB[45][31] , \SUMB[45][30] , \SUMB[45][29] , \SUMB[45][28] ,
         \SUMB[45][27] , \SUMB[45][26] , \SUMB[45][25] , \SUMB[45][24] ,
         \SUMB[45][23] , \SUMB[45][22] , \SUMB[45][21] , \SUMB[45][20] ,
         \SUMB[45][19] , \SUMB[45][18] , \SUMB[45][17] , \SUMB[45][16] ,
         \SUMB[45][15] , \SUMB[45][14] , \SUMB[45][13] , \SUMB[45][12] ,
         \SUMB[45][11] , \SUMB[45][10] , \SUMB[45][9] , \SUMB[45][8] ,
         \SUMB[45][7] , \SUMB[45][6] , \SUMB[45][5] , \SUMB[45][4] ,
         \SUMB[45][3] , \SUMB[45][2] , \SUMB[45][1] , \SUMB[44][46] ,
         \SUMB[44][45] , \SUMB[44][44] , \SUMB[44][43] , \SUMB[44][42] ,
         \SUMB[44][41] , \SUMB[44][40] , \SUMB[44][39] , \SUMB[44][38] ,
         \SUMB[44][37] , \SUMB[44][36] , \SUMB[44][35] , \SUMB[44][34] ,
         \SUMB[44][33] , \SUMB[44][32] , \SUMB[44][31] , \SUMB[44][30] ,
         \SUMB[44][29] , \SUMB[44][28] , \SUMB[44][27] , \SUMB[44][26] ,
         \SUMB[44][25] , \SUMB[44][24] , \SUMB[44][23] , \SUMB[44][22] ,
         \SUMB[44][21] , \SUMB[44][20] , \SUMB[44][19] , \SUMB[44][18] ,
         \SUMB[44][17] , \SUMB[44][16] , \SUMB[44][15] , \SUMB[44][14] ,
         \SUMB[44][13] , \SUMB[44][12] , \SUMB[44][11] , \SUMB[44][10] ,
         \SUMB[44][9] , \SUMB[44][8] , \SUMB[44][7] , \SUMB[44][6] ,
         \SUMB[44][5] , \SUMB[44][4] , \SUMB[44][3] , \SUMB[44][2] ,
         \SUMB[44][1] , \SUMB[43][46] , \SUMB[43][45] , \SUMB[43][44] ,
         \SUMB[43][43] , \SUMB[43][42] , \SUMB[43][41] , \SUMB[43][40] ,
         \SUMB[43][39] , \SUMB[43][38] , \SUMB[43][37] , \SUMB[43][36] ,
         \SUMB[43][35] , \SUMB[43][34] , \SUMB[43][33] , \SUMB[43][32] ,
         \SUMB[43][31] , \SUMB[43][30] , \SUMB[43][29] , \SUMB[43][28] ,
         \SUMB[43][27] , \SUMB[43][26] , \SUMB[43][25] , \SUMB[43][24] ,
         \SUMB[43][23] , \SUMB[43][22] , \SUMB[43][21] , \SUMB[43][20] ,
         \SUMB[43][19] , \SUMB[43][18] , \SUMB[43][17] , \SUMB[43][16] ,
         \SUMB[43][15] , \SUMB[43][14] , \SUMB[43][13] , \SUMB[43][12] ,
         \SUMB[43][11] , \SUMB[43][10] , \SUMB[43][9] , \SUMB[43][8] ,
         \SUMB[43][7] , \SUMB[43][6] , \SUMB[43][5] , \SUMB[43][4] ,
         \SUMB[43][3] , \SUMB[43][2] , \SUMB[43][1] , \SUMB[42][46] ,
         \SUMB[42][45] , \SUMB[42][44] , \SUMB[42][43] , \SUMB[42][42] ,
         \SUMB[42][41] , \SUMB[42][40] , \SUMB[42][39] , \SUMB[42][38] ,
         \SUMB[42][37] , \SUMB[42][36] , \SUMB[42][35] , \SUMB[42][34] ,
         \SUMB[42][33] , \SUMB[42][32] , \SUMB[42][31] , \SUMB[42][30] ,
         \SUMB[42][29] , \SUMB[42][28] , \SUMB[42][27] , \SUMB[42][26] ,
         \SUMB[42][25] , \SUMB[42][24] , \SUMB[42][23] , \SUMB[42][22] ,
         \SUMB[42][21] , \SUMB[42][20] , \SUMB[42][19] , \SUMB[42][18] ,
         \SUMB[42][17] , \SUMB[42][16] , \SUMB[42][15] , \SUMB[42][14] ,
         \SUMB[42][13] , \SUMB[42][12] , \SUMB[42][11] , \SUMB[42][10] ,
         \SUMB[42][9] , \SUMB[42][8] , \SUMB[42][7] , \SUMB[42][6] ,
         \SUMB[42][5] , \SUMB[42][4] , \SUMB[42][3] , \SUMB[42][2] ,
         \SUMB[42][1] , \SUMB[41][46] , \SUMB[41][45] , \SUMB[41][44] ,
         \SUMB[41][43] , \SUMB[41][42] , \SUMB[41][41] , \SUMB[41][40] ,
         \SUMB[41][39] , \SUMB[41][38] , \SUMB[41][37] , \SUMB[41][36] ,
         \SUMB[41][35] , \SUMB[41][34] , \SUMB[41][33] , \SUMB[41][32] ,
         \SUMB[41][31] , \SUMB[41][30] , \SUMB[41][29] , \SUMB[41][28] ,
         \SUMB[41][27] , \SUMB[41][26] , \SUMB[41][25] , \SUMB[41][24] ,
         \SUMB[41][23] , \SUMB[41][22] , \SUMB[41][21] , \SUMB[41][20] ,
         \SUMB[41][19] , \SUMB[41][18] , \SUMB[41][17] , \SUMB[41][16] ,
         \SUMB[41][15] , \SUMB[41][14] , \SUMB[41][13] , \SUMB[41][12] ,
         \SUMB[41][11] , \SUMB[41][10] , \SUMB[41][9] , \SUMB[41][8] ,
         \SUMB[41][7] , \SUMB[41][6] , \SUMB[41][5] , \SUMB[41][4] ,
         \SUMB[41][3] , \SUMB[41][2] , \SUMB[41][1] , \SUMB[40][46] ,
         \SUMB[40][45] , \SUMB[40][44] , \SUMB[40][43] , \SUMB[40][42] ,
         \SUMB[40][41] , \SUMB[40][40] , \SUMB[40][39] , \SUMB[40][38] ,
         \SUMB[40][37] , \SUMB[40][36] , \SUMB[40][35] , \SUMB[40][34] ,
         \SUMB[40][33] , \SUMB[40][32] , \SUMB[40][31] , \SUMB[40][30] ,
         \SUMB[40][29] , \SUMB[40][28] , \SUMB[40][27] , \SUMB[40][26] ,
         \SUMB[40][25] , \SUMB[40][24] , \SUMB[40][23] , \SUMB[40][22] ,
         \SUMB[40][21] , \SUMB[40][20] , \SUMB[40][19] , \SUMB[40][18] ,
         \SUMB[40][17] , \SUMB[40][16] , \SUMB[40][15] , \SUMB[40][14] ,
         \SUMB[40][13] , \SUMB[40][12] , \SUMB[40][11] , \SUMB[40][10] ,
         \SUMB[40][9] , \SUMB[40][8] , \SUMB[40][7] , \SUMB[40][6] ,
         \SUMB[40][5] , \SUMB[40][4] , \SUMB[40][3] , \SUMB[40][2] ,
         \SUMB[40][1] , \SUMB[39][46] , \SUMB[39][45] , \SUMB[39][44] ,
         \SUMB[39][43] , \SUMB[39][42] , \SUMB[39][41] , \SUMB[39][40] ,
         \SUMB[39][39] , \SUMB[39][38] , \SUMB[39][37] , \SUMB[39][36] ,
         \SUMB[39][35] , \SUMB[39][34] , \SUMB[39][33] , \SUMB[39][32] ,
         \SUMB[39][31] , \SUMB[39][30] , \SUMB[39][29] , \SUMB[39][28] ,
         \SUMB[39][27] , \SUMB[39][26] , \SUMB[39][25] , \SUMB[39][24] ,
         \SUMB[39][23] , \SUMB[39][22] , \SUMB[39][21] , \SUMB[39][20] ,
         \SUMB[39][19] , \SUMB[39][18] , \SUMB[39][17] , \SUMB[39][16] ,
         \SUMB[39][15] , \SUMB[39][14] , \SUMB[39][13] , \SUMB[39][12] ,
         \SUMB[39][11] , \SUMB[39][10] , \SUMB[39][9] , \SUMB[39][8] ,
         \SUMB[39][7] , \SUMB[39][6] , \SUMB[39][5] , \SUMB[39][4] ,
         \SUMB[39][3] , \SUMB[39][2] , \SUMB[39][1] , \SUMB[38][46] ,
         \SUMB[38][45] , \SUMB[38][44] , \SUMB[38][43] , \SUMB[38][42] ,
         \SUMB[38][41] , \SUMB[38][40] , \SUMB[38][39] , \SUMB[38][38] ,
         \SUMB[38][37] , \SUMB[38][36] , \SUMB[38][35] , \SUMB[38][34] ,
         \SUMB[38][33] , \SUMB[38][32] , \SUMB[38][31] , \SUMB[38][30] ,
         \SUMB[38][29] , \SUMB[38][28] , \SUMB[38][27] , \SUMB[38][26] ,
         \SUMB[38][25] , \SUMB[38][24] , \SUMB[38][23] , \SUMB[38][22] ,
         \SUMB[38][21] , \SUMB[38][20] , \SUMB[38][19] , \SUMB[38][18] ,
         \SUMB[38][17] , \SUMB[38][16] , \SUMB[38][15] , \SUMB[38][14] ,
         \SUMB[38][13] , \SUMB[38][12] , \SUMB[38][11] , \SUMB[38][10] ,
         \SUMB[38][9] , \SUMB[38][8] , \SUMB[38][7] , \SUMB[38][6] ,
         \SUMB[38][5] , \SUMB[38][4] , \SUMB[38][3] , \SUMB[38][2] ,
         \SUMB[38][1] , \SUMB[37][46] , \SUMB[37][45] , \SUMB[37][44] ,
         \SUMB[37][43] , \SUMB[37][42] , \SUMB[37][41] , \SUMB[37][40] ,
         \SUMB[37][39] , \SUMB[37][38] , \SUMB[37][37] , \SUMB[37][36] ,
         \SUMB[37][35] , \SUMB[37][34] , \SUMB[37][33] , \SUMB[37][32] ,
         \SUMB[37][31] , \SUMB[37][30] , \SUMB[37][29] , \SUMB[37][28] ,
         \SUMB[37][27] , \SUMB[37][26] , \SUMB[37][25] , \SUMB[37][24] ,
         \SUMB[37][23] , \SUMB[37][22] , \SUMB[37][21] , \SUMB[37][20] ,
         \SUMB[37][19] , \SUMB[37][18] , \SUMB[37][17] , \SUMB[37][16] ,
         \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] ,
         \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] ,
         \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] ,
         \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] ,
         \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] ,
         \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] ,
         \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[44] , \A1[43] ,
         \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] ,
         \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] ,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] ,
         \A2[87] , \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] ,
         \A2[80] , \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] ,
         \A2[73] , \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] ,
         \A2[66] , \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] ,
         \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] ,
         \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n651, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n736, n738, n739, n740,
         n741, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1395, n1396,
         n1397, n1398, n1399, n1400, n1403, n1404, n1405, n1408, n1409, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1422,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535;
  assign PRODUCT[0] = \B[0] ;
  assign \B[0]  = B[0];
  assign \ab[47][47]  = B[47];
  assign \ab[46][46]  = B[46];
  assign \ab[45][45]  = B[45];
  assign \ab[44][44]  = B[44];
  assign \ab[43][43]  = B[43];
  assign \ab[42][42]  = B[42];
  assign \ab[41][41]  = B[41];
  assign \ab[40][40]  = B[40];
  assign \ab[39][39]  = B[39];
  assign \ab[38][38]  = B[38];
  assign \ab[37][37]  = B[37];
  assign \ab[36][36]  = B[36];
  assign \ab[35][35]  = B[35];
  assign \ab[34][34]  = B[34];
  assign \ab[33][33]  = B[33];
  assign \ab[32][32]  = B[32];
  assign \ab[31][31]  = B[31];
  assign \ab[30][30]  = B[30];
  assign \ab[29][29]  = B[29];
  assign \ab[28][28]  = B[28];
  assign \ab[27][27]  = B[27];
  assign \ab[26][26]  = B[26];
  assign \ab[25][25]  = B[25];
  assign \ab[24][24]  = B[24];
  assign \ab[23][23]  = B[23];
  assign \ab[22][22]  = B[22];
  assign \ab[21][21]  = B[21];
  assign \ab[20][20]  = B[20];
  assign \ab[19][19]  = B[19];
  assign \ab[18][18]  = B[18];
  assign \ab[17][17]  = B[17];
  assign \ab[16][16]  = B[16];
  assign \ab[15][15]  = B[15];
  assign \ab[14][14]  = B[14];
  assign \ab[13][13]  = B[13];
  assign \ab[12][12]  = B[12];
  assign \ab[11][11]  = B[11];
  assign \ab[10][10]  = B[10];
  assign \ab[9][9]  = B[9];
  assign \ab[8][8]  = B[8];
  assign \ab[7][7]  = B[7];
  assign \ab[6][6]  = B[6];
  assign \ab[5][5]  = B[5];
  assign \ab[4][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[1][1]  = B[1];

  FA1AP S4_37 ( .A(\ab[47][37] ), .B(\CARRYB[46][37] ), .CI(\SUMB[46][38] ), 
        .CO(\CARRYB[47][37] ), .S(\SUMB[47][37] ) );
  FA1AP S2_45_15 ( .A(\ab[45][15] ), .B(\CARRYB[44][15] ), .CI(\SUMB[44][16] ), 
        .CO(\CARRYB[45][15] ), .S(\SUMB[45][15] ) );
  FA1AP S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA1AP S2_7_36 ( .A(n470), .B(\CARRYB[6][36] ), .CI(\SUMB[6][37] ), .CO(
        \CARRYB[7][36] ), .S(\SUMB[7][36] ) );
  FA1AP S2_3_16 ( .A(n1321), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), .CO(
        \CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1AP S2_2_38 ( .A(n1312), .B(\CARRYB[1][38] ), .CI(\SUMB[1][39] ), .CO(
        \CARRYB[2][38] ), .S(\SUMB[2][38] ) );
  LOG_POLY_DW01_add_5 FS_1 ( .A({1'b0, \A1[92] , \A1[91] , \A1[90] , \A1[89] , 
        \A1[88] , \A1[87] , \A1[86] , \A1[85] , \A1[84] , \A1[83] , \A1[82] , 
        \A1[81] , \A1[80] , \A1[79] , \A1[78] , \A1[77] , \A1[76] , \A1[75] , 
        \A1[74] , \A1[73] , \A1[72] , \A1[71] , \A1[70] , \A1[69] , \A1[68] , 
        \A1[67] , \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] , \A1[61] , 
        \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , 
        \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , 
        \A1[46] , \SUMB[47][0] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , 
        \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[93] , 
        \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] , \A2[86] , 
        \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] , \A2[79] , 
        \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] , \A2[72] , 
        \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] , \A2[65] , 
        \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , 
        \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , 
        \A2[50] , \A2[49] , \A2[48] , \A2[47] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[95:2])
         );
  FA1P S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA1P S2_41_10 ( .A(\ab[41][10] ), .B(\CARRYB[40][10] ), .CI(\SUMB[40][11] ), 
        .CO(\CARRYB[41][10] ), .S(\SUMB[41][10] ) );
  FA1A S2_9_1 ( .A(n1378), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1P S2_41_8 ( .A(n519), .B(\CARRYB[40][8] ), .CI(\SUMB[40][9] ), .CO(
        \CARRYB[41][8] ), .S(\SUMB[41][8] ) );
  FA1 S2_8_28 ( .A(\CARRYB[7][28] ), .B(n277), .CI(\SUMB[7][29] ), .CO(
        \CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA1P S2_39_4 ( .A(n355), .B(\CARRYB[38][4] ), .CI(\SUMB[38][5] ), .CO(
        \CARRYB[39][4] ), .S(\SUMB[39][4] ) );
  FA1P S2_40_22 ( .A(\ab[40][22] ), .B(\CARRYB[39][22] ), .CI(\SUMB[39][23] ), 
        .CO(\CARRYB[40][22] ), .S(\SUMB[40][22] ) );
  FA1P S2_11_32 ( .A(n577), .B(\CARRYB[10][32] ), .CI(\SUMB[10][33] ), .CO(
        \CARRYB[11][32] ), .S(\SUMB[11][32] ) );
  FA1P S2_12_25 ( .A(\CARRYB[11][25] ), .B(n610), .CI(\SUMB[11][26] ), .CO(
        \CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA1P S2_42_15 ( .A(\ab[42][15] ), .B(\CARRYB[41][15] ), .CI(\SUMB[41][16] ), 
        .CO(\CARRYB[42][15] ), .S(\SUMB[42][15] ) );
  FA1P S2_26_30 ( .A(\ab[30][26] ), .B(\CARRYB[25][30] ), .CI(\SUMB[25][31] ), 
        .CO(\CARRYB[26][30] ), .S(\SUMB[26][30] ) );
  FA1P S2_18_14 ( .A(n644), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), .CO(
        \CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA1P S2_19_14 ( .A(n636), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), .CO(
        \CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA1P S2_28_14 ( .A(\CARRYB[27][14] ), .B(\ab[28][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA1A S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA1P S2_15_40 ( .A(\ab[40][15] ), .B(\CARRYB[14][40] ), .CI(\SUMB[14][41] ), 
        .CO(\CARRYB[15][40] ), .S(\SUMB[15][40] ) );
  FA1P S2_15_41 ( .A(\ab[41][15] ), .B(\CARRYB[14][41] ), .CI(\SUMB[14][42] ), 
        .CO(\CARRYB[15][41] ), .S(\SUMB[15][41] ) );
  FA1P S2_16_40 ( .A(\ab[40][16] ), .B(\CARRYB[15][40] ), .CI(\SUMB[15][41] ), 
        .CO(\CARRYB[16][40] ), .S(\SUMB[16][40] ) );
  FA1P S2_37_6 ( .A(n1286), .B(\CARRYB[36][6] ), .CI(\SUMB[36][7] ), .CO(
        \CARRYB[37][6] ), .S(\SUMB[37][6] ) );
  FA1P S2_35_6 ( .A(n409), .B(\CARRYB[34][6] ), .CI(\SUMB[34][7] ), .CO(
        \CARRYB[35][6] ), .S(\SUMB[35][6] ) );
  FA1P S2_36_6 ( .A(n436), .B(\CARRYB[35][6] ), .CI(\SUMB[35][7] ), .CO(
        \CARRYB[36][6] ), .S(\SUMB[36][6] ) );
  FA1P S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA1A S2_8_1 ( .A(n1353), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_8_2 ( .A(n340), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S1_10_0 ( .A(n1385), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1P S2_9_26 ( .A(\SUMB[8][27] ), .B(n523), .CI(\CARRYB[8][26] ), .CO(
        \CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA1P S2_23_26 ( .A(\CARRYB[22][26] ), .B(\ab[26][23] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA1P S4_12 ( .A(\ab[47][12] ), .B(\CARRYB[46][12] ), .CI(\SUMB[46][13] ), 
        .CO(\CARRYB[47][12] ), .S(\SUMB[47][12] ) );
  FA1P S2_30_12 ( .A(n598), .B(\CARRYB[29][12] ), .CI(\SUMB[29][13] ), .CO(
        \CARRYB[30][12] ), .S(\SUMB[30][12] ) );
  FA1P S2_40_8 ( .A(n454), .B(\CARRYB[39][8] ), .CI(\SUMB[39][9] ), .CO(
        \CARRYB[40][8] ), .S(\SUMB[40][8] ) );
  FA1P S2_20_10 ( .A(n549), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), .CO(
        \CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA1P S2_6_31 ( .A(n453), .B(\CARRYB[5][31] ), .CI(\SUMB[5][32] ), .CO(
        \CARRYB[6][31] ), .S(\SUMB[6][31] ) );
  FA1P S2_36_17 ( .A(\ab[36][17] ), .B(\CARRYB[35][17] ), .CI(\SUMB[35][18] ), 
        .CO(\CARRYB[36][17] ), .S(\SUMB[36][17] ) );
  FA1P S2_37_17 ( .A(\ab[37][17] ), .B(\CARRYB[36][17] ), .CI(\SUMB[36][18] ), 
        .CO(\CARRYB[37][17] ), .S(\SUMB[37][17] ) );
  FA1P S2_39_3 ( .A(n269), .B(\CARRYB[38][3] ), .CI(\SUMB[38][4] ), .CO(
        \CARRYB[39][3] ), .S(\SUMB[39][3] ) );
  FA1P S2_40_3 ( .A(n288), .B(\CARRYB[39][3] ), .CI(\SUMB[39][4] ), .CO(
        \CARRYB[40][3] ), .S(\SUMB[40][3] ) );
  FA1P S2_14_41 ( .A(\ab[41][14] ), .B(\CARRYB[13][41] ), .CI(\SUMB[13][42] ), 
        .CO(\CARRYB[14][41] ), .S(\SUMB[14][41] ) );
  FA1P S2_13_41 ( .A(\ab[41][13] ), .B(\CARRYB[12][41] ), .CI(\SUMB[12][42] ), 
        .CO(\CARRYB[13][41] ), .S(\SUMB[13][41] ) );
  FA1A S2_34_44 ( .A(\ab[44][34] ), .B(\CARRYB[33][44] ), .CI(\SUMB[33][45] ), 
        .CO(\CARRYB[34][44] ), .S(\SUMB[34][44] ) );
  FA1P S2_10_43 ( .A(\ab[43][10] ), .B(\CARRYB[9][43] ), .CI(\SUMB[9][44] ), 
        .CO(\CARRYB[10][43] ), .S(\SUMB[10][43] ) );
  FA1P S2_38_5 ( .A(n1273), .B(\CARRYB[37][5] ), .CI(\SUMB[37][6] ), .CO(
        \CARRYB[38][5] ), .S(\SUMB[38][5] ) );
  FA1P S2_39_5 ( .A(n384), .B(\CARRYB[38][5] ), .CI(\SUMB[38][6] ), .CO(
        \CARRYB[39][5] ), .S(\SUMB[39][5] ) );
  FA1P S2_11_20 ( .A(n1322), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), .CO(
        \CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1P S2_29_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA1P S2_27_30 ( .A(\CARRYB[26][30] ), .B(\ab[30][27] ), .CI(\SUMB[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA1P S2_17_33 ( .A(\ab[33][17] ), .B(\CARRYB[16][33] ), .CI(\SUMB[16][34] ), 
        .CO(\CARRYB[17][33] ), .S(\SUMB[17][33] ) );
  FA1P S2_16_33 ( .A(\ab[33][16] ), .B(\CARRYB[15][33] ), .CI(\SUMB[15][34] ), 
        .CO(\CARRYB[16][33] ), .S(\SUMB[16][33] ) );
  FA1P S2_38_9 ( .A(n522), .B(\CARRYB[37][9] ), .CI(\SUMB[37][10] ), .CO(
        \CARRYB[38][9] ), .S(\SUMB[38][9] ) );
  FA1P S2_31_7 ( .A(n460), .B(\CARRYB[30][7] ), .CI(\SUMB[30][8] ), .CO(
        \CARRYB[31][7] ), .S(\SUMB[31][7] ) );
  FA1P S2_40_5 ( .A(n377), .B(\CARRYB[39][5] ), .CI(\SUMB[39][6] ), .CO(
        \CARRYB[40][5] ), .S(\SUMB[40][5] ) );
  FA1P S2_11_15 ( .A(n585), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), .CO(
        \CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1P S2_41_15 ( .A(\ab[41][15] ), .B(\CARRYB[40][15] ), .CI(\SUMB[40][16] ), 
        .CO(\CARRYB[41][15] ), .S(\SUMB[41][15] ) );
  FA1P S2_12_37 ( .A(\CARRYB[11][37] ), .B(\ab[37][12] ), .CI(\SUMB[11][38] ), 
        .CO(\CARRYB[12][37] ), .S(\SUMB[12][37] ) );
  FA1P S2_14_43 ( .A(\ab[43][14] ), .B(\CARRYB[13][43] ), .CI(\SUMB[13][44] ), 
        .CO(\CARRYB[14][43] ), .S(\SUMB[14][43] ) );
  FA1P S2_32_9 ( .A(n501), .B(\CARRYB[31][9] ), .CI(\SUMB[31][10] ), .CO(
        \CARRYB[32][9] ), .S(\SUMB[32][9] ) );
  FA1P S2_7_24 ( .A(n1285), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), .CO(
        \CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA1P S2_30_23 ( .A(\ab[30][23] ), .B(\CARRYB[29][23] ), .CI(\SUMB[29][24] ), 
        .CO(\CARRYB[30][23] ), .S(\SUMB[30][23] ) );
  FA1P S2_31_23 ( .A(\ab[31][23] ), .B(\CARRYB[30][23] ), .CI(\SUMB[30][24] ), 
        .CO(\CARRYB[31][23] ), .S(\SUMB[31][23] ) );
  FA1P S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA1P S2_19_10 ( .A(n560), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), .CO(
        \CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA1P S2_30_25 ( .A(\ab[30][25] ), .B(\CARRYB[29][25] ), .CI(\SUMB[29][26] ), 
        .CO(\CARRYB[30][25] ), .S(\SUMB[30][25] ) );
  FA1P S2_31_25 ( .A(\ab[31][25] ), .B(\CARRYB[30][25] ), .CI(\SUMB[30][26] ), 
        .CO(\CARRYB[31][25] ), .S(\SUMB[31][25] ) );
  FA1P S2_14_29 ( .A(\ab[29][14] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA1P S2_11_36 ( .A(\CARRYB[10][36] ), .B(\ab[36][11] ), .CI(\SUMB[10][37] ), 
        .CO(\CARRYB[11][36] ), .S(\SUMB[11][36] ) );
  FA1P S2_39_16 ( .A(\ab[39][16] ), .B(\CARRYB[38][16] ), .CI(\SUMB[38][17] ), 
        .CO(\CARRYB[39][16] ), .S(\SUMB[39][16] ) );
  FA1P S2_38_16 ( .A(\ab[38][16] ), .B(\CARRYB[37][16] ), .CI(\SUMB[37][17] ), 
        .CO(\CARRYB[38][16] ), .S(\SUMB[38][16] ) );
  FA1P S2_14_17 ( .A(n643), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), .CO(
        \CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA1P S2_6_22 ( .A(n408), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), .CO(
        \CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA1P S2_37_5 ( .A(n1281), .B(\CARRYB[36][5] ), .CI(\SUMB[36][6] ), .CO(
        \CARRYB[37][5] ), .S(\SUMB[37][5] ) );
  FA1P S2_38_6 ( .A(n1280), .B(\CARRYB[37][6] ), .CI(\SUMB[37][7] ), .CO(
        \CARRYB[38][6] ), .S(\SUMB[38][6] ) );
  FA1P S2_37_10 ( .A(n567), .B(\CARRYB[36][10] ), .CI(\SUMB[36][11] ), .CO(
        \CARRYB[37][10] ), .S(\SUMB[37][10] ) );
  FA1P S2_13_19 ( .A(n630), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), .CO(
        \CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA1P S2_36_10 ( .A(n574), .B(\CARRYB[35][10] ), .CI(\SUMB[35][11] ), .CO(
        \CARRYB[36][10] ), .S(\SUMB[36][10] ) );
  FA1P S4_2 ( .A(n271), .B(\CARRYB[46][2] ), .CI(\SUMB[46][3] ), .CO(
        \CARRYB[47][2] ), .S(\SUMB[47][2] ) );
  FA1P S2_40_15 ( .A(\ab[40][15] ), .B(\CARRYB[39][15] ), .CI(\SUMB[39][16] ), 
        .CO(\CARRYB[40][15] ), .S(\SUMB[40][15] ) );
  FA1P S2_39_15 ( .A(\ab[39][15] ), .B(\CARRYB[38][15] ), .CI(\SUMB[38][16] ), 
        .CO(\CARRYB[39][15] ), .S(\SUMB[39][15] ) );
  FA1P S2_37_27 ( .A(\ab[37][27] ), .B(\CARRYB[36][27] ), .CI(\SUMB[36][28] ), 
        .CO(\CARRYB[37][27] ), .S(\SUMB[37][27] ) );
  FA1P S2_29_27 ( .A(\ab[29][27] ), .B(\CARRYB[28][27] ), .CI(\SUMB[28][28] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA1P S2_27_27 ( .A(n1483), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), .CO(
        \CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA1P S2_9_16 ( .A(n535), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), .CO(
        \CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1P S2_29_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA1P S2_17_27 ( .A(\ab[27][17] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA1P S2_9_36 ( .A(n537), .B(\CARRYB[8][36] ), .CI(\SUMB[8][37] ), .CO(
        \CARRYB[9][36] ), .S(\SUMB[9][36] ) );
  FA1P S2_4_32 ( .A(n376), .B(\CARRYB[3][32] ), .CI(\SUMB[3][33] ), .CO(
        \CARRYB[4][32] ), .S(\SUMB[4][32] ) );
  FA1P S2_5_32 ( .A(n390), .B(\CARRYB[4][32] ), .CI(\SUMB[4][33] ), .CO(
        \CARRYB[5][32] ), .S(\SUMB[5][32] ) );
  FA1P S2_14_32 ( .A(\ab[32][14] ), .B(\CARRYB[13][32] ), .CI(\SUMB[13][33] ), 
        .CO(\CARRYB[14][32] ), .S(\SUMB[14][32] ) );
  FA1P S2_15_32 ( .A(\ab[32][15] ), .B(\CARRYB[14][32] ), .CI(\SUMB[14][33] ), 
        .CO(\CARRYB[15][32] ), .S(\SUMB[15][32] ) );
  FA1P S2_15_18 ( .A(\ab[18][15] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA1P S2_33_8 ( .A(n489), .B(\CARRYB[32][8] ), .CI(\SUMB[32][9] ), .CO(
        \CARRYB[33][8] ), .S(\SUMB[33][8] ) );
  FA1P S2_34_8 ( .A(n488), .B(\CARRYB[33][8] ), .CI(\SUMB[33][9] ), .CO(
        \CARRYB[34][8] ), .S(\SUMB[34][8] ) );
  FA1P S2_28_10 ( .A(n548), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), .CO(
        \CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA1P S2_43_32 ( .A(\ab[43][32] ), .B(\CARRYB[42][32] ), .CI(\SUMB[42][33] ), 
        .CO(\CARRYB[43][32] ), .S(\SUMB[43][32] ) );
  FA1P S2_15_43 ( .A(\ab[43][15] ), .B(\CARRYB[14][43] ), .CI(\SUMB[14][44] ), 
        .CO(\CARRYB[15][43] ), .S(\SUMB[15][43] ) );
  FA1P S2_12_29 ( .A(\CARRYB[11][29] ), .B(n609), .CI(\SUMB[11][30] ), .CO(
        \CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA1P S2_39_23 ( .A(\ab[39][23] ), .B(\CARRYB[38][23] ), .CI(\SUMB[38][24] ), 
        .CO(\CARRYB[39][23] ), .S(\SUMB[39][23] ) );
  FA1P S2_33_6 ( .A(n434), .B(\CARRYB[32][6] ), .CI(\SUMB[32][7] ), .CO(
        \CARRYB[33][6] ), .S(\SUMB[33][6] ) );
  FA1P S2_34_6 ( .A(n430), .B(\CARRYB[33][6] ), .CI(\SUMB[33][7] ), .CO(
        \CARRYB[34][6] ), .S(\SUMB[34][6] ) );
  FA1P S4_5 ( .A(n274), .B(\CARRYB[46][5] ), .CI(\SUMB[46][6] ), .CO(
        \CARRYB[47][5] ), .S(\SUMB[47][5] ) );
  FA1P S2_11_42 ( .A(\ab[42][11] ), .B(\CARRYB[10][42] ), .CI(\SUMB[10][43] ), 
        .CO(\CARRYB[11][42] ), .S(\SUMB[11][42] ) );
  FA1P S2_12_42 ( .A(\ab[42][12] ), .B(\CARRYB[11][42] ), .CI(\SUMB[11][43] ), 
        .CO(\CARRYB[12][42] ), .S(\SUMB[12][42] ) );
  FA1P S2_9_43 ( .A(\ab[9][43] ), .B(\CARRYB[8][43] ), .CI(\SUMB[8][44] ), 
        .CO(\CARRYB[9][43] ), .S(\SUMB[9][43] ) );
  FA1P S2_10_42 ( .A(\ab[42][10] ), .B(\CARRYB[9][42] ), .CI(\SUMB[9][43] ), 
        .CO(\CARRYB[10][42] ), .S(\SUMB[10][42] ) );
  FA1P S2_44_25 ( .A(\ab[44][25] ), .B(\CARRYB[43][25] ), .CI(\SUMB[43][26] ), 
        .CO(\CARRYB[44][25] ), .S(\SUMB[44][25] ) );
  FA1P S2_46_12 ( .A(\ab[46][12] ), .B(\CARRYB[45][12] ), .CI(\SUMB[45][13] ), 
        .CO(\CARRYB[46][12] ), .S(\SUMB[46][12] ) );
  FA1P S2_9_21 ( .A(n512), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), .CO(
        \CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA1A S4_32 ( .A(\ab[47][32] ), .B(\CARRYB[46][32] ), .CI(\SUMB[46][33] ), 
        .CO(\CARRYB[47][32] ), .S(\SUMB[47][32] ) );
  FA1P S1_45_0 ( .A(n1416), .B(\CARRYB[44][0] ), .CI(\SUMB[44][1] ), .CO(
        \CARRYB[45][0] ), .S(\A1[43] ) );
  FA1A S2_7_1 ( .A(n1381), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1P S2_20_26 ( .A(\ab[26][20] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA1P S2_38_23 ( .A(\ab[38][23] ), .B(\CARRYB[37][23] ), .CI(\SUMB[37][24] ), 
        .CO(\CARRYB[38][23] ), .S(\SUMB[38][23] ) );
  FA1P S2_6_44 ( .A(n273), .B(\CARRYB[5][44] ), .CI(\SUMB[5][45] ), .CO(
        \CARRYB[6][44] ), .S(\SUMB[6][44] ) );
  FA1P S2_7_44 ( .A(n467), .B(\CARRYB[6][44] ), .CI(\SUMB[6][45] ), .CO(
        \CARRYB[7][44] ), .S(\SUMB[7][44] ) );
  FA1P S2_13_43 ( .A(\ab[43][13] ), .B(\CARRYB[12][43] ), .CI(\SUMB[12][44] ), 
        .CO(\CARRYB[13][43] ), .S(\SUMB[13][43] ) );
  FA1P S2_12_41 ( .A(\ab[41][12] ), .B(\CARRYB[11][41] ), .CI(\SUMB[11][42] ), 
        .CO(\CARRYB[12][41] ), .S(\SUMB[12][41] ) );
  FA1P S2_12_44 ( .A(\ab[44][12] ), .B(\CARRYB[11][44] ), .CI(\SUMB[11][45] ), 
        .CO(\CARRYB[12][44] ), .S(\SUMB[12][44] ) );
  FA1P S2_13_44 ( .A(\ab[44][13] ), .B(\CARRYB[12][44] ), .CI(\SUMB[12][45] ), 
        .CO(\CARRYB[13][44] ), .S(\SUMB[13][44] ) );
  FA1P S2_36_5 ( .A(n407), .B(\CARRYB[35][5] ), .CI(\SUMB[35][6] ), .CO(
        \CARRYB[36][5] ), .S(\SUMB[36][5] ) );
  FA1P S2_11_37 ( .A(\ab[37][11] ), .B(\CARRYB[10][37] ), .CI(\SUMB[10][38] ), 
        .CO(\CARRYB[11][37] ), .S(\SUMB[11][37] ) );
  FA1P S2_20_21 ( .A(\ab[21][20] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA1P S2_21_21 ( .A(A[21]), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), .CO(
        \CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA1P S2_38_19 ( .A(\ab[38][19] ), .B(\CARRYB[37][19] ), .CI(\SUMB[37][20] ), 
        .CO(\CARRYB[38][19] ), .S(\SUMB[38][19] ) );
  FA1P S2_5_25 ( .A(n406), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), .CO(
        \CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA1P S2_6_25 ( .A(n405), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), .CO(
        \CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA1P S2_23_29 ( .A(\ab[29][23] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA1P S2_17_39 ( .A(\ab[39][17] ), .B(\CARRYB[16][39] ), .CI(\SUMB[16][40] ), 
        .CO(\CARRYB[17][39] ), .S(\SUMB[17][39] ) );
  FA1A S2_16_3 ( .A(n1321), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), .CO(
        \CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1P S2_21_10 ( .A(n547), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), .CO(
        \CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1P S2_36_23 ( .A(\ab[36][23] ), .B(\CARRYB[35][23] ), .CI(\SUMB[35][24] ), 
        .CO(\CARRYB[36][23] ), .S(\SUMB[36][23] ) );
  FA1P S2_37_23 ( .A(\ab[37][23] ), .B(\CARRYB[36][23] ), .CI(\SUMB[36][24] ), 
        .CO(\CARRYB[37][23] ), .S(\SUMB[37][23] ) );
  FA1P S2_37_4 ( .A(n1274), .B(\CARRYB[36][4] ), .CI(\SUMB[36][5] ), .CO(
        \CARRYB[37][4] ), .S(\SUMB[37][4] ) );
  FA1P S2_5_26 ( .A(n389), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), .CO(
        \CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA1AP S2_7_34 ( .A(n477), .B(\CARRYB[6][34] ), .CI(\SUMB[6][35] ), .CO(
        \CARRYB[7][34] ), .S(\SUMB[7][34] ) );
  FA1P S2_8_43 ( .A(n511), .B(\CARRYB[7][43] ), .CI(\SUMB[7][44] ), .CO(
        \CARRYB[8][43] ), .S(\SUMB[8][43] ) );
  FA1P S2_20_14 ( .A(n637), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), .CO(
        \CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA1P S2_32_12 ( .A(n601), .B(\CARRYB[31][12] ), .CI(\SUMB[31][13] ), .CO(
        \CARRYB[32][12] ), .S(\SUMB[32][12] ) );
  FA1 S2_46_32 ( .A(\ab[46][32] ), .B(\CARRYB[45][32] ), .CI(\SUMB[45][33] ), 
        .CO(\CARRYB[46][32] ), .S(\SUMB[46][32] ) );
  FA1A S2_8_22 ( .A(\CARRYB[7][22] ), .B(n452), .CI(\SUMB[7][23] ), .CO(
        \CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA1P S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), 
        .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FA1P S2_31_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FA1P S2_17_42 ( .A(\ab[42][17] ), .B(\CARRYB[16][42] ), .CI(\SUMB[16][43] ), 
        .CO(\CARRYB[17][42] ), .S(\SUMB[17][42] ) );
  FA1 S2_43_41 ( .A(\ab[43][41] ), .B(\CARRYB[42][41] ), .CI(\SUMB[42][42] ), 
        .CO(\CARRYB[43][41] ), .S(\SUMB[43][41] ) );
  FA1A S2_44_41 ( .A(\ab[44][41] ), .B(\CARRYB[43][41] ), .CI(\SUMB[43][42] ), 
        .CO(\CARRYB[44][41] ), .S(\SUMB[44][41] ) );
  FA1P S2_19_19 ( .A(n1468), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), .CO(
        \CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA1P S2_42_4 ( .A(n322), .B(\CARRYB[41][4] ), .CI(\SUMB[41][5] ), .CO(
        \CARRYB[42][4] ), .S(\SUMB[42][4] ) );
  FA1P S2_43_4 ( .A(n337), .B(\CARRYB[42][4] ), .CI(\SUMB[42][5] ), .CO(
        \CARRYB[43][4] ), .S(\SUMB[43][4] ) );
  FA1P S2_36_20 ( .A(\ab[36][20] ), .B(\CARRYB[35][20] ), .CI(\SUMB[35][21] ), 
        .CO(\CARRYB[36][20] ), .S(\SUMB[36][20] ) );
  FA1P S2_3_26 ( .A(n336), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), .CO(
        \CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA1P S2_10_15 ( .A(n558), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), .CO(
        \CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1 S2_21_24 ( .A(\ab[24][21] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA1 S2_41_9 ( .A(\ab[9][41] ), .B(\CARRYB[40][9] ), .CI(\SUMB[40][10] ), 
        .CO(\CARRYB[41][9] ), .S(\SUMB[41][9] ) );
  FA1P S2_35_41 ( .A(\ab[41][35] ), .B(\CARRYB[34][41] ), .CI(\SUMB[34][42] ), 
        .CO(\CARRYB[35][41] ), .S(\SUMB[35][41] ) );
  FA1P S2_6_35 ( .A(n409), .B(\CARRYB[5][35] ), .CI(\SUMB[5][36] ), .CO(
        \CARRYB[6][35] ), .S(\SUMB[6][35] ) );
  FA1P S2_18_32 ( .A(\ab[32][18] ), .B(\CARRYB[17][32] ), .CI(\SUMB[17][33] ), 
        .CO(\CARRYB[18][32] ), .S(\SUMB[18][32] ) );
  FA1P S2_38_34 ( .A(\ab[38][34] ), .B(\CARRYB[37][34] ), .CI(\SUMB[37][35] ), 
        .CO(\CARRYB[38][34] ), .S(\SUMB[38][34] ) );
  FA1P S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA1P S2_38_4 ( .A(n335), .B(\CARRYB[37][4] ), .CI(\SUMB[37][5] ), .CO(
        \CARRYB[38][4] ), .S(\SUMB[38][4] ) );
  FA1P S2_11_33 ( .A(n573), .B(\CARRYB[10][33] ), .CI(\SUMB[10][34] ), .CO(
        \CARRYB[11][33] ), .S(\SUMB[11][33] ) );
  FA1P S2_3_39 ( .A(n269), .B(\CARRYB[2][39] ), .CI(\SUMB[2][40] ), .CO(
        \CARRYB[3][39] ), .S(\SUMB[3][39] ) );
  FA1P S2_13_42 ( .A(\ab[42][13] ), .B(\CARRYB[12][42] ), .CI(\SUMB[12][43] ), 
        .CO(\CARRYB[13][42] ), .S(\SUMB[13][42] ) );
  FA1P S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA1P S2_29_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA1 S2_45_36 ( .A(\ab[45][36] ), .B(\CARRYB[44][36] ), .CI(\SUMB[44][37] ), 
        .CO(\CARRYB[45][36] ), .S(\SUMB[45][36] ) );
  FA1P S2_36_34 ( .A(\ab[36][34] ), .B(\CARRYB[35][34] ), .CI(\SUMB[35][35] ), 
        .CO(\CARRYB[36][34] ), .S(\SUMB[36][34] ) );
  FA1P S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA1P S2_11_44 ( .A(\ab[44][11] ), .B(\CARRYB[10][44] ), .CI(\SUMB[10][45] ), 
        .CO(\CARRYB[11][44] ), .S(\SUMB[11][44] ) );
  FA1P S3_3_46 ( .A(n295), .B(\CARRYB[2][46] ), .CI(n271), .CO(\CARRYB[3][46] ), .S(\SUMB[3][46] ) );
  FA1 S2_22_11 ( .A(n565), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), .CO(
        \CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA1P S2_41_7 ( .A(n463), .B(\CARRYB[40][7] ), .CI(\SUMB[40][8] ), .CO(
        \CARRYB[41][7] ), .S(\SUMB[41][7] ) );
  FA1P S2_6_17 ( .A(n1292), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), .CO(
        \CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1P S2_7_17 ( .A(n448), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), .CO(
        \CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1P S2_35_5 ( .A(n382), .B(\CARRYB[34][5] ), .CI(\SUMB[34][6] ), .CO(
        \CARRYB[35][5] ), .S(\SUMB[35][5] ) );
  FA1P S2_35_10 ( .A(n532), .B(\CARRYB[34][10] ), .CI(\SUMB[34][11] ), .CO(
        \CARRYB[35][10] ), .S(\SUMB[35][10] ) );
  FA1P S2_11_43 ( .A(\ab[43][11] ), .B(\CARRYB[10][43] ), .CI(\SUMB[10][44] ), 
        .CO(\CARRYB[11][43] ), .S(\SUMB[11][43] ) );
  FA1P S2_4_44 ( .A(n354), .B(\CARRYB[3][44] ), .CI(\SUMB[3][45] ), .CO(
        \CARRYB[4][44] ), .S(\SUMB[4][44] ) );
  FA1P S2_5_44 ( .A(n415), .B(\CARRYB[4][44] ), .CI(\SUMB[4][45] ), .CO(
        \CARRYB[5][44] ), .S(\SUMB[5][44] ) );
  FA1P S2_8_13 ( .A(n487), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), .CO(
        \CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1P S2_39_6 ( .A(n432), .B(\CARRYB[38][6] ), .CI(\SUMB[38][7] ), .CO(
        \CARRYB[39][6] ), .S(\SUMB[39][6] ) );
  FA1P S2_5_31 ( .A(n403), .B(\CARRYB[4][31] ), .CI(\SUMB[4][32] ), .CO(
        \CARRYB[5][31] ), .S(\SUMB[5][31] ) );
  FA1 S2_2_17 ( .A(n294), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), .CO(
        \CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_11_26 ( .A(\CARRYB[10][26] ), .B(n578), .CI(\SUMB[10][27] ), .CO(
        \CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA1P S2_43_6 ( .A(n447), .B(\CARRYB[42][6] ), .CI(\SUMB[42][7] ), .CO(
        \CARRYB[43][6] ), .S(\SUMB[43][6] ) );
  FA1P S2_42_5 ( .A(n402), .B(\CARRYB[41][5] ), .CI(\SUMB[41][6] ), .CO(
        \CARRYB[42][5] ), .S(\SUMB[42][5] ) );
  FA1P S1_46_0 ( .A(n1336), .B(\CARRYB[45][0] ), .CI(\SUMB[45][1] ), .CO(
        \CARRYB[46][0] ), .S(\A1[44] ) );
  FA1A S2_11_4 ( .A(n381), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(
        \CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1P S2_10_33 ( .A(n542), .B(\CARRYB[9][33] ), .CI(\SUMB[9][34] ), .CO(
        \CARRYB[10][33] ), .S(\SUMB[10][33] ) );
  FA1P S2_23_40 ( .A(\ab[40][23] ), .B(\CARRYB[22][40] ), .CI(\SUMB[22][41] ), 
        .CO(\CARRYB[23][40] ), .S(\SUMB[23][40] ) );
  FA1P S2_36_38 ( .A(\ab[38][36] ), .B(\CARRYB[35][38] ), .CI(\SUMB[35][39] ), 
        .CO(\CARRYB[36][38] ), .S(\SUMB[36][38] ) );
  FA1P S2_37_37 ( .A(n1505), .B(\CARRYB[36][37] ), .CI(\SUMB[36][38] ), .CO(
        \CARRYB[37][37] ), .S(\SUMB[37][37] ) );
  FA1P S2_22_27 ( .A(\CARRYB[21][27] ), .B(\ab[27][22] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA1P S2_32_2 ( .A(n1315), .B(\CARRYB[31][2] ), .CI(\SUMB[31][3] ), .CO(
        \CARRYB[32][2] ), .S(\SUMB[32][2] ) );
  FA1A S2_3_1 ( .A(n1529), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_4_1 ( .A(n1533), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S1_18_0 ( .A(n1428), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), .CO(
        \CARRYB[18][0] ), .S(\A1[16] ) );
  FA1A S2_44_40 ( .A(\ab[44][40] ), .B(\CARRYB[43][40] ), .CI(\SUMB[43][41] ), 
        .CO(\CARRYB[44][40] ), .S(\SUMB[44][40] ) );
  FA1P S2_40_9 ( .A(\ab[9][40] ), .B(\CARRYB[39][9] ), .CI(\SUMB[39][10] ), 
        .CO(\CARRYB[40][9] ), .S(\SUMB[40][9] ) );
  FA1P S2_30_17 ( .A(\ab[30][17] ), .B(\CARRYB[29][17] ), .CI(\SUMB[29][18] ), 
        .CO(\CARRYB[30][17] ), .S(\SUMB[30][17] ) );
  FA1A S2_25_41 ( .A(\ab[41][25] ), .B(\CARRYB[24][41] ), .CI(\SUMB[24][42] ), 
        .CO(\CARRYB[25][41] ), .S(\SUMB[25][41] ) );
  FA1P S2_8_37 ( .A(n486), .B(\CARRYB[7][37] ), .CI(\SUMB[7][38] ), .CO(
        \CARRYB[8][37] ), .S(\SUMB[8][37] ) );
  FA1P S2_4_27 ( .A(\CARRYB[3][27] ), .B(n356), .CI(\SUMB[3][28] ), .CO(
        \CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA1A S2_17_19 ( .A(\CARRYB[16][19] ), .B(\ab[19][17] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA1A S2_44_15 ( .A(\ab[44][15] ), .B(\CARRYB[43][15] ), .CI(\SUMB[43][16] ), 
        .CO(\CARRYB[44][15] ), .S(\SUMB[44][15] ) );
  FA1P S2_35_11 ( .A(\ab[35][11] ), .B(\CARRYB[34][11] ), .CI(\SUMB[34][12] ), 
        .CO(\CARRYB[35][11] ), .S(\SUMB[35][11] ) );
  FA1P S2_40_7 ( .A(n418), .B(\CARRYB[39][7] ), .CI(\SUMB[39][8] ), .CO(
        \CARRYB[40][7] ), .S(\SUMB[40][7] ) );
  FA1P S2_33_5 ( .A(n386), .B(\CARRYB[32][5] ), .CI(\SUMB[32][6] ), .CO(
        \CARRYB[33][5] ), .S(\SUMB[33][5] ) );
  FA1P S2_34_5 ( .A(n392), .B(\CARRYB[33][5] ), .CI(\SUMB[33][6] ), .CO(
        \CARRYB[34][5] ), .S(\SUMB[34][5] ) );
  FA1P S2_10_44 ( .A(\ab[44][10] ), .B(\CARRYB[9][44] ), .CI(\SUMB[9][45] ), 
        .CO(\CARRYB[10][44] ), .S(\SUMB[10][44] ) );
  FA1P S2_9_19 ( .A(n531), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), .CO(
        \CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1P S2_33_12 ( .A(\ab[33][12] ), .B(\CARRYB[32][12] ), .CI(\SUMB[32][13] ), 
        .CO(\CARRYB[33][12] ), .S(\SUMB[33][12] ) );
  FA1P S2_42_32 ( .A(\ab[42][32] ), .B(\CARRYB[41][32] ), .CI(\SUMB[41][33] ), 
        .CO(\CARRYB[42][32] ), .S(\SUMB[42][32] ) );
  FA1P S2_35_23 ( .A(\ab[35][23] ), .B(\CARRYB[34][23] ), .CI(\SUMB[34][24] ), 
        .CO(\CARRYB[35][23] ), .S(\SUMB[35][23] ) );
  FA1P S2_34_23 ( .A(\CARRYB[33][23] ), .B(\ab[34][23] ), .CI(\SUMB[33][24] ), 
        .CO(\CARRYB[34][23] ), .S(\SUMB[34][23] ) );
  FA1P S1_43_0 ( .A(n1418), .B(\CARRYB[42][0] ), .CI(\SUMB[42][1] ), .CO(
        \CARRYB[43][0] ), .S(\A1[41] ) );
  FA1P S2_42_30 ( .A(\ab[42][30] ), .B(\CARRYB[41][30] ), .CI(\SUMB[41][31] ), 
        .CO(\CARRYB[42][30] ), .S(\SUMB[42][30] ) );
  FA1P S2_40_33 ( .A(\ab[40][33] ), .B(\CARRYB[39][33] ), .CI(\SUMB[39][34] ), 
        .CO(\CARRYB[40][33] ), .S(\SUMB[40][33] ) );
  FA1P S2_15_16 ( .A(\ab[16][15] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA1P S2_26_40 ( .A(\ab[40][26] ), .B(\CARRYB[25][40] ), .CI(\SUMB[25][41] ), 
        .CO(\CARRYB[26][40] ), .S(\SUMB[26][40] ) );
  FA1P S2_18_41 ( .A(\ab[41][18] ), .B(\CARRYB[17][41] ), .CI(\SUMB[17][42] ), 
        .CO(\CARRYB[18][41] ), .S(\SUMB[18][41] ) );
  FA1P S2_3_32 ( .A(n321), .B(\CARRYB[2][32] ), .CI(\SUMB[2][33] ), .CO(
        \CARRYB[3][32] ), .S(\SUMB[3][32] ) );
  FA1P S2_12_43 ( .A(\ab[43][12] ), .B(\CARRYB[11][43] ), .CI(\SUMB[11][44] ), 
        .CO(\CARRYB[12][43] ), .S(\SUMB[12][43] ) );
  FA1P S2_4_26 ( .A(n364), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), .CO(
        \CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA1P S2_41_3 ( .A(n282), .B(\CARRYB[40][3] ), .CI(\SUMB[40][4] ), .CO(
        \CARRYB[41][3] ), .S(\SUMB[41][3] ) );
  FA1P S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA1P S2_14_21 ( .A(n639), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), .CO(
        \CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA1A S2_21_6 ( .A(n439), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), .CO(
        \CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA1 S2_9_13 ( .A(n530), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), .CO(
        \CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1P S2_28_8 ( .A(n277), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), .CO(
        \CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA1P S2_16_27 ( .A(\ab[27][16] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA1P S2_3_15 ( .A(n1318), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), .CO(
        \CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1P S2_36_15 ( .A(\ab[36][15] ), .B(\CARRYB[35][15] ), .CI(\SUMB[35][16] ), 
        .CO(\CARRYB[36][15] ), .S(\SUMB[36][15] ) );
  FA1P S2_19_11 ( .A(n572), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), .CO(
        \CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA1P S2_41_30 ( .A(\ab[41][30] ), .B(\CARRYB[40][30] ), .CI(\SUMB[40][31] ), 
        .CO(\CARRYB[41][30] ), .S(\SUMB[41][30] ) );
  FA1P S2_32_25 ( .A(\ab[32][25] ), .B(\CARRYB[31][25] ), .CI(\SUMB[31][26] ), 
        .CO(\CARRYB[32][25] ), .S(\SUMB[32][25] ) );
  FA1P S2_8_16 ( .A(n518), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), .CO(
        \CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1P S2_19_30 ( .A(\ab[30][19] ), .B(\CARRYB[18][30] ), .CI(\SUMB[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA1 S2_8_31 ( .A(n485), .B(\CARRYB[7][31] ), .CI(\SUMB[7][32] ), .CO(
        \CARRYB[8][31] ), .S(\SUMB[8][31] ) );
  FA1 S2_20_16 ( .A(\CARRYB[19][16] ), .B(\ab[20][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA1P S2_37_34 ( .A(\ab[37][34] ), .B(\CARRYB[36][34] ), .CI(\SUMB[36][35] ), 
        .CO(\CARRYB[37][34] ), .S(\SUMB[37][34] ) );
  FA1P S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA1P S2_19_39 ( .A(\ab[39][19] ), .B(\CARRYB[18][39] ), .CI(\SUMB[18][40] ), 
        .CO(\CARRYB[19][39] ), .S(\SUMB[19][39] ) );
  FA1A S2_17_30 ( .A(\ab[30][17] ), .B(\CARRYB[16][30] ), .CI(\SUMB[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA1P S2_43_12 ( .A(\ab[43][12] ), .B(\CARRYB[42][12] ), .CI(\SUMB[42][13] ), 
        .CO(\CARRYB[43][12] ), .S(\SUMB[43][12] ) );
  FA1P S2_39_33 ( .A(\ab[39][33] ), .B(\CARRYB[38][33] ), .CI(\SUMB[38][34] ), 
        .CO(\CARRYB[39][33] ), .S(\SUMB[39][33] ) );
  FA1P S2_20_39 ( .A(\ab[39][20] ), .B(\CARRYB[19][39] ), .CI(\SUMB[19][40] ), 
        .CO(\CARRYB[20][39] ), .S(\SUMB[20][39] ) );
  FA1P S2_22_28 ( .A(\ab[28][22] ), .B(\CARRYB[21][28] ), .CI(\SUMB[21][29] ), 
        .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FA1P S2_29_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA1A S2_30_24 ( .A(\ab[30][24] ), .B(\CARRYB[29][24] ), .CI(\SUMB[29][25] ), 
        .CO(\CARRYB[30][24] ), .S(\SUMB[30][24] ) );
  FA1P S2_16_16 ( .A(A[16]), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), .CO(
        \CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA1P S2_39_9 ( .A(n529), .B(\CARRYB[38][9] ), .CI(\SUMB[38][10] ), .CO(
        \CARRYB[39][9] ), .S(\SUMB[39][9] ) );
  FA1 S2_7_22 ( .A(n416), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), .CO(
        \CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA1P S2_18_42 ( .A(\ab[42][18] ), .B(\CARRYB[17][42] ), .CI(\SUMB[17][43] ), 
        .CO(\CARRYB[18][42] ), .S(\SUMB[18][42] ) );
  FA1P S2_19_42 ( .A(\ab[42][19] ), .B(\CARRYB[18][42] ), .CI(\SUMB[18][43] ), 
        .CO(\CARRYB[19][42] ), .S(\SUMB[19][42] ) );
  FA1P S2_13_17 ( .A(n629), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), .CO(
        \CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA1P S2_31_30 ( .A(\ab[31][30] ), .B(\CARRYB[30][30] ), .CI(\SUMB[30][31] ), 
        .CO(\CARRYB[31][30] ), .S(\SUMB[31][30] ) );
  FA1A S2_46_37 ( .A(\ab[46][37] ), .B(\CARRYB[45][37] ), .CI(\SUMB[45][38] ), 
        .CO(\CARRYB[46][37] ), .S(\SUMB[46][37] ) );
  FA1P S2_39_31 ( .A(\ab[39][31] ), .B(\CARRYB[38][31] ), .CI(\SUMB[38][32] ), 
        .CO(\CARRYB[39][31] ), .S(\SUMB[39][31] ) );
  FA1P S2_19_40 ( .A(\ab[40][19] ), .B(\CARRYB[18][40] ), .CI(\SUMB[18][41] ), 
        .CO(\CARRYB[19][40] ), .S(\SUMB[19][40] ) );
  FA1P S2_20_40 ( .A(\ab[40][20] ), .B(\CARRYB[19][40] ), .CI(\SUMB[19][41] ), 
        .CO(\CARRYB[20][40] ), .S(\SUMB[20][40] ) );
  FA1 S2_4_29 ( .A(\CARRYB[3][29] ), .B(n1271), .CI(\SUMB[3][30] ), .CO(
        \CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA1P S2_31_26 ( .A(\ab[31][26] ), .B(\CARRYB[30][26] ), .CI(\SUMB[30][27] ), 
        .CO(\CARRYB[31][26] ), .S(\SUMB[31][26] ) );
  FA1P S2_18_29 ( .A(\ab[29][18] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA1P S2_3_33 ( .A(n318), .B(\CARRYB[2][33] ), .CI(\SUMB[2][34] ), .CO(
        \CARRYB[3][33] ), .S(\SUMB[3][33] ) );
  FA1P S2_37_9 ( .A(n546), .B(\CARRYB[36][9] ), .CI(\SUMB[36][10] ), .CO(
        \CARRYB[37][9] ), .S(\SUMB[37][9] ) );
  FA1P S2_27_15 ( .A(\CARRYB[26][15] ), .B(\ab[27][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA1P S2_21_39 ( .A(\ab[39][21] ), .B(\CARRYB[20][39] ), .CI(\SUMB[20][40] ), 
        .CO(\CARRYB[21][39] ), .S(\SUMB[21][39] ) );
  FA1A S2_41_16 ( .A(\ab[41][16] ), .B(\CARRYB[40][16] ), .CI(\SUMB[40][17] ), 
        .CO(\CARRYB[41][16] ), .S(\SUMB[41][16] ) );
  FA1P S2_29_13 ( .A(n621), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), .CO(
        \CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA1P S2_15_17 ( .A(\ab[17][15] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA1P S2_29_36 ( .A(\ab[36][29] ), .B(\CARRYB[28][36] ), .CI(\SUMB[28][37] ), 
        .CO(\CARRYB[29][36] ), .S(\SUMB[29][36] ) );
  FA1 S2_12_20 ( .A(\SUMB[11][21] ), .B(\CARRYB[11][20] ), .CI(n597), .CO(
        \CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA1P S2_29_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA1P S2_17_32 ( .A(\ab[32][17] ), .B(\CARRYB[16][32] ), .CI(\SUMB[16][33] ), 
        .CO(\CARRYB[17][32] ), .S(\SUMB[17][32] ) );
  FA1 S2_3_38 ( .A(n343), .B(\CARRYB[2][38] ), .CI(\SUMB[2][39] ), .CO(
        \CARRYB[3][38] ), .S(\SUMB[3][38] ) );
  FA1A S2_32_13 ( .A(\ab[32][13] ), .B(\CARRYB[31][13] ), .CI(\SUMB[31][14] ), 
        .CO(\CARRYB[32][13] ), .S(\SUMB[32][13] ) );
  FA1 S2_31_13 ( .A(\ab[31][13] ), .B(\CARRYB[30][13] ), .CI(\SUMB[30][14] ), 
        .CO(\CARRYB[31][13] ), .S(\SUMB[31][13] ) );
  FA1 S2_8_35 ( .A(n276), .B(\CARRYB[7][35] ), .CI(\SUMB[7][36] ), .CO(
        \CARRYB[8][35] ), .S(\SUMB[8][35] ) );
  FA1P S2_8_36 ( .A(n517), .B(\CARRYB[7][36] ), .CI(\SUMB[7][37] ), .CO(
        \CARRYB[8][36] ), .S(\SUMB[8][36] ) );
  FA1P S2_18_10 ( .A(n557), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), .CO(
        \CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA1A S2_9_33 ( .A(n516), .B(\CARRYB[8][33] ), .CI(\SUMB[8][34] ), .CO(
        \CARRYB[9][33] ), .S(\SUMB[9][33] ) );
  FA1P S2_31_19 ( .A(\ab[31][19] ), .B(\CARRYB[30][19] ), .CI(\SUMB[30][20] ), 
        .CO(\CARRYB[31][19] ), .S(\SUMB[31][19] ) );
  FA1P S2_42_26 ( .A(\ab[42][26] ), .B(\CARRYB[41][26] ), .CI(\SUMB[41][27] ), 
        .CO(\CARRYB[42][26] ), .S(\SUMB[42][26] ) );
  FA1P S2_15_19 ( .A(\ab[19][15] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA1P S2_2_34 ( .A(n1307), .B(\CARRYB[1][34] ), .CI(\SUMB[1][35] ), .CO(
        \CARRYB[2][34] ), .S(\SUMB[2][34] ) );
  FA1A S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA1P S2_29_40 ( .A(\ab[40][29] ), .B(\CARRYB[28][40] ), .CI(\SUMB[28][41] ), 
        .CO(\CARRYB[29][40] ), .S(\SUMB[29][40] ) );
  FA1P S2_30_40 ( .A(\ab[40][30] ), .B(\CARRYB[29][40] ), .CI(\SUMB[29][41] ), 
        .CO(\CARRYB[30][40] ), .S(\SUMB[30][40] ) );
  FA1A S2_43_10 ( .A(\ab[43][10] ), .B(\CARRYB[42][10] ), .CI(\SUMB[42][11] ), 
        .CO(\CARRYB[43][10] ), .S(\SUMB[43][10] ) );
  FA1A S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA1A S2_5_9 ( .A(n427), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S1_20_0 ( .A(n1375), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), .CO(
        \CARRYB[20][0] ), .S(\A1[18] ) );
  FA1AP S2_2_31 ( .A(n1340), .B(\CARRYB[1][31] ), .CI(\SUMB[1][32] ), .CO(
        \CARRYB[2][31] ), .S(\SUMB[2][31] ) );
  FA1P S2_5_36 ( .A(n407), .B(\CARRYB[4][36] ), .CI(\SUMB[4][37] ), .CO(
        \CARRYB[5][36] ), .S(\SUMB[5][36] ) );
  FA1P S2_35_38 ( .A(\ab[38][35] ), .B(\CARRYB[34][38] ), .CI(\SUMB[34][39] ), 
        .CO(\CARRYB[35][38] ), .S(\SUMB[35][38] ) );
  FA1P S2_3_13 ( .A(n360), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), .CO(
        \CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1 S2_42_10 ( .A(\ab[42][10] ), .B(\CARRYB[41][10] ), .CI(\SUMB[41][11] ), 
        .CO(\CARRYB[42][10] ), .S(\SUMB[42][10] ) );
  FA1 S2_34_12 ( .A(\ab[34][12] ), .B(\CARRYB[33][12] ), .CI(\SUMB[33][13] ), 
        .CO(\CARRYB[34][12] ), .S(\SUMB[34][12] ) );
  FA1P S2_2_22 ( .A(\CARRYB[1][22] ), .B(n1301), .CI(\SUMB[1][23] ), .CO(
        \CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA1A S2_41_31 ( .A(\ab[41][31] ), .B(\CARRYB[40][31] ), .CI(\SUMB[40][32] ), 
        .CO(\CARRYB[41][31] ), .S(\SUMB[41][31] ) );
  FA1P S2_6_20 ( .A(\CARRYB[5][20] ), .B(n429), .CI(\SUMB[5][21] ), .CO(
        \CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1 S2_40_31 ( .A(\ab[40][31] ), .B(\CARRYB[39][31] ), .CI(\SUMB[39][32] ), 
        .CO(\CARRYB[40][31] ), .S(\SUMB[40][31] ) );
  FA1P S2_30_9 ( .A(n462), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), .CO(
        \CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA1A S4_20 ( .A(\ab[47][20] ), .B(\CARRYB[46][20] ), .CI(\SUMB[46][21] ), 
        .CO(\CARRYB[47][20] ), .S(\SUMB[47][20] ) );
  FA1P S2_45_20 ( .A(\ab[45][20] ), .B(\CARRYB[44][20] ), .CI(\SUMB[44][21] ), 
        .CO(\CARRYB[45][20] ), .S(\SUMB[45][20] ) );
  FA1P S2_31_11 ( .A(n579), .B(\CARRYB[30][11] ), .CI(\SUMB[30][12] ), .CO(
        \CARRYB[31][11] ), .S(\SUMB[31][11] ) );
  FA1A S2_27_40 ( .A(\ab[40][27] ), .B(\CARRYB[26][40] ), .CI(\SUMB[26][41] ), 
        .CO(\CARRYB[27][40] ), .S(\SUMB[27][40] ) );
  FA1A S2_2_1 ( .A(n1535), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S1_15_0 ( .A(n1432), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\A1[13] ) );
  FA1A S1_2_0 ( .A(n1390), .B(\ab[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_9_0 ( .A(n1368), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_8_0 ( .A(n1386), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S1_7_0 ( .A(n1392), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_5_0 ( .A(n1389), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S1_4_0 ( .A(n1388), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S2_12_1 ( .A(n1354), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), .CO(
        \CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S1_22_0 ( .A(n310), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), .CO(
        \CARRYB[22][0] ), .S(\A1[20] ) );
  FA1A S2_13_1 ( .A(n1370), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), .CO(
        \CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_21_1 ( .A(n268), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), .CO(
        \CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_15_1 ( .A(n267), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1A S2_2_4 ( .A(n370), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_2_7 ( .A(n348), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_5_1 ( .A(n1377), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S1_12_0 ( .A(n1384), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), .CO(
        \CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S2_10_1 ( .A(n1346), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S1_23_0 ( .A(n1338), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), .CO(
        \CARRYB[23][0] ), .S(\A1[21] ) );
  FA1A S2_28_1 ( .A(n1331), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), .CO(
        \CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA1A S2_27_1 ( .A(n1330), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), .CO(
        \CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA1A S1_14_0 ( .A(n1351), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(
        \CARRYB[14][0] ), .S(\A1[12] ) );
  FA1A S1_17_0 ( .A(n1429), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), .CO(
        \CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S2_2_10 ( .A(n303), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), .CO(
        \CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S2_36_18 ( .A(\CARRYB[35][18] ), .B(\ab[36][18] ), .CI(\SUMB[35][19] ), 
        .CO(\CARRYB[36][18] ), .S(\SUMB[36][18] ) );
  FA1A S2_3_3 ( .A(n1435), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_21_3 ( .A(n330), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), .CO(
        \CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1A S2_41_41 ( .A(A[41]), .B(\CARRYB[40][41] ), .CI(\SUMB[40][42] ), .CO(
        \CARRYB[41][41] ), .S(\SUMB[41][41] ) );
  FA1A S2_3_10 ( .A(n328), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), .CO(
        \CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_4_2 ( .A(n370), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_7_4 ( .A(n369), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_12_4 ( .A(n380), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), .CO(
        \CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_9_3 ( .A(n347), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_4_7 ( .A(n369), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_15_4 ( .A(n362), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1A S2_5_4 ( .A(n379), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_5_2 ( .A(n359), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_11_6 ( .A(n457), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(
        \CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_23_2 ( .A(n302), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), .CO(
        \CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA1A S2_13_5 ( .A(n421), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), .CO(
        \CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_4_3 ( .A(n358), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_14_4 ( .A(n366), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(
        \CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_22_2 ( .A(n1301), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), .CO(
        \CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA1A S2_6_7 ( .A(n480), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_13_6 ( .A(n450), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), .CO(
        \CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_12_6 ( .A(n476), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), .CO(
        \CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_6_11 ( .A(n457), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), .CO(
        \CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_7_2 ( .A(n348), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_17_3 ( .A(n333), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), .CO(
        \CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1A S2_33_45 ( .A(\ab[45][33] ), .B(\CARRYB[32][45] ), .CI(\SUMB[32][46] ), 
        .CO(\CARRYB[33][45] ), .S(\SUMB[33][45] ) );
  FA1A S2_17_8 ( .A(n500), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), .CO(
        \CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1A S2_37_43 ( .A(\ab[43][37] ), .B(\CARRYB[36][43] ), .CI(\SUMB[36][44] ), 
        .CO(\CARRYB[37][43] ), .S(\SUMB[37][43] ) );
  FA1A S2_42_39 ( .A(\ab[42][39] ), .B(\CARRYB[41][39] ), .CI(\SUMB[41][40] ), 
        .CO(\CARRYB[42][39] ), .S(\SUMB[42][39] ) );
  FA1A S3_43_46 ( .A(\ab[46][43] ), .B(\CARRYB[42][46] ), .CI(\ab[47][42] ), 
        .CO(\CARRYB[43][46] ), .S(\SUMB[43][46] ) );
  FA1A S2_24_45 ( .A(\ab[45][24] ), .B(\CARRYB[23][45] ), .CI(\SUMB[23][46] ), 
        .CO(\CARRYB[24][45] ), .S(\SUMB[24][45] ) );
  FA1AP S4_30 ( .A(\ab[47][30] ), .B(\CARRYB[46][30] ), .CI(\SUMB[46][31] ), 
        .CO(\CARRYB[47][30] ), .S(\SUMB[47][30] ) );
  FA1A S2_24_3 ( .A(n307), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), .CO(
        \CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA1A S2_26_3 ( .A(n336), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), .CO(
        \CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA1A S2_23_5 ( .A(n394), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), .CO(
        \CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA1A S2_11_7 ( .A(n494), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(
        \CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_36_45 ( .A(\ab[45][36] ), .B(\CARRYB[35][45] ), .CI(\SUMB[35][46] ), 
        .CO(\CARRYB[36][45] ), .S(\SUMB[36][45] ) );
  FA1A S2_34_45 ( .A(\ab[45][34] ), .B(\CARRYB[33][45] ), .CI(\SUMB[33][46] ), 
        .CO(\CARRYB[34][45] ), .S(\SUMB[34][45] ) );
  FA1A S2_43_42 ( .A(\ab[43][42] ), .B(\CARRYB[42][42] ), .CI(\SUMB[42][43] ), 
        .CO(\CARRYB[43][42] ), .S(\SUMB[43][42] ) );
  FA1A S2_38_41 ( .A(\ab[41][38] ), .B(\CARRYB[37][41] ), .CI(\SUMB[37][42] ), 
        .CO(\CARRYB[38][41] ), .S(\SUMB[38][41] ) );
  FA1A S2_21_35 ( .A(\ab[35][21] ), .B(\CARRYB[20][35] ), .CI(\SUMB[20][36] ), 
        .CO(\CARRYB[21][35] ), .S(\SUMB[21][35] ) );
  FA1A S2_29_43 ( .A(\ab[43][29] ), .B(\CARRYB[28][43] ), .CI(\SUMB[28][44] ), 
        .CO(\CARRYB[29][43] ), .S(\SUMB[29][43] ) );
  FA1A S2_39_40 ( .A(\ab[40][39] ), .B(\CARRYB[38][40] ), .CI(\SUMB[38][41] ), 
        .CO(\CARRYB[39][40] ), .S(\SUMB[39][40] ) );
  FA1A S2_45_27 ( .A(\ab[45][27] ), .B(\CARRYB[44][27] ), .CI(\SUMB[44][28] ), 
        .CO(\CARRYB[45][27] ), .S(\SUMB[45][27] ) );
  FA1A S2_40_24 ( .A(\ab[40][24] ), .B(\CARRYB[39][24] ), .CI(\SUMB[39][25] ), 
        .CO(\CARRYB[40][24] ), .S(\SUMB[40][24] ) );
  FA1A S2_37_41 ( .A(\ab[41][37] ), .B(\CARRYB[36][41] ), .CI(\SUMB[36][42] ), 
        .CO(\CARRYB[37][41] ), .S(\SUMB[37][41] ) );
  FA1A S2_32_44 ( .A(\ab[44][32] ), .B(\CARRYB[31][44] ), .CI(\SUMB[31][45] ), 
        .CO(\CARRYB[32][44] ), .S(\SUMB[32][44] ) );
  FA1AP S2_17_11 ( .A(n581), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), .CO(
        \CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA1A S2_25_45 ( .A(\ab[45][25] ), .B(\CARRYB[24][45] ), .CI(\SUMB[24][46] ), 
        .CO(\CARRYB[25][45] ), .S(\SUMB[25][45] ) );
  FA1A S2_36_42 ( .A(\ab[42][36] ), .B(\CARRYB[35][42] ), .CI(\SUMB[35][43] ), 
        .CO(\CARRYB[36][42] ), .S(\SUMB[36][42] ) );
  FA1A S2_13_30 ( .A(n614), .B(\CARRYB[12][30] ), .CI(\SUMB[12][31] ), .CO(
        \CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA1AP S4_22 ( .A(\CARRYB[46][22] ), .B(\ab[47][22] ), .CI(\SUMB[46][23] ), 
        .CO(\CARRYB[47][22] ), .S(\SUMB[47][22] ) );
  FA1A S2_36_41 ( .A(\ab[41][36] ), .B(\CARRYB[35][41] ), .CI(\SUMB[35][42] ), 
        .CO(\CARRYB[36][41] ), .S(\SUMB[36][41] ) );
  FA1A S2_35_43 ( .A(\ab[43][35] ), .B(\CARRYB[34][43] ), .CI(\SUMB[34][44] ), 
        .CO(\CARRYB[35][43] ), .S(\SUMB[35][43] ) );
  FA1A S2_35_31 ( .A(\ab[35][31] ), .B(\CARRYB[34][31] ), .CI(\SUMB[34][32] ), 
        .CO(\CARRYB[35][31] ), .S(\SUMB[35][31] ) );
  FA1A S3_34_46 ( .A(\ab[46][34] ), .B(\CARRYB[33][46] ), .CI(\ab[47][33] ), 
        .CO(\CARRYB[34][46] ), .S(\SUMB[34][46] ) );
  FA1A S3_32_46 ( .A(\ab[46][32] ), .B(\CARRYB[31][46] ), .CI(\ab[47][31] ), 
        .CO(\CARRYB[32][46] ), .S(\SUMB[32][46] ) );
  FA1A S3_21_46 ( .A(\ab[46][21] ), .B(\CARRYB[20][46] ), .CI(\ab[47][20] ), 
        .CO(\CARRYB[21][46] ), .S(\SUMB[21][46] ) );
  FA1AP S4_15 ( .A(\ab[47][15] ), .B(\CARRYB[46][15] ), .CI(\SUMB[46][16] ), 
        .CO(\CARRYB[47][15] ), .S(\SUMB[47][15] ) );
  FA1AP S4_10 ( .A(\CARRYB[46][10] ), .B(\ab[47][10] ), .CI(\SUMB[46][11] ), 
        .CO(\CARRYB[47][10] ), .S(\SUMB[47][10] ) );
  FA1A S2_45_38 ( .A(\ab[45][38] ), .B(\CARRYB[44][38] ), .CI(\SUMB[44][39] ), 
        .CO(\CARRYB[45][38] ), .S(\SUMB[45][38] ) );
  FA1A S2_34_40 ( .A(\ab[40][34] ), .B(\CARRYB[33][40] ), .CI(\SUMB[33][41] ), 
        .CO(\CARRYB[34][40] ), .S(\SUMB[34][40] ) );
  FA1A S2_44_30 ( .A(\ab[44][30] ), .B(\CARRYB[43][30] ), .CI(\SUMB[43][31] ), 
        .CO(\CARRYB[44][30] ), .S(\SUMB[44][30] ) );
  FA1A S2_36_30 ( .A(\ab[36][30] ), .B(\CARRYB[35][30] ), .CI(\SUMB[35][31] ), 
        .CO(\CARRYB[36][30] ), .S(\SUMB[36][30] ) );
  FA1A S2_25_42 ( .A(\ab[42][25] ), .B(\CARRYB[24][42] ), .CI(\SUMB[24][43] ), 
        .CO(\CARRYB[25][42] ), .S(\SUMB[25][42] ) );
  FA1A S2_44_38 ( .A(\ab[44][38] ), .B(\CARRYB[43][38] ), .CI(\SUMB[43][39] ), 
        .CO(\CARRYB[44][38] ), .S(\SUMB[44][38] ) );
  FA1A S3_27_46 ( .A(\ab[46][27] ), .B(\CARRYB[26][46] ), .CI(\ab[47][26] ), 
        .CO(\CARRYB[27][46] ), .S(\SUMB[27][46] ) );
  FA1A S2_46_10 ( .A(\ab[46][10] ), .B(\CARRYB[45][10] ), .CI(\SUMB[45][11] ), 
        .CO(\CARRYB[46][10] ), .S(\SUMB[46][10] ) );
  FA1A S2_23_10 ( .A(n561), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), .CO(
        \CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA1A S2_10_25 ( .A(\CARRYB[9][25] ), .B(n540), .CI(\SUMB[9][26] ), .CO(
        \CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA1A S2_17_13 ( .A(n629), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), .CO(
        \CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA1AP S2_22_14 ( .A(n646), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), .CO(
        \CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA1A S2_35_19 ( .A(\CARRYB[34][19] ), .B(\ab[35][19] ), .CI(\SUMB[34][20] ), 
        .CO(\CARRYB[35][19] ), .S(\SUMB[35][19] ) );
  FA1A S2_35_36 ( .A(\ab[36][35] ), .B(\CARRYB[34][36] ), .CI(\SUMB[34][37] ), 
        .CO(\CARRYB[35][36] ), .S(\SUMB[35][36] ) );
  FA1A S3_31_46 ( .A(\ab[46][31] ), .B(\CARRYB[30][46] ), .CI(\ab[47][30] ), 
        .CO(\CARRYB[31][46] ), .S(\SUMB[31][46] ) );
  FA1A S2_5_23 ( .A(n394), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), .CO(
        \CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA1A S2_32_20 ( .A(\ab[32][20] ), .B(\CARRYB[31][20] ), .CI(\SUMB[31][21] ), 
        .CO(\CARRYB[32][20] ), .S(\SUMB[32][20] ) );
  FA1P S2_46_5 ( .A(n388), .B(\CARRYB[45][5] ), .CI(\SUMB[45][6] ), .CO(
        \CARRYB[46][5] ), .S(\SUMB[46][5] ) );
  FA1P S2_41_5 ( .A(n385), .B(\CARRYB[40][5] ), .CI(\SUMB[40][6] ), .CO(
        \CARRYB[41][5] ), .S(\SUMB[41][5] ) );
  FA1P S1_44_0 ( .A(n306), .B(\CARRYB[43][0] ), .CI(\SUMB[43][1] ), .CO(
        \CARRYB[44][0] ), .S(\A1[42] ) );
  FA1 S2_46_17 ( .A(\ab[46][17] ), .B(\CARRYB[45][17] ), .CI(\SUMB[45][18] ), 
        .CO(\CARRYB[46][17] ), .S(\SUMB[46][17] ) );
  FA1 S2_43_40 ( .A(\ab[43][40] ), .B(\CARRYB[42][40] ), .CI(\SUMB[42][41] ), 
        .CO(\CARRYB[43][40] ), .S(\SUMB[43][40] ) );
  FA1AP S2_24_39 ( .A(\ab[39][24] ), .B(\CARRYB[23][39] ), .CI(\SUMB[23][40] ), 
        .CO(\CARRYB[24][39] ), .S(\SUMB[24][39] ) );
  FA1A S2_33_42 ( .A(\ab[42][33] ), .B(\CARRYB[32][42] ), .CI(\SUMB[32][43] ), 
        .CO(\CARRYB[33][42] ), .S(\SUMB[33][42] ) );
  FA1A S2_35_42 ( .A(\ab[42][35] ), .B(\CARRYB[34][42] ), .CI(\SUMB[34][43] ), 
        .CO(\CARRYB[35][42] ), .S(\SUMB[35][42] ) );
  FA1A S2_33_43 ( .A(\ab[43][33] ), .B(\CARRYB[32][43] ), .CI(\SUMB[32][44] ), 
        .CO(\CARRYB[33][43] ), .S(\SUMB[33][43] ) );
  FA1 S2_46_7 ( .A(\ab[7][46] ), .B(\CARRYB[45][7] ), .CI(\SUMB[45][8] ), .CO(
        \CARRYB[46][7] ), .S(\SUMB[46][7] ) );
  FA1P S2_9_44 ( .A(\ab[9][44] ), .B(\CARRYB[8][44] ), .CI(\SUMB[8][45] ), 
        .CO(\CARRYB[9][44] ), .S(\SUMB[9][44] ) );
  FA1A S2_20_30 ( .A(\ab[30][20] ), .B(\CARRYB[19][30] ), .CI(\SUMB[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA1 S2_40_13 ( .A(\ab[40][13] ), .B(\CARRYB[39][13] ), .CI(\SUMB[39][14] ), 
        .CO(\CARRYB[40][13] ), .S(\SUMB[40][13] ) );
  FA1A S2_24_13 ( .A(\CARRYB[23][13] ), .B(n631), .CI(\SUMB[23][14] ), .CO(
        \CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA1P S2_46_13 ( .A(\ab[46][13] ), .B(\CARRYB[45][13] ), .CI(\SUMB[45][14] ), 
        .CO(\CARRYB[46][13] ), .S(\SUMB[46][13] ) );
  FA1 S2_46_20 ( .A(\ab[46][20] ), .B(\CARRYB[45][20] ), .CI(\SUMB[45][21] ), 
        .CO(\CARRYB[46][20] ), .S(\SUMB[46][20] ) );
  FA1 S2_38_13 ( .A(\SUMB[37][14] ), .B(\CARRYB[37][13] ), .CI(\ab[38][13] ), 
        .CO(\CARRYB[38][13] ), .S(\SUMB[38][13] ) );
  FA1 S2_25_37 ( .A(\ab[37][25] ), .B(\CARRYB[24][37] ), .CI(\SUMB[24][38] ), 
        .CO(\CARRYB[25][37] ), .S(\SUMB[25][37] ) );
  FA1 S2_14_28 ( .A(\ab[28][14] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA1P S2_28_26 ( .A(\ab[28][26] ), .B(\CARRYB[27][26] ), .CI(\SUMB[27][27] ), 
        .CO(\CARRYB[28][26] ), .S(\SUMB[28][26] ) );
  FA1P S2_16_28 ( .A(\ab[28][16] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA1 S2_8_3 ( .A(n326), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1P S2_28_2 ( .A(n1309), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), .CO(
        \CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA1 S2_22_5 ( .A(n371), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), .CO(
        \CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA1A S2_18_3 ( .A(n1391), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), .CO(
        \CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1AP S4_17 ( .A(\ab[47][17] ), .B(\CARRYB[46][17] ), .CI(\SUMB[46][18] ), 
        .CO(\CARRYB[47][17] ), .S(\SUMB[47][17] ) );
  FA1A S2_3_8 ( .A(n326), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_6_2 ( .A(n325), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_3_2 ( .A(n301), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1P S2_29_10 ( .A(n555), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), .CO(
        \CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA1 S2_40_21 ( .A(\ab[40][21] ), .B(\CARRYB[39][21] ), .CI(\SUMB[39][22] ), 
        .CO(\CARRYB[40][21] ), .S(\SUMB[40][21] ) );
  FA1P S2_34_37 ( .A(\ab[37][34] ), .B(\CARRYB[33][37] ), .CI(\SUMB[33][38] ), 
        .CO(\CARRYB[34][37] ), .S(\SUMB[34][37] ) );
  FA1P S2_38_42 ( .A(\ab[42][38] ), .B(\CARRYB[37][42] ), .CI(\SUMB[37][43] ), 
        .CO(\CARRYB[38][42] ), .S(\SUMB[38][42] ) );
  FA1 S2_28_37 ( .A(\ab[37][28] ), .B(\CARRYB[27][37] ), .CI(\SUMB[27][38] ), 
        .CO(\CARRYB[28][37] ), .S(\SUMB[28][37] ) );
  FA1A S2_6_9 ( .A(n449), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1P S2_15_2 ( .A(n1304), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_15_3 ( .A(n1318), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1AP S4_4 ( .A(n272), .B(\CARRYB[46][4] ), .CI(\SUMB[46][5] ), .CO(
        \CARRYB[47][4] ), .S(\SUMB[47][4] ) );
  FA1A S2_5_3 ( .A(n324), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1 S2_26_1 ( .A(n1409), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), .CO(
        \CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA1A S2_8_8 ( .A(A[8]), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S3_33_46 ( .A(\ab[46][33] ), .B(\CARRYB[32][46] ), .CI(\ab[47][32] ), 
        .CO(\CARRYB[33][46] ), .S(\SUMB[33][46] ) );
  FA1 S2_10_3 ( .A(n328), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_19_4 ( .A(n1277), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), .CO(
        \CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1P S2_40_18 ( .A(\ab[40][18] ), .B(\CARRYB[39][18] ), .CI(\SUMB[39][19] ), 
        .CO(\CARRYB[40][18] ), .S(\SUMB[40][18] ) );
  FA1A S2_8_5 ( .A(n425), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_10_5 ( .A(n437), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_12_5 ( .A(n441), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), .CO(
        \CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1 S2_19_1 ( .A(n1344), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), .CO(
        \CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1A S2_5_35 ( .A(n382), .B(\CARRYB[4][35] ), .CI(\SUMB[4][36] ), .CO(
        \CARRYB[5][35] ), .S(\SUMB[5][35] ) );
  FA1P S2_8_42 ( .A(n534), .B(\CARRYB[7][42] ), .CI(\SUMB[7][43] ), .CO(
        \CARRYB[8][42] ), .S(\SUMB[8][42] ) );
  FA1P S2_25_30 ( .A(\ab[30][25] ), .B(\CARRYB[24][30] ), .CI(\SUMB[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA1P S2_44_4 ( .A(n354), .B(\CARRYB[43][4] ), .CI(\SUMB[43][5] ), .CO(
        \CARRYB[44][4] ), .S(\SUMB[44][4] ) );
  FA1AP S2_16_35 ( .A(\ab[35][16] ), .B(\CARRYB[15][35] ), .CI(\SUMB[15][36] ), 
        .CO(\CARRYB[16][35] ), .S(\SUMB[16][35] ) );
  FA1P S2_22_1 ( .A(n1393), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), .CO(
        \CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA1P S2_17_1 ( .A(n1430), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), .CO(
        \CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1P S2_12_35 ( .A(\ab[35][12] ), .B(\CARRYB[11][35] ), .CI(\SUMB[11][36] ), 
        .CO(\CARRYB[12][35] ), .S(\SUMB[12][35] ) );
  FA1AP S2_22_31 ( .A(\ab[31][22] ), .B(\CARRYB[21][31] ), .CI(\SUMB[21][32] ), 
        .CO(\CARRYB[22][31] ), .S(\SUMB[22][31] ) );
  FA1P S2_22_30 ( .A(\ab[30][22] ), .B(\CARRYB[21][30] ), .CI(\SUMB[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA1 S2_36_2 ( .A(n293), .B(\CARRYB[35][2] ), .CI(\SUMB[35][3] ), .CO(
        \CARRYB[36][2] ), .S(\SUMB[36][2] ) );
  FA1P S2_36_37 ( .A(\ab[37][36] ), .B(\CARRYB[35][37] ), .CI(\SUMB[35][38] ), 
        .CO(\CARRYB[36][37] ), .S(\SUMB[36][37] ) );
  FA1P S2_4_39 ( .A(n355), .B(\CARRYB[3][39] ), .CI(\SUMB[3][40] ), .CO(
        \CARRYB[4][39] ), .S(\SUMB[4][39] ) );
  FA1 S2_6_4 ( .A(n315), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_13_3 ( .A(n360), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), .CO(
        \CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1P S2_6_38 ( .A(n1280), .B(\CARRYB[5][38] ), .CI(\SUMB[5][39] ), .CO(
        \CARRYB[6][38] ), .S(\SUMB[6][38] ) );
  FA1P S2_5_40 ( .A(n377), .B(\CARRYB[4][40] ), .CI(\SUMB[4][41] ), .CO(
        \CARRYB[5][40] ), .S(\SUMB[5][40] ) );
  FA1P S2_6_40 ( .A(n387), .B(\CARRYB[5][40] ), .CI(\SUMB[5][41] ), .CO(
        \CARRYB[6][40] ), .S(\SUMB[6][40] ) );
  FA1 S2_39_35 ( .A(\ab[39][35] ), .B(\CARRYB[38][35] ), .CI(\SUMB[38][36] ), 
        .CO(\CARRYB[39][35] ), .S(\SUMB[39][35] ) );
  FA1P S2_2_6 ( .A(n325), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1P S2_11_35 ( .A(\ab[35][11] ), .B(\CARRYB[10][35] ), .CI(\SUMB[10][36] ), 
        .CO(\CARRYB[11][35] ), .S(\SUMB[11][35] ) );
  FA1AP S2_4_40 ( .A(n323), .B(\CARRYB[3][40] ), .CI(\SUMB[3][41] ), .CO(
        \CARRYB[4][40] ), .S(\SUMB[4][40] ) );
  FA1P S2_33_41 ( .A(\ab[41][33] ), .B(\CARRYB[32][41] ), .CI(\SUMB[32][42] ), 
        .CO(\CARRYB[33][41] ), .S(\SUMB[33][41] ) );
  FA1 S2_34_41 ( .A(\ab[41][34] ), .B(\CARRYB[33][41] ), .CI(\SUMB[33][42] ), 
        .CO(\CARRYB[34][41] ), .S(\SUMB[34][41] ) );
  FA1P S2_32_18 ( .A(\ab[32][18] ), .B(\CARRYB[31][18] ), .CI(\SUMB[31][19] ), 
        .CO(\CARRYB[32][18] ), .S(\SUMB[32][18] ) );
  FA1P S2_7_37 ( .A(n461), .B(\CARRYB[6][37] ), .CI(\SUMB[6][38] ), .CO(
        \CARRYB[7][37] ), .S(\SUMB[7][37] ) );
  FA1P S2_44_20 ( .A(\ab[44][20] ), .B(\CARRYB[43][20] ), .CI(\SUMB[43][21] ), 
        .CO(\CARRYB[44][20] ), .S(\SUMB[44][20] ) );
  FA1P S2_15_42 ( .A(\ab[42][15] ), .B(\CARRYB[14][42] ), .CI(\SUMB[14][43] ), 
        .CO(\CARRYB[15][42] ), .S(\SUMB[15][42] ) );
  FA1P S2_16_42 ( .A(\ab[42][16] ), .B(\CARRYB[15][42] ), .CI(\SUMB[15][43] ), 
        .CO(\CARRYB[16][42] ), .S(\SUMB[16][42] ) );
  FA1P S4_27 ( .A(\ab[47][27] ), .B(\CARRYB[46][27] ), .CI(\SUMB[46][28] ), 
        .CO(\CARRYB[47][27] ), .S(\SUMB[47][27] ) );
  FA1P S2_33_18 ( .A(\ab[33][18] ), .B(\CARRYB[32][18] ), .CI(\SUMB[32][19] ), 
        .CO(\CARRYB[33][18] ), .S(\SUMB[33][18] ) );
  FA1 S2_33_40 ( .A(\ab[40][33] ), .B(\CARRYB[32][40] ), .CI(\SUMB[32][41] ), 
        .CO(\CARRYB[33][40] ), .S(\SUMB[33][40] ) );
  FA1P S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA1 S2_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\SUMB[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA1P S2_40_30 ( .A(\ab[40][30] ), .B(\CARRYB[39][30] ), .CI(\SUMB[39][31] ), 
        .CO(\CARRYB[40][30] ), .S(\SUMB[40][30] ) );
  FA1AP S2_44_5 ( .A(n415), .B(\CARRYB[43][5] ), .CI(\SUMB[43][6] ), .CO(
        \CARRYB[44][5] ), .S(\SUMB[44][5] ) );
  FA1P S2_45_5 ( .A(n401), .B(\CARRYB[44][5] ), .CI(\SUMB[44][6] ), .CO(
        \CARRYB[45][5] ), .S(\SUMB[45][5] ) );
  FA1P S2_44_13 ( .A(\ab[44][13] ), .B(\CARRYB[43][13] ), .CI(\SUMB[43][14] ), 
        .CO(\CARRYB[44][13] ), .S(\SUMB[44][13] ) );
  FA1P S2_45_13 ( .A(\ab[45][13] ), .B(\CARRYB[44][13] ), .CI(\SUMB[44][14] ), 
        .CO(\CARRYB[45][13] ), .S(\SUMB[45][13] ) );
  FA1P S2_18_23 ( .A(\ab[23][18] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA1P S2_35_17 ( .A(\ab[35][17] ), .B(\CARRYB[34][17] ), .CI(\SUMB[34][18] ), 
        .CO(\CARRYB[35][17] ), .S(\SUMB[35][17] ) );
  FA1P S2_19_22 ( .A(\ab[22][19] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA1P S2_20_22 ( .A(\ab[22][20] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA1P S2_44_27 ( .A(\ab[44][27] ), .B(\CARRYB[43][27] ), .CI(\SUMB[43][28] ), 
        .CO(\CARRYB[44][27] ), .S(\SUMB[44][27] ) );
  FA1 S2_27_3 ( .A(n292), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), .CO(
        \CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA1P S2_42_2 ( .A(n1328), .B(\CARRYB[41][2] ), .CI(\SUMB[41][3] ), .CO(
        \CARRYB[42][2] ), .S(\SUMB[42][2] ) );
  FA1P S2_9_42 ( .A(\ab[9][42] ), .B(\CARRYB[8][42] ), .CI(\SUMB[8][43] ), 
        .CO(\CARRYB[9][42] ), .S(\SUMB[9][42] ) );
  FA1P S2_35_37 ( .A(\ab[37][35] ), .B(\CARRYB[34][37] ), .CI(\SUMB[34][38] ), 
        .CO(\CARRYB[35][37] ), .S(\SUMB[35][37] ) );
  FA1 S2_43_5 ( .A(n399), .B(\CARRYB[42][5] ), .CI(\SUMB[42][6] ), .CO(
        \CARRYB[43][5] ), .S(\SUMB[43][5] ) );
  FA1P S2_40_23 ( .A(\ab[40][23] ), .B(\CARRYB[39][23] ), .CI(\SUMB[39][24] ), 
        .CO(\CARRYB[40][23] ), .S(\SUMB[40][23] ) );
  FA1 S2_37_7 ( .A(n461), .B(\CARRYB[36][7] ), .CI(\SUMB[36][8] ), .CO(
        \CARRYB[37][7] ), .S(\SUMB[37][7] ) );
  FA1P S2_42_25 ( .A(\ab[42][25] ), .B(\CARRYB[41][25] ), .CI(\SUMB[41][26] ), 
        .CO(\CARRYB[42][25] ), .S(\SUMB[42][25] ) );
  FA1 S2_38_12 ( .A(\CARRYB[37][12] ), .B(\ab[38][12] ), .CI(\SUMB[37][13] ), 
        .CO(\CARRYB[38][12] ), .S(\SUMB[38][12] ) );
  FA1AP S2_45_31 ( .A(\ab[45][31] ), .B(\CARRYB[44][31] ), .CI(\SUMB[44][32] ), 
        .CO(\CARRYB[45][31] ), .S(\SUMB[45][31] ) );
  FA1P S2_9_34 ( .A(n539), .B(\CARRYB[8][34] ), .CI(\SUMB[8][35] ), .CO(
        \CARRYB[9][34] ), .S(\SUMB[9][34] ) );
  FA1P S2_10_34 ( .A(n564), .B(\CARRYB[9][34] ), .CI(\SUMB[9][35] ), .CO(
        \CARRYB[10][34] ), .S(\SUMB[10][34] ) );
  FA1A S2_29_41 ( .A(\ab[41][29] ), .B(\CARRYB[28][41] ), .CI(\SUMB[28][42] ), 
        .CO(\CARRYB[29][41] ), .S(\SUMB[29][41] ) );
  FA1A S2_45_22 ( .A(\ab[45][22] ), .B(\CARRYB[44][22] ), .CI(\SUMB[44][23] ), 
        .CO(\CARRYB[45][22] ), .S(\SUMB[45][22] ) );
  FA1AP S2_23_11 ( .A(n582), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), .CO(
        \CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA1P S2_35_28 ( .A(\CARRYB[34][28] ), .B(\ab[35][28] ), .CI(\SUMB[34][29] ), 
        .CO(\CARRYB[35][28] ), .S(\SUMB[35][28] ) );
  FA1P S2_2_23 ( .A(n302), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), .CO(
        \CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA1 S2_24_42 ( .A(\ab[42][24] ), .B(\CARRYB[23][42] ), .CI(\SUMB[23][43] ), 
        .CO(\CARRYB[24][42] ), .S(\SUMB[24][42] ) );
  FA1P S2_7_43 ( .A(n279), .B(\CARRYB[6][43] ), .CI(\SUMB[6][44] ), .CO(
        \CARRYB[7][43] ), .S(\SUMB[7][43] ) );
  FA1P S2_8_44 ( .A(\ab[8][44] ), .B(\CARRYB[7][44] ), .CI(\SUMB[7][45] ), 
        .CO(\CARRYB[8][44] ), .S(\SUMB[8][44] ) );
  FA1P S2_33_24 ( .A(\ab[33][24] ), .B(\CARRYB[32][24] ), .CI(\SUMB[32][25] ), 
        .CO(\CARRYB[33][24] ), .S(\SUMB[33][24] ) );
  FA1P S2_18_12 ( .A(n599), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), .CO(
        \CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA1P S2_21_17 ( .A(\SUMB[20][18] ), .B(\CARRYB[20][17] ), .CI(\ab[21][17] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA1P S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA1P S2_33_1 ( .A(n1372), .B(\CARRYB[32][1] ), .CI(\SUMB[32][2] ), .CO(
        \CARRYB[33][1] ), .S(\SUMB[33][1] ) );
  FA1P S2_17_17 ( .A(n1464), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), .CO(
        \CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA1P S2_37_38 ( .A(\ab[38][37] ), .B(\CARRYB[36][38] ), .CI(\SUMB[36][39] ), 
        .CO(\CARRYB[37][38] ), .S(\SUMB[37][38] ) );
  FA1P S2_31_8 ( .A(n485), .B(\CARRYB[30][8] ), .CI(\SUMB[30][9] ), .CO(
        \CARRYB[31][8] ), .S(\SUMB[31][8] ) );
  FA1P S2_32_8 ( .A(n278), .B(\CARRYB[31][8] ), .CI(\SUMB[31][9] ), .CO(
        \CARRYB[32][8] ), .S(\SUMB[32][8] ) );
  FA1P S2_24_37 ( .A(\ab[37][24] ), .B(\CARRYB[23][37] ), .CI(\SUMB[23][38] ), 
        .CO(\CARRYB[24][37] ), .S(\SUMB[24][37] ) );
  FA1 S2_12_39 ( .A(\SUMB[11][40] ), .B(\CARRYB[11][39] ), .CI(\ab[39][12] ), 
        .CO(\CARRYB[12][39] ), .S(\SUMB[12][39] ) );
  FA1P S2_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\SUMB[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA1P S2_34_7 ( .A(n477), .B(\CARRYB[33][7] ), .CI(\SUMB[33][8] ), .CO(
        \CARRYB[34][7] ), .S(\SUMB[34][7] ) );
  FA1P S2_35_7 ( .A(n417), .B(\CARRYB[34][7] ), .CI(\SUMB[34][8] ), .CO(
        \CARRYB[35][7] ), .S(\SUMB[35][7] ) );
  FA1P S2_26_32 ( .A(\ab[32][26] ), .B(\CARRYB[25][32] ), .CI(\SUMB[25][33] ), 
        .CO(\CARRYB[26][32] ), .S(\SUMB[26][32] ) );
  FA1A S2_13_26 ( .A(n616), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), .CO(
        \CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA1AP S2_14_26 ( .A(n645), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), .CO(
        \CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA1P S2_40_4 ( .A(n323), .B(\CARRYB[39][4] ), .CI(\SUMB[39][5] ), .CO(
        \CARRYB[40][4] ), .S(\SUMB[40][4] ) );
  FA1P S2_41_4 ( .A(n320), .B(\CARRYB[40][4] ), .CI(\SUMB[40][5] ), .CO(
        \CARRYB[41][4] ), .S(\SUMB[41][4] ) );
  FA1P S2_11_18 ( .A(n584), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), .CO(
        \CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1P S2_46_19 ( .A(\ab[46][19] ), .B(\CARRYB[45][19] ), .CI(\SUMB[45][20] ), 
        .CO(\CARRYB[46][19] ), .S(\SUMB[46][19] ) );
  FA1P S4_19 ( .A(\ab[47][19] ), .B(\CARRYB[46][19] ), .CI(\SUMB[46][20] ), 
        .CO(\CARRYB[47][19] ), .S(\SUMB[47][19] ) );
  FA1 S2_17_35 ( .A(\ab[35][17] ), .B(\CARRYB[16][35] ), .CI(\SUMB[16][36] ), 
        .CO(\CARRYB[17][35] ), .S(\SUMB[17][35] ) );
  FA1 S2_22_10 ( .A(n281), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), .CO(
        \CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA1 S2_2_45 ( .A(n1314), .B(\CARRYB[1][45] ), .CI(\SUMB[1][46] ), .CO(
        \CARRYB[2][45] ), .S(\SUMB[2][45] ) );
  FA1P S2_7_40 ( .A(n418), .B(\CARRYB[6][40] ), .CI(\SUMB[6][41] ), .CO(
        \CARRYB[7][40] ), .S(\SUMB[7][40] ) );
  FA1P S2_6_43 ( .A(n447), .B(\CARRYB[5][43] ), .CI(\SUMB[5][44] ), .CO(
        \CARRYB[6][43] ), .S(\SUMB[6][43] ) );
  FA1P S2_24_36 ( .A(\ab[36][24] ), .B(\CARRYB[23][36] ), .CI(\SUMB[23][37] ), 
        .CO(\CARRYB[24][36] ), .S(\SUMB[24][36] ) );
  FA1P S2_30_2 ( .A(n290), .B(\CARRYB[29][2] ), .CI(\SUMB[29][3] ), .CO(
        \CARRYB[30][2] ), .S(\SUMB[30][2] ) );
  FA1P S2_31_2 ( .A(n1340), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), .CO(
        \CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FA1 S2_25_3 ( .A(n284), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), .CO(
        \CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA1AP S2_2_26 ( .A(n299), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), .CO(
        \CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA1AP S2_19_36 ( .A(\CARRYB[18][36] ), .B(\ab[36][19] ), .CI(\SUMB[18][37] ), 
        .CO(\CARRYB[19][36] ), .S(\SUMB[19][36] ) );
  FA1AP S2_13_20 ( .A(n615), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), .CO(
        \CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA1P S2_18_19 ( .A(\SUMB[17][20] ), .B(\CARRYB[17][19] ), .CI(\ab[19][18] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA1AP S2_22_16 ( .A(\CARRYB[21][16] ), .B(\ab[22][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA1P S2_45_32 ( .A(\ab[45][32] ), .B(\CARRYB[44][32] ), .CI(\SUMB[44][33] ), 
        .CO(\CARRYB[45][32] ), .S(\SUMB[45][32] ) );
  FA1AP S2_14_35 ( .A(\ab[35][14] ), .B(\CARRYB[13][35] ), .CI(\SUMB[13][36] ), 
        .CO(\CARRYB[14][35] ), .S(\SUMB[14][35] ) );
  FA1 S2_34_18 ( .A(\ab[34][18] ), .B(\CARRYB[33][18] ), .CI(\SUMB[33][19] ), 
        .CO(\CARRYB[34][18] ), .S(\SUMB[34][18] ) );
  FA1AP S2_17_38 ( .A(\ab[38][17] ), .B(\CARRYB[16][38] ), .CI(\SUMB[16][39] ), 
        .CO(\CARRYB[17][38] ), .S(\SUMB[17][38] ) );
  FA1P S2_32_11 ( .A(n577), .B(\CARRYB[31][11] ), .CI(\SUMB[31][12] ), .CO(
        \CARRYB[32][11] ), .S(\SUMB[32][11] ) );
  FA1AP S4_14 ( .A(\ab[47][14] ), .B(\CARRYB[46][14] ), .CI(\SUMB[46][15] ), 
        .CO(\CARRYB[47][14] ), .S(\SUMB[47][14] ) );
  FA1P S2_11_24 ( .A(n588), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), .CO(
        \CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA1 S2_8_33 ( .A(n489), .B(\CARRYB[7][33] ), .CI(\SUMB[7][34] ), .CO(
        \CARRYB[8][33] ), .S(\SUMB[8][33] ) );
  FA1 S2_38_26 ( .A(\SUMB[37][27] ), .B(\CARRYB[37][26] ), .CI(\ab[38][26] ), 
        .CO(\CARRYB[38][26] ), .S(\SUMB[38][26] ) );
  FA1 S2_31_42 ( .A(\ab[42][31] ), .B(\CARRYB[30][42] ), .CI(\SUMB[30][43] ), 
        .CO(\CARRYB[31][42] ), .S(\SUMB[31][42] ) );
  FA1P S2_32_42 ( .A(\ab[42][32] ), .B(\CARRYB[31][42] ), .CI(\SUMB[31][43] ), 
        .CO(\CARRYB[32][42] ), .S(\SUMB[32][42] ) );
  FA1 S2_40_41 ( .A(\ab[41][40] ), .B(\CARRYB[39][41] ), .CI(\SUMB[39][42] ), 
        .CO(\CARRYB[40][41] ), .S(\SUMB[40][41] ) );
  FA1P S2_25_11 ( .A(n563), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), .CO(
        \CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA1 S2_45_10 ( .A(\ab[45][10] ), .B(\CARRYB[44][10] ), .CI(\SUMB[44][11] ), 
        .CO(\CARRYB[45][10] ), .S(\SUMB[45][10] ) );
  FA1A S2_6_30 ( .A(n373), .B(\CARRYB[5][30] ), .CI(\SUMB[5][31] ), .CO(
        \CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA1P S2_15_28 ( .A(\ab[28][15] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA1P S2_16_6 ( .A(n431), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), .CO(
        \CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1P S2_39_27 ( .A(\ab[39][27] ), .B(\CARRYB[38][27] ), .CI(\SUMB[38][28] ), 
        .CO(\CARRYB[39][27] ), .S(\SUMB[39][27] ) );
  FA1A S2_33_19 ( .A(\ab[33][19] ), .B(\CARRYB[32][19] ), .CI(\SUMB[32][20] ), 
        .CO(\CARRYB[33][19] ), .S(\SUMB[33][19] ) );
  FA1P S2_45_17 ( .A(\ab[45][17] ), .B(\CARRYB[44][17] ), .CI(\SUMB[44][18] ), 
        .CO(\CARRYB[45][17] ), .S(\SUMB[45][17] ) );
  FA1P S2_9_15 ( .A(n527), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), .CO(
        \CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1P S2_24_11 ( .A(n588), .B(\CARRYB[23][11] ), .CI(\SUMB[23][12] ), .CO(
        \CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA1P S4_3 ( .A(n270), .B(\CARRYB[46][3] ), .CI(\SUMB[46][4] ), .CO(
        \CARRYB[47][3] ), .S(\SUMB[47][3] ) );
  FA1P S2_27_10 ( .A(n520), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), .CO(
        \CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA1A S2_9_35 ( .A(n496), .B(\CARRYB[8][35] ), .CI(\SUMB[8][36] ), .CO(
        \CARRYB[9][35] ), .S(\SUMB[9][35] ) );
  FA1P S2_14_34 ( .A(\ab[34][14] ), .B(\CARRYB[13][34] ), .CI(\SUMB[13][35] ), 
        .CO(\CARRYB[14][34] ), .S(\SUMB[14][34] ) );
  FA1AP S2_37_30 ( .A(\CARRYB[36][30] ), .B(\ab[37][30] ), .CI(\SUMB[36][31] ), 
        .CO(\CARRYB[37][30] ), .S(\SUMB[37][30] ) );
  FA1 S2_32_19 ( .A(\ab[32][19] ), .B(\CARRYB[31][19] ), .CI(\SUMB[31][20] ), 
        .CO(\CARRYB[32][19] ), .S(\SUMB[32][19] ) );
  FA1P S2_41_18 ( .A(\ab[41][18] ), .B(\CARRYB[40][18] ), .CI(\SUMB[40][19] ), 
        .CO(\CARRYB[41][18] ), .S(\SUMB[41][18] ) );
  FA1P S2_20_13 ( .A(n615), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), .CO(
        \CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA1P S2_21_13 ( .A(n626), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), .CO(
        \CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA1P S2_45_16 ( .A(\ab[45][16] ), .B(\CARRYB[44][16] ), .CI(\SUMB[44][17] ), 
        .CO(\CARRYB[45][16] ), .S(\SUMB[45][16] ) );
  FA1 S2_9_40 ( .A(\ab[9][40] ), .B(\CARRYB[8][40] ), .CI(\SUMB[8][41] ), .CO(
        \CARRYB[9][40] ), .S(\SUMB[9][40] ) );
  FA1P S2_44_16 ( .A(\ab[44][16] ), .B(\CARRYB[43][16] ), .CI(\SUMB[43][17] ), 
        .CO(\CARRYB[44][16] ), .S(\SUMB[44][16] ) );
  FA1P S2_35_29 ( .A(\ab[35][29] ), .B(\CARRYB[34][29] ), .CI(\SUMB[34][30] ), 
        .CO(\CARRYB[35][29] ), .S(\SUMB[35][29] ) );
  FA1P S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA1P S2_35_20 ( .A(\ab[35][20] ), .B(\CARRYB[34][20] ), .CI(\SUMB[34][21] ), 
        .CO(\CARRYB[35][20] ), .S(\SUMB[35][20] ) );
  FA1 S2_34_13 ( .A(\CARRYB[33][13] ), .B(\ab[34][13] ), .CI(\SUMB[33][14] ), 
        .CO(\CARRYB[34][13] ), .S(\SUMB[34][13] ) );
  FA1P S2_44_10 ( .A(\ab[44][10] ), .B(\CARRYB[43][10] ), .CI(\SUMB[43][11] ), 
        .CO(\CARRYB[44][10] ), .S(\SUMB[44][10] ) );
  FA1P S2_36_27 ( .A(\SUMB[35][28] ), .B(\CARRYB[35][27] ), .CI(\ab[36][27] ), 
        .CO(\CARRYB[36][27] ), .S(\SUMB[36][27] ) );
  FA1P S2_45_25 ( .A(\ab[45][25] ), .B(\CARRYB[44][25] ), .CI(\SUMB[44][26] ), 
        .CO(\CARRYB[45][25] ), .S(\SUMB[45][25] ) );
  FA1P S2_13_18 ( .A(n623), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), .CO(
        \CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA1A S2_46_4 ( .A(n334), .B(\CARRYB[45][4] ), .CI(\SUMB[45][5] ), .CO(
        \CARRYB[46][4] ), .S(\SUMB[46][4] ) );
  FA1P S2_37_24 ( .A(\ab[37][24] ), .B(\CARRYB[36][24] ), .CI(\SUMB[36][25] ), 
        .CO(\CARRYB[37][24] ), .S(\SUMB[37][24] ) );
  FA1P S2_30_26 ( .A(\ab[30][26] ), .B(\CARRYB[29][26] ), .CI(\SUMB[29][27] ), 
        .CO(\CARRYB[30][26] ), .S(\SUMB[30][26] ) );
  FA1P S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA1P S2_38_24 ( .A(\ab[38][24] ), .B(\CARRYB[37][24] ), .CI(\SUMB[37][25] ), 
        .CO(\CARRYB[38][24] ), .S(\SUMB[38][24] ) );
  FA1 S1_27_0 ( .A(n1367), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), .CO(
        \CARRYB[27][0] ), .S(\A1[25] ) );
  FA1P S2_16_1 ( .A(n1427), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), .CO(
        \CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1AP S2_33_13 ( .A(\ab[33][13] ), .B(\CARRYB[32][13] ), .CI(\SUMB[32][14] ), 
        .CO(\CARRYB[33][13] ), .S(\SUMB[33][13] ) );
  FA1 S2_12_21 ( .A(\CARRYB[11][21] ), .B(n596), .CI(\SUMB[11][22] ), .CO(
        \CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA1P S2_37_31 ( .A(\ab[37][31] ), .B(\CARRYB[36][31] ), .CI(\SUMB[36][32] ), 
        .CO(\CARRYB[37][31] ), .S(\SUMB[37][31] ) );
  FA1 S2_43_30 ( .A(\ab[43][30] ), .B(\CARRYB[42][30] ), .CI(\SUMB[42][31] ), 
        .CO(\CARRYB[43][30] ), .S(\SUMB[43][30] ) );
  FA1P S2_22_40 ( .A(\ab[40][22] ), .B(\CARRYB[21][40] ), .CI(\SUMB[21][41] ), 
        .CO(\CARRYB[22][40] ), .S(\SUMB[22][40] ) );
  FA1P S2_22_39 ( .A(\ab[39][22] ), .B(\CARRYB[21][39] ), .CI(\SUMB[21][40] ), 
        .CO(\CARRYB[22][39] ), .S(\SUMB[22][39] ) );
  FA1AP S2_39_13 ( .A(\ab[39][13] ), .B(\CARRYB[38][13] ), .CI(\SUMB[38][14] ), 
        .CO(\CARRYB[39][13] ), .S(\SUMB[39][13] ) );
  FA1 S2_40_12 ( .A(\ab[40][12] ), .B(\CARRYB[39][12] ), .CI(\SUMB[39][13] ), 
        .CO(\CARRYB[40][12] ), .S(\SUMB[40][12] ) );
  FA1P S2_9_20 ( .A(n525), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), .CO(
        \CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1P S2_14_20 ( .A(n637), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), .CO(
        \CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA1P S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA1P S2_16_36 ( .A(\ab[36][16] ), .B(\CARRYB[15][36] ), .CI(\SUMB[15][37] ), 
        .CO(\CARRYB[16][36] ), .S(\SUMB[16][36] ) );
  FA1A S2_8_38 ( .A(n1293), .B(\CARRYB[7][38] ), .CI(\SUMB[7][39] ), .CO(
        \CARRYB[8][38] ), .S(\SUMB[8][38] ) );
  FA1AP S4_25 ( .A(\ab[47][25] ), .B(\CARRYB[46][25] ), .CI(\SUMB[46][26] ), 
        .CO(\CARRYB[47][25] ), .S(\SUMB[47][25] ) );
  FA1P S2_46_2 ( .A(n1308), .B(\CARRYB[45][2] ), .CI(\SUMB[45][3] ), .CO(
        \CARRYB[46][2] ), .S(\SUMB[46][2] ) );
  FA1 S2_30_20 ( .A(\ab[30][20] ), .B(\CARRYB[29][20] ), .CI(\SUMB[29][21] ), 
        .CO(\CARRYB[30][20] ), .S(\SUMB[30][20] ) );
  FA1AP S2_31_20 ( .A(\ab[31][20] ), .B(\CARRYB[30][20] ), .CI(\SUMB[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FA1AP S2_29_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA1P S2_21_27 ( .A(\ab[27][21] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA1P S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA1P S2_43_13 ( .A(\ab[43][13] ), .B(\CARRYB[42][13] ), .CI(\SUMB[42][14] ), 
        .CO(\CARRYB[43][13] ), .S(\SUMB[43][13] ) );
  FA1 S2_12_30 ( .A(\SUMB[11][31] ), .B(\CARRYB[11][30] ), .CI(n598), .CO(
        \CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA1AP S2_18_25 ( .A(\ab[25][18] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA1AP S2_37_18 ( .A(\ab[37][18] ), .B(\CARRYB[36][18] ), .CI(\SUMB[36][19] ), 
        .CO(\CARRYB[37][18] ), .S(\SUMB[37][18] ) );
  FA1 S2_40_16 ( .A(\ab[40][16] ), .B(\CARRYB[39][16] ), .CI(\SUMB[39][17] ), 
        .CO(\CARRYB[40][16] ), .S(\SUMB[40][16] ) );
  FA1 S2_25_22 ( .A(\CARRYB[24][22] ), .B(\ab[25][22] ), .CI(\SUMB[24][23] ), 
        .CO(\CARRYB[25][22] ), .S(\SUMB[25][22] ) );
  FA1P S2_7_19 ( .A(n451), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), .CO(
        \CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1P S2_16_18 ( .A(\ab[18][16] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA1AP S2_20_23 ( .A(\CARRYB[19][23] ), .B(\ab[23][20] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA1P S2_38_27 ( .A(\ab[38][27] ), .B(\CARRYB[37][27] ), .CI(\SUMB[37][28] ), 
        .CO(\CARRYB[38][27] ), .S(\SUMB[38][27] ) );
  FA1 S2_38_17 ( .A(\ab[38][17] ), .B(\CARRYB[37][17] ), .CI(\SUMB[37][18] ), 
        .CO(\CARRYB[38][17] ), .S(\SUMB[38][17] ) );
  FA1 S2_30_16 ( .A(\CARRYB[29][16] ), .B(\ab[30][16] ), .CI(\SUMB[29][17] ), 
        .CO(\CARRYB[30][16] ), .S(\SUMB[30][16] ) );
  FA1P S2_45_12 ( .A(\ab[45][12] ), .B(\CARRYB[44][12] ), .CI(\SUMB[44][13] ), 
        .CO(\CARRYB[45][12] ), .S(\SUMB[45][12] ) );
  FA1P S2_44_12 ( .A(\ab[44][12] ), .B(\CARRYB[43][12] ), .CI(\SUMB[43][13] ), 
        .CO(\CARRYB[44][12] ), .S(\SUMB[44][12] ) );
  FA1P S2_44_24 ( .A(\ab[44][24] ), .B(\CARRYB[43][24] ), .CI(\SUMB[43][25] ), 
        .CO(\CARRYB[44][24] ), .S(\SUMB[44][24] ) );
  FA1P S2_46_24 ( .A(\ab[46][24] ), .B(\CARRYB[45][24] ), .CI(\SUMB[45][25] ), 
        .CO(\CARRYB[46][24] ), .S(\SUMB[46][24] ) );
  FA1P S2_8_7 ( .A(n493), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1P S2_32_6 ( .A(n395), .B(\CARRYB[31][6] ), .CI(\SUMB[31][7] ), .CO(
        \CARRYB[32][6] ), .S(\SUMB[32][6] ) );
  FA1P S2_12_7 ( .A(n510), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), .CO(
        \CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1P S2_13_7 ( .A(n465), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), .CO(
        \CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1P S2_43_27 ( .A(\ab[43][27] ), .B(\CARRYB[42][27] ), .CI(\SUMB[42][28] ), 
        .CO(\CARRYB[43][27] ), .S(\SUMB[43][27] ) );
  FA1P S2_11_39 ( .A(\ab[39][11] ), .B(\CARRYB[10][39] ), .CI(\SUMB[10][40] ), 
        .CO(\CARRYB[11][39] ), .S(\SUMB[11][39] ) );
  FA1A S2_12_38 ( .A(\ab[38][12] ), .B(\CARRYB[11][38] ), .CI(\SUMB[11][39] ), 
        .CO(\CARRYB[12][38] ), .S(\SUMB[12][38] ) );
  FA1 S2_32_23 ( .A(\ab[32][23] ), .B(\CARRYB[31][23] ), .CI(\SUMB[31][24] ), 
        .CO(\CARRYB[32][23] ), .S(\SUMB[32][23] ) );
  FA1 S2_11_38 ( .A(\SUMB[10][39] ), .B(\CARRYB[10][38] ), .CI(\ab[38][11] ), 
        .CO(\CARRYB[11][38] ), .S(\SUMB[11][38] ) );
  FA1 S2_15_25 ( .A(\CARRYB[14][25] ), .B(\ab[25][15] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA1A S2_33_23 ( .A(\ab[33][23] ), .B(\CARRYB[32][23] ), .CI(\SUMB[32][24] ), 
        .CO(\CARRYB[33][23] ), .S(\SUMB[33][23] ) );
  FA1AP S2_19_34 ( .A(\ab[34][19] ), .B(\CARRYB[18][34] ), .CI(\SUMB[18][35] ), 
        .CO(\CARRYB[19][34] ), .S(\SUMB[19][34] ) );
  FA1P S2_14_31 ( .A(\ab[31][14] ), .B(\CARRYB[13][31] ), .CI(\SUMB[13][32] ), 
        .CO(\CARRYB[14][31] ), .S(\SUMB[14][31] ) );
  FA1 S2_5_24 ( .A(\CARRYB[4][24] ), .B(n1275), .CI(\SUMB[4][25] ), .CO(
        \CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA1A S2_4_36 ( .A(n367), .B(\CARRYB[3][36] ), .CI(\SUMB[3][37] ), .CO(
        \CARRYB[4][36] ), .S(\SUMB[4][36] ) );
  FA1P S2_9_2 ( .A(n316), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1 S2_10_2 ( .A(n303), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1AP S2_37_14 ( .A(\ab[37][14] ), .B(\CARRYB[36][14] ), .CI(\SUMB[36][15] ), 
        .CO(\CARRYB[37][14] ), .S(\SUMB[37][14] ) );
  FA1P S2_43_26 ( .A(\ab[43][26] ), .B(\CARRYB[42][26] ), .CI(\SUMB[42][27] ), 
        .CO(\CARRYB[43][26] ), .S(\SUMB[43][26] ) );
  FA1P S2_34_30 ( .A(\ab[34][30] ), .B(\CARRYB[33][30] ), .CI(\SUMB[33][31] ), 
        .CO(\CARRYB[34][30] ), .S(\SUMB[34][30] ) );
  FA1 S2_7_15 ( .A(n471), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), .CO(
        \CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1 S2_36_12 ( .A(\ab[36][12] ), .B(\CARRYB[35][12] ), .CI(\SUMB[35][13] ), 
        .CO(\CARRYB[36][12] ), .S(\SUMB[36][12] ) );
  FA1P S2_36_24 ( .A(\ab[36][24] ), .B(\CARRYB[35][24] ), .CI(\SUMB[35][25] ), 
        .CO(\CARRYB[36][24] ), .S(\SUMB[36][24] ) );
  FA1P S2_42_22 ( .A(\ab[42][22] ), .B(\CARRYB[41][22] ), .CI(\SUMB[41][23] ), 
        .CO(\CARRYB[42][22] ), .S(\SUMB[42][22] ) );
  FA1P S2_43_22 ( .A(\ab[43][22] ), .B(\CARRYB[42][22] ), .CI(\SUMB[42][23] ), 
        .CO(\CARRYB[43][22] ), .S(\SUMB[43][22] ) );
  FA1P S2_9_37 ( .A(n546), .B(\CARRYB[8][37] ), .CI(\SUMB[8][38] ), .CO(
        \CARRYB[9][37] ), .S(\SUMB[9][37] ) );
  FA1 S2_21_31 ( .A(\ab[31][21] ), .B(\CARRYB[20][31] ), .CI(\SUMB[20][32] ), 
        .CO(\CARRYB[21][31] ), .S(\SUMB[21][31] ) );
  FA1 S2_8_29 ( .A(\CARRYB[7][29] ), .B(n1290), .CI(\SUMB[7][30] ), .CO(
        \CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA1AP S2_42_13 ( .A(\ab[42][13] ), .B(\CARRYB[41][13] ), .CI(\SUMB[41][14] ), 
        .CO(\CARRYB[42][13] ), .S(\SUMB[42][13] ) );
  FA1A S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA1P S2_29_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA1 S2_16_26 ( .A(\CARRYB[15][26] ), .B(\ab[26][16] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA1 S2_15_29 ( .A(\CARRYB[14][29] ), .B(\ab[29][15] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA1A S2_41_11 ( .A(\ab[41][11] ), .B(\CARRYB[40][11] ), .CI(\SUMB[40][12] ), 
        .CO(\CARRYB[41][11] ), .S(\SUMB[41][11] ) );
  FA1P S2_15_39 ( .A(\CARRYB[14][39] ), .B(\ab[39][15] ), .CI(\SUMB[14][40] ), 
        .CO(\CARRYB[15][39] ), .S(\SUMB[15][39] ) );
  FA1P S2_39_14 ( .A(\ab[39][14] ), .B(\CARRYB[38][14] ), .CI(\SUMB[38][15] ), 
        .CO(\CARRYB[39][14] ), .S(\SUMB[39][14] ) );
  FA1 S2_29_14 ( .A(\CARRYB[28][14] ), .B(\ab[29][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA1P S2_5_18 ( .A(n398), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), .CO(
        \CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1P S2_6_18 ( .A(n428), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), .CO(
        \CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1P S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA1A S2_26_21 ( .A(\CARRYB[25][21] ), .B(\ab[26][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA1 S2_36_14 ( .A(\ab[36][14] ), .B(\CARRYB[35][14] ), .CI(\SUMB[35][15] ), 
        .CO(\CARRYB[36][14] ), .S(\SUMB[36][14] ) );
  FA1A S2_23_42 ( .A(\ab[42][23] ), .B(\CARRYB[22][42] ), .CI(\SUMB[22][43] ), 
        .CO(\CARRYB[23][42] ), .S(\SUMB[23][42] ) );
  FA1A S2_32_40 ( .A(\ab[40][32] ), .B(\CARRYB[31][40] ), .CI(\SUMB[31][41] ), 
        .CO(\CARRYB[32][40] ), .S(\SUMB[32][40] ) );
  FA1AP S2_11_40 ( .A(\ab[40][11] ), .B(\CARRYB[10][40] ), .CI(\SUMB[10][41] ), 
        .CO(\CARRYB[11][40] ), .S(\SUMB[11][40] ) );
  FA1 S2_6_29 ( .A(\CARRYB[5][29] ), .B(n1279), .CI(\SUMB[5][30] ), .CO(
        \CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA1P S2_11_19 ( .A(n572), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), .CO(
        \CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1P S2_39_28 ( .A(\ab[39][28] ), .B(\CARRYB[38][28] ), .CI(\SUMB[38][29] ), 
        .CO(\CARRYB[39][28] ), .S(\SUMB[39][28] ) );
  FA1A S2_10_37 ( .A(n567), .B(\CARRYB[9][37] ), .CI(\SUMB[9][38] ), .CO(
        \CARRYB[10][37] ), .S(\SUMB[10][37] ) );
  FA1A S2_21_33 ( .A(\ab[33][21] ), .B(\CARRYB[20][33] ), .CI(\SUMB[20][34] ), 
        .CO(\CARRYB[21][33] ), .S(\SUMB[21][33] ) );
  FA1 S2_10_30 ( .A(n507), .B(\CARRYB[9][30] ), .CI(\SUMB[9][31] ), .CO(
        \CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA1A S2_15_37 ( .A(\ab[37][15] ), .B(\CARRYB[14][37] ), .CI(\SUMB[14][38] ), 
        .CO(\CARRYB[15][37] ), .S(\SUMB[15][37] ) );
  FA1 S2_37_15 ( .A(\ab[37][15] ), .B(\CARRYB[36][15] ), .CI(\SUMB[36][16] ), 
        .CO(\CARRYB[37][15] ), .S(\SUMB[37][15] ) );
  FA1P S2_25_31 ( .A(\ab[31][25] ), .B(\CARRYB[24][31] ), .CI(\SUMB[24][32] ), 
        .CO(\CARRYB[25][31] ), .S(\SUMB[25][31] ) );
  FA1P S2_36_29 ( .A(\ab[36][29] ), .B(\CARRYB[35][29] ), .CI(\SUMB[35][30] ), 
        .CO(\CARRYB[36][29] ), .S(\SUMB[36][29] ) );
  FA1P S2_13_25 ( .A(n625), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), .CO(
        \CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA1P S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA1P S2_14_25 ( .A(\CARRYB[13][25] ), .B(n635), .CI(\SUMB[13][26] ), .CO(
        \CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA1A S2_39_26 ( .A(\ab[39][26] ), .B(\CARRYB[38][26] ), .CI(\SUMB[38][27] ), 
        .CO(\CARRYB[39][26] ), .S(\SUMB[39][26] ) );
  FA1P S2_16_12 ( .A(n612), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), .CO(
        \CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA1P S2_31_9 ( .A(n524), .B(\CARRYB[30][9] ), .CI(\SUMB[30][10] ), .CO(
        \CARRYB[31][9] ), .S(\SUMB[31][9] ) );
  FA1P S2_21_26 ( .A(\ab[26][21] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA1P S2_22_26 ( .A(\ab[26][22] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA1P S2_6_34 ( .A(\CARRYB[5][34] ), .B(n430), .CI(\SUMB[5][35] ), .CO(
        \CARRYB[6][34] ), .S(\SUMB[6][34] ) );
  FA1 S2_34_15 ( .A(\ab[34][15] ), .B(\CARRYB[33][15] ), .CI(\SUMB[33][16] ), 
        .CO(\CARRYB[34][15] ), .S(\SUMB[34][15] ) );
  FA1A S2_39_11 ( .A(\ab[39][11] ), .B(\CARRYB[38][11] ), .CI(\SUMB[38][12] ), 
        .CO(\CARRYB[39][11] ), .S(\SUMB[39][11] ) );
  FA1A S2_39_12 ( .A(\CARRYB[38][12] ), .B(\ab[39][12] ), .CI(\SUMB[38][13] ), 
        .CO(\CARRYB[39][12] ), .S(\SUMB[39][12] ) );
  FA1A S2_37_12 ( .A(\ab[37][12] ), .B(\CARRYB[36][12] ), .CI(\SUMB[36][13] ), 
        .CO(\CARRYB[37][12] ), .S(\SUMB[37][12] ) );
  FA1P S2_9_18 ( .A(n528), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), .CO(
        \CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1AP S2_30_11 ( .A(n550), .B(\CARRYB[29][11] ), .CI(\SUMB[29][12] ), .CO(
        \CARRYB[30][11] ), .S(\SUMB[30][11] ) );
  FA1P S2_12_18 ( .A(n599), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), .CO(
        \CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA1P S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA1P S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA1P S2_45_39 ( .A(\ab[45][39] ), .B(\CARRYB[44][39] ), .CI(\SUMB[44][40] ), 
        .CO(\CARRYB[45][39] ), .S(\SUMB[45][39] ) );
  FA1A S2_34_16 ( .A(\ab[34][16] ), .B(\CARRYB[33][16] ), .CI(\SUMB[33][17] ), 
        .CO(\CARRYB[34][16] ), .S(\SUMB[34][16] ) );
  FA1AP S2_32_17 ( .A(\ab[32][17] ), .B(\CARRYB[31][17] ), .CI(\SUMB[31][18] ), 
        .CO(\CARRYB[32][17] ), .S(\SUMB[32][17] ) );
  FA1 S2_32_16 ( .A(\ab[32][16] ), .B(\CARRYB[31][16] ), .CI(\SUMB[31][17] ), 
        .CO(\CARRYB[32][16] ), .S(\SUMB[32][16] ) );
  FA1P S2_10_19 ( .A(n560), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), .CO(
        \CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1P S2_8_18 ( .A(n506), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), .CO(
        \CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1 S2_15_35 ( .A(\ab[35][15] ), .B(\CARRYB[14][35] ), .CI(\SUMB[14][36] ), 
        .CO(\CARRYB[15][35] ), .S(\SUMB[15][35] ) );
  FA1P S2_44_36 ( .A(\ab[44][36] ), .B(\CARRYB[43][36] ), .CI(\SUMB[43][37] ), 
        .CO(\CARRYB[44][36] ), .S(\SUMB[44][36] ) );
  FA1 S2_24_41 ( .A(\ab[41][24] ), .B(\CARRYB[23][41] ), .CI(\SUMB[23][42] ), 
        .CO(\CARRYB[24][41] ), .S(\SUMB[24][41] ) );
  FA1 S2_28_41 ( .A(\ab[41][28] ), .B(\CARRYB[27][41] ), .CI(\SUMB[27][42] ), 
        .CO(\CARRYB[28][41] ), .S(\SUMB[28][41] ) );
  FA1P S2_27_41 ( .A(\ab[41][27] ), .B(\CARRYB[26][41] ), .CI(\SUMB[26][42] ), 
        .CO(\CARRYB[27][41] ), .S(\SUMB[27][41] ) );
  FA1A S2_24_4 ( .A(n1272), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), .CO(
        \CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA1P S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA1A S2_15_20 ( .A(\ab[20][15] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA1P S2_2_30 ( .A(n290), .B(\CARRYB[1][30] ), .CI(\SUMB[1][31] ), .CO(
        \CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  FA1P S2_26_10 ( .A(n544), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), .CO(
        \CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA1P S2_15_13 ( .A(n628), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), .CO(
        \CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA1P S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA1P S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA1 S2_25_33 ( .A(\CARRYB[24][33] ), .B(\ab[33][25] ), .CI(\SUMB[24][34] ), 
        .CO(\CARRYB[25][33] ), .S(\SUMB[25][33] ) );
  FA1P S2_9_30 ( .A(n462), .B(\CARRYB[8][30] ), .CI(\SUMB[8][31] ), .CO(
        \CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA1 S2_32_15 ( .A(\SUMB[31][16] ), .B(\CARRYB[31][15] ), .CI(\ab[32][15] ), 
        .CO(\CARRYB[32][15] ), .S(\SUMB[32][15] ) );
  FA1 S2_4_28 ( .A(\CARRYB[3][28] ), .B(n351), .CI(\SUMB[3][29] ), .CO(
        \CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA1P S2_3_34 ( .A(n305), .B(\CARRYB[2][34] ), .CI(\SUMB[2][35] ), .CO(
        \CARRYB[3][34] ), .S(\SUMB[3][34] ) );
  FA1 S2_4_34 ( .A(n352), .B(\CARRYB[3][34] ), .CI(\SUMB[3][35] ), .CO(
        \CARRYB[4][34] ), .S(\SUMB[4][34] ) );
  FA1A S2_5_34 ( .A(n392), .B(\CARRYB[4][34] ), .CI(\SUMB[4][35] ), .CO(
        \CARRYB[5][34] ), .S(\SUMB[5][34] ) );
  FA1 S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA1 S2_36_13 ( .A(\CARRYB[35][13] ), .B(\ab[36][13] ), .CI(\SUMB[35][14] ), 
        .CO(\CARRYB[36][13] ), .S(\SUMB[36][13] ) );
  FA1AP S2_18_26 ( .A(\ab[26][18] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA1 S2_24_14 ( .A(n640), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), .CO(
        \CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA1P S2_17_41 ( .A(\ab[41][17] ), .B(\CARRYB[16][41] ), .CI(\SUMB[16][42] ), 
        .CO(\CARRYB[17][41] ), .S(\SUMB[17][41] ) );
  FA1P S2_36_31 ( .A(\ab[36][31] ), .B(\CARRYB[35][31] ), .CI(\SUMB[35][32] ), 
        .CO(\CARRYB[36][31] ), .S(\SUMB[36][31] ) );
  FA1P S2_14_14 ( .A(n1459), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), .CO(
        \CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1AP S2_29_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA1 S2_6_27 ( .A(\CARRYB[5][27] ), .B(n397), .CI(\SUMB[5][28] ), .CO(
        \CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA1 S2_10_27 ( .A(\CARRYB[9][27] ), .B(n520), .CI(\SUMB[9][28] ), .CO(
        \CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA1P S2_6_19 ( .A(n1289), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), .CO(
        \CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1P S2_19_21 ( .A(\ab[21][19] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA1P S2_22_36 ( .A(\CARRYB[21][36] ), .B(\ab[36][22] ), .CI(\SUMB[21][37] ), 
        .CO(\CARRYB[22][36] ), .S(\SUMB[22][36] ) );
  FA1AP S2_3_24 ( .A(\CARRYB[2][24] ), .B(n307), .CI(\SUMB[2][25] ), .CO(
        \CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA1 S2_34_1 ( .A(n1359), .B(\CARRYB[33][1] ), .CI(\SUMB[33][2] ), .CO(
        \CARRYB[34][1] ), .S(\SUMB[34][1] ) );
  FA1 S2_10_41 ( .A(\ab[41][10] ), .B(\CARRYB[9][41] ), .CI(\SUMB[9][42] ), 
        .CO(\CARRYB[10][41] ), .S(\SUMB[10][41] ) );
  FA1AP S2_3_35 ( .A(\CARRYB[2][35] ), .B(n298), .CI(\SUMB[2][36] ), .CO(
        \CARRYB[3][35] ), .S(\SUMB[3][35] ) );
  FA1 S2_2_35 ( .A(n1316), .B(\CARRYB[1][35] ), .CI(\SUMB[1][36] ), .CO(
        \CARRYB[2][35] ), .S(\SUMB[2][35] ) );
  FA1 S2_2_29 ( .A(\CARRYB[1][29] ), .B(n1303), .CI(\SUMB[1][30] ), .CO(
        \CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA1P S2_5_22 ( .A(\CARRYB[4][22] ), .B(n371), .CI(\SUMB[4][23] ), .CO(
        \CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA1P S2_5_37 ( .A(n1281), .B(\CARRYB[4][37] ), .CI(\SUMB[4][38] ), .CO(
        \CARRYB[5][37] ), .S(\SUMB[5][37] ) );
  FA1P S2_10_24 ( .A(n554), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), .CO(
        \CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA1 S2_10_21 ( .A(n547), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), .CO(
        \CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA1A S2_26_27 ( .A(\ab[27][26] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), 
        .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FA1P S2_3_19 ( .A(n329), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), .CO(
        \CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1 S2_12_31 ( .A(n591), .B(\CARRYB[11][31] ), .CI(\SUMB[11][32] ), .CO(
        \CARRYB[12][31] ), .S(\SUMB[12][31] ) );
  FA1A S2_4_38 ( .A(n335), .B(\CARRYB[3][38] ), .CI(\SUMB[3][39] ), .CO(
        \CARRYB[4][38] ), .S(\SUMB[4][38] ) );
  FA1 S2_9_31 ( .A(n524), .B(\CARRYB[8][31] ), .CI(\SUMB[8][32] ), .CO(
        \CARRYB[9][31] ), .S(\SUMB[9][31] ) );
  FA1 S2_9_6 ( .A(n449), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1P S2_10_6 ( .A(n464), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1P S2_9_23 ( .A(\CARRYB[8][23] ), .B(n521), .CI(\SUMB[8][24] ), .CO(
        \CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA1A S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA1P S2_18_30 ( .A(\ab[30][18] ), .B(\CARRYB[17][30] ), .CI(\SUMB[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA1P S2_7_35 ( .A(n417), .B(\CARRYB[6][35] ), .CI(\SUMB[6][36] ), .CO(
        \CARRYB[7][35] ), .S(\SUMB[7][35] ) );
  FA1A S2_12_13 ( .A(n604), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), .CO(
        \CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_2_39 ( .A(n1313), .B(\CARRYB[1][39] ), .CI(\SUMB[1][40] ), .CO(
        \CARRYB[2][39] ), .S(\SUMB[2][39] ) );
  FA1A S2_9_27 ( .A(n491), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), .CO(
        \CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA1A S2_29_30 ( .A(\ab[30][29] ), .B(\CARRYB[28][30] ), .CI(\SUMB[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FA1P S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA1A S2_12_19 ( .A(n605), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), .CO(
        \CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA1P S2_10_20 ( .A(n549), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), .CO(
        \CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1 S2_11_13 ( .A(n587), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), .CO(
        \CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_7_27 ( .A(\CARRYB[6][27] ), .B(n423), .CI(\SUMB[6][28] ), .CO(
        \CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA1A S2_11_21 ( .A(n580), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), .CO(
        \CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA1 S2_5_27 ( .A(n374), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), .CO(
        \CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA1P S2_8_34 ( .A(n488), .B(\CARRYB[7][34] ), .CI(\SUMB[7][35] ), .CO(
        \CARRYB[8][34] ), .S(\SUMB[8][34] ) );
  FA1 S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA1 S2_23_28 ( .A(\ab[28][23] ), .B(\CARRYB[22][28] ), .CI(\SUMB[22][29] ), 
        .CO(\CARRYB[23][28] ), .S(\SUMB[23][28] ) );
  FA1 S2_3_28 ( .A(n286), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), .CO(
        \CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA1P S2_41_22 ( .A(\ab[41][22] ), .B(\CARRYB[40][22] ), .CI(\SUMB[40][23] ), 
        .CO(\CARRYB[41][22] ), .S(\SUMB[41][22] ) );
  FA1A S2_29_2 ( .A(n1303), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), .CO(
        \CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA1P S2_10_35 ( .A(n532), .B(\CARRYB[9][35] ), .CI(\SUMB[9][36] ), .CO(
        \CARRYB[10][35] ), .S(\SUMB[10][35] ) );
  FA1P S2_41_33 ( .A(\ab[41][33] ), .B(\CARRYB[40][33] ), .CI(\SUMB[40][34] ), 
        .CO(\CARRYB[41][33] ), .S(\SUMB[41][33] ) );
  FA1A S2_14_18 ( .A(n644), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), .CO(
        \CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA1P S2_8_21 ( .A(n490), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), .CO(
        \CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA1A S2_30_3 ( .A(n300), .B(\CARRYB[29][3] ), .CI(\SUMB[29][4] ), .CO(
        \CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA1A S2_23_14 ( .A(n642), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), .CO(
        \CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA1P S2_26_13 ( .A(n616), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), .CO(
        \CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA1 S2_46_15 ( .A(\ab[46][15] ), .B(\CARRYB[45][15] ), .CI(\SUMB[45][16] ), 
        .CO(\CARRYB[46][15] ), .S(\SUMB[46][15] ) );
  FA1P S2_20_29 ( .A(\ab[29][20] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA1 S2_32_29 ( .A(\ab[32][29] ), .B(\CARRYB[31][29] ), .CI(\SUMB[31][30] ), 
        .CO(\CARRYB[32][29] ), .S(\SUMB[32][29] ) );
  FA1AP S2_8_20 ( .A(n478), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), .CO(
        \CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA1AP S2_8_26 ( .A(n497), .B(\SUMB[7][27] ), .CI(\CARRYB[7][26] ), .CO(
        \CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA1AP S2_24_28 ( .A(\ab[28][24] ), .B(\CARRYB[23][28] ), .CI(\SUMB[23][29] ), 
        .CO(\CARRYB[24][28] ), .S(\SUMB[24][28] ) );
  FA1 S2_29_11 ( .A(n571), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), .CO(
        \CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA1AP S2_26_31 ( .A(\ab[31][26] ), .B(\CARRYB[25][31] ), .CI(\SUMB[25][32] ), 
        .CO(\CARRYB[26][31] ), .S(\SUMB[26][31] ) );
  FA1A S2_28_30 ( .A(\ab[30][28] ), .B(\CARRYB[27][30] ), .CI(\SUMB[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA1P S2_16_39 ( .A(\ab[39][16] ), .B(\CARRYB[15][39] ), .CI(\SUMB[15][40] ), 
        .CO(\CARRYB[16][39] ), .S(\SUMB[16][39] ) );
  FA1P S2_22_37 ( .A(\ab[37][22] ), .B(\CARRYB[21][37] ), .CI(\SUMB[21][38] ), 
        .CO(\CARRYB[22][37] ), .S(\SUMB[22][37] ) );
  FA1P S2_23_37 ( .A(\ab[37][23] ), .B(\CARRYB[22][37] ), .CI(\SUMB[22][38] ), 
        .CO(\CARRYB[23][37] ), .S(\SUMB[23][37] ) );
  FA1P S2_29_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA1A S2_22_29 ( .A(\ab[29][22] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA1P S2_24_38 ( .A(\ab[38][24] ), .B(\CARRYB[23][38] ), .CI(\SUMB[23][39] ), 
        .CO(\CARRYB[24][38] ), .S(\SUMB[24][38] ) );
  FA1P S2_44_32 ( .A(\ab[44][32] ), .B(\CARRYB[43][32] ), .CI(\SUMB[43][33] ), 
        .CO(\CARRYB[44][32] ), .S(\SUMB[44][32] ) );
  FA1 S2_33_36 ( .A(\ab[36][33] ), .B(\CARRYB[32][36] ), .CI(\SUMB[32][37] ), 
        .CO(\CARRYB[33][36] ), .S(\SUMB[33][36] ) );
  FA1 S2_25_27 ( .A(\ab[27][25] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA1 S2_22_15 ( .A(\CARRYB[21][15] ), .B(\ab[22][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA1A S2_25_26 ( .A(\ab[26][25] ), .B(\CARRYB[24][26] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA1P S2_28_11 ( .A(n562), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), .CO(
        \CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA1AP S2_12_36 ( .A(\ab[36][12] ), .B(\CARRYB[11][36] ), .CI(\SUMB[11][37] ), 
        .CO(\CARRYB[12][36] ), .S(\SUMB[12][36] ) );
  FA1 S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA1 S2_3_42 ( .A(n1380), .B(\CARRYB[2][42] ), .CI(\SUMB[2][43] ), .CO(
        \CARRYB[3][42] ), .S(\SUMB[3][42] ) );
  FA1A S2_4_42 ( .A(\CARRYB[3][42] ), .B(n322), .CI(\SUMB[3][43] ), .CO(
        \CARRYB[4][42] ), .S(\SUMB[4][42] ) );
  FA1A S2_3_20 ( .A(n1379), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), .CO(
        \CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1 S2_7_39 ( .A(n475), .B(\CARRYB[6][39] ), .CI(\SUMB[6][40] ), .CO(
        \CARRYB[7][39] ), .S(\SUMB[7][39] ) );
  FA1A S2_38_15 ( .A(\ab[38][15] ), .B(\CARRYB[37][15] ), .CI(\SUMB[37][16] ), 
        .CO(\CARRYB[38][15] ), .S(\SUMB[38][15] ) );
  FA1A S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA1AP S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), 
        .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FA1 S2_31_17 ( .A(\ab[31][17] ), .B(\CARRYB[30][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FA1 S2_2_16 ( .A(n1299), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), .CO(
        \CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1P S2_13_37 ( .A(\ab[37][13] ), .B(\CARRYB[12][37] ), .CI(\SUMB[12][38] ), 
        .CO(\CARRYB[13][37] ), .S(\SUMB[13][37] ) );
  FA1A S2_34_17 ( .A(\ab[34][17] ), .B(\CARRYB[33][17] ), .CI(\SUMB[33][18] ), 
        .CO(\CARRYB[34][17] ), .S(\SUMB[34][17] ) );
  FA1 S2_33_17 ( .A(\ab[33][17] ), .B(\CARRYB[32][17] ), .CI(\SUMB[32][18] ), 
        .CO(\CARRYB[33][17] ), .S(\SUMB[33][17] ) );
  FA1AP S2_24_22 ( .A(\ab[24][22] ), .B(\CARRYB[23][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA1A S1_6_0 ( .A(n1387), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_16_0 ( .A(n1395), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), .CO(
        \CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S1_19_0 ( .A(n1334), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), .CO(
        \CARRYB[19][0] ), .S(\A1[17] ) );
  FA1A S1_21_0 ( .A(n651), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), .CO(
        \CARRYB[21][0] ), .S(\A1[19] ) );
  FA1A S2_6_1 ( .A(n1383), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_14_1 ( .A(n1376), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(
        \CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_17_2 ( .A(n294), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), .CO(
        \CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1A S2_20_1 ( .A(n1414), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), .CO(
        \CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1A S2_13_2 ( .A(n317), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), .CO(
        \CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_18_2 ( .A(n1339), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), .CO(
        \CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1A S2_19_2 ( .A(n291), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), .CO(
        \CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1A S2_21_4 ( .A(n363), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), .CO(
        \CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1A S4_36 ( .A(\ab[47][36] ), .B(\CARRYB[46][36] ), .CI(\SUMB[46][37] ), 
        .CO(\CARRYB[47][36] ), .S(\SUMB[47][36] ) );
  FA1A S4_40 ( .A(\ab[47][40] ), .B(\CARRYB[46][40] ), .CI(\SUMB[46][41] ), 
        .CO(\CARRYB[47][40] ), .S(\SUMB[47][40] ) );
  FA1A S4_26 ( .A(\ab[47][26] ), .B(\CARRYB[46][26] ), .CI(\SUMB[46][27] ), 
        .CO(\CARRYB[47][26] ), .S(\SUMB[47][26] ) );
  FA1A S3_46_46 ( .A(n1525), .B(\CARRYB[45][46] ), .CI(\ab[47][45] ), .CO(
        \CARRYB[46][46] ), .S(\SUMB[46][46] ) );
  FA1A S4_41 ( .A(\ab[47][41] ), .B(\CARRYB[46][41] ), .CI(\SUMB[46][42] ), 
        .CO(\CARRYB[47][41] ), .S(\SUMB[47][41] ) );
  FA1A S4_31 ( .A(\ab[47][31] ), .B(\CARRYB[46][31] ), .CI(\SUMB[46][32] ), 
        .CO(\CARRYB[47][31] ), .S(\SUMB[47][31] ) );
  FA1A S2_46_38 ( .A(\ab[46][38] ), .B(\CARRYB[45][38] ), .CI(\SUMB[45][39] ), 
        .CO(\CARRYB[46][38] ), .S(\SUMB[46][38] ) );
  FA1A S2_46_33 ( .A(\ab[46][33] ), .B(\CARRYB[45][33] ), .CI(\SUMB[45][34] ), 
        .CO(\CARRYB[46][33] ), .S(\SUMB[46][33] ) );
  FA1A S2_46_40 ( .A(\ab[46][40] ), .B(\CARRYB[45][40] ), .CI(\SUMB[45][41] ), 
        .CO(\CARRYB[46][40] ), .S(\SUMB[46][40] ) );
  FA1A S2_46_41 ( .A(\ab[46][41] ), .B(\CARRYB[45][41] ), .CI(\SUMB[45][42] ), 
        .CO(\CARRYB[46][41] ), .S(\SUMB[46][41] ) );
  FA1A S2_46_26 ( .A(\ab[46][26] ), .B(\CARRYB[45][26] ), .CI(\SUMB[45][27] ), 
        .CO(\CARRYB[46][26] ), .S(\SUMB[46][26] ) );
  FA1A S2_4_5 ( .A(n379), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_4_6 ( .A(n315), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_11_5 ( .A(n412), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(
        \CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_17_7 ( .A(n448), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), .CO(
        \CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1A S2_18_7 ( .A(n474), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), .CO(
        \CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1A S2_21_5 ( .A(n400), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), .CO(
        \CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1A S2_23_4 ( .A(n311), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), .CO(
        \CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA1A S2_29_4 ( .A(n1271), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), .CO(
        \CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA1A S2_45_14 ( .A(\ab[45][14] ), .B(\CARRYB[44][14] ), .CI(\SUMB[44][15] ), 
        .CO(\CARRYB[45][14] ), .S(\SUMB[45][14] ) );
  FA1A S2_45_33 ( .A(\ab[45][33] ), .B(\CARRYB[44][33] ), .CI(\SUMB[44][34] ), 
        .CO(\CARRYB[45][33] ), .S(\SUMB[45][33] ) );
  FA1A S2_45_40 ( .A(\ab[45][40] ), .B(\CARRYB[44][40] ), .CI(\SUMB[44][41] ), 
        .CO(\CARRYB[45][40] ), .S(\SUMB[45][40] ) );
  FA1A S2_45_41 ( .A(\ab[45][41] ), .B(\CARRYB[44][41] ), .CI(\SUMB[44][42] ), 
        .CO(\CARRYB[45][41] ), .S(\SUMB[45][41] ) );
  FA1A S2_45_45 ( .A(n1523), .B(\CARRYB[44][45] ), .CI(\SUMB[44][46] ), .CO(
        \CARRYB[45][45] ), .S(\SUMB[45][45] ) );
  FA1A S2_6_5 ( .A(n410), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_20_6 ( .A(n429), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), .CO(
        \CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1A S2_24_5 ( .A(n1275), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), .CO(
        \CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA1A S2_25_7 ( .A(n419), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), .CO(
        \CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA1A S2_28_6 ( .A(n396), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), .CO(
        \CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA1A S2_44_33 ( .A(\ab[44][33] ), .B(\CARRYB[43][33] ), .CI(\SUMB[43][34] ), 
        .CO(\CARRYB[44][33] ), .S(\SUMB[44][33] ) );
  FA1A S2_44_35 ( .A(\ab[44][35] ), .B(\CARRYB[43][35] ), .CI(\SUMB[43][36] ), 
        .CO(\CARRYB[44][35] ), .S(\SUMB[44][35] ) );
  FA1A S2_44_34 ( .A(\ab[44][34] ), .B(\CARRYB[43][34] ), .CI(\SUMB[43][35] ), 
        .CO(\CARRYB[44][34] ), .S(\SUMB[44][34] ) );
  FA1A S2_44_42 ( .A(\ab[44][42] ), .B(\CARRYB[43][42] ), .CI(\SUMB[43][43] ), 
        .CO(\CARRYB[44][42] ), .S(\SUMB[44][42] ) );
  FA1A S2_2_8 ( .A(n340), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_9_7 ( .A(n514), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_14_8 ( .A(n495), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), .CO(
        \CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_22_6 ( .A(n408), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), .CO(
        \CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA1A S2_23_6 ( .A(n422), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), .CO(
        \CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA1A S2_23_7 ( .A(n466), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), .CO(
        \CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA1A S2_43_34 ( .A(\ab[43][34] ), .B(\CARRYB[42][34] ), .CI(\SUMB[42][35] ), 
        .CO(\CARRYB[43][34] ), .S(\SUMB[43][34] ) );
  FA1A S2_43_38 ( .A(\ab[43][38] ), .B(\CARRYB[42][38] ), .CI(\SUMB[42][39] ), 
        .CO(\CARRYB[43][38] ), .S(\SUMB[43][38] ) );
  FA1A S2_43_36 ( .A(\ab[43][36] ), .B(\CARRYB[42][36] ), .CI(\SUMB[42][37] ), 
        .CO(\CARRYB[43][36] ), .S(\SUMB[43][36] ) );
  FA1A S2_43_35 ( .A(\ab[43][35] ), .B(\CARRYB[42][35] ), .CI(\SUMB[42][36] ), 
        .CO(\CARRYB[43][35] ), .S(\SUMB[43][35] ) );
  FA1A S3_42_46 ( .A(\ab[46][42] ), .B(\CARRYB[41][46] ), .CI(\ab[47][41] ), 
        .CO(\CARRYB[42][46] ), .S(\SUMB[42][46] ) );
  FA1A S2_21_8 ( .A(n490), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), .CO(
        \CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1A S2_22_8 ( .A(n452), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), .CO(
        \CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA1A S2_43_9 ( .A(\ab[9][43] ), .B(\CARRYB[42][9] ), .CI(\SUMB[42][10] ), 
        .CO(\CARRYB[43][9] ), .S(\SUMB[43][9] ) );
  FA1A S2_42_35 ( .A(\ab[42][35] ), .B(\CARRYB[41][35] ), .CI(\SUMB[41][36] ), 
        .CO(\CARRYB[42][35] ), .S(\SUMB[42][35] ) );
  FA1A S2_42_38 ( .A(\ab[42][38] ), .B(\CARRYB[41][38] ), .CI(\SUMB[41][39] ), 
        .CO(\CARRYB[42][38] ), .S(\SUMB[42][38] ) );
  FA1A S2_42_37 ( .A(\ab[42][37] ), .B(\CARRYB[41][37] ), .CI(\SUMB[41][38] ), 
        .CO(\CARRYB[42][37] ), .S(\SUMB[42][37] ) );
  FA1A S2_42_36 ( .A(\ab[42][36] ), .B(\CARRYB[41][36] ), .CI(\SUMB[41][37] ), 
        .CO(\CARRYB[42][36] ), .S(\SUMB[42][36] ) );
  FA1A S2_41_35 ( .A(\ab[41][35] ), .B(\CARRYB[40][35] ), .CI(\SUMB[40][36] ), 
        .CO(\CARRYB[41][35] ), .S(\SUMB[41][35] ) );
  FA1A S3_41_46 ( .A(\ab[46][41] ), .B(\CARRYB[40][46] ), .CI(\ab[47][40] ), 
        .CO(\CARRYB[41][46] ), .S(\SUMB[41][46] ) );
  FA1A S2_4_9 ( .A(n375), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_14_11 ( .A(n586), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), .CO(
        \CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_41_36 ( .A(\ab[41][36] ), .B(\CARRYB[40][36] ), .CI(\SUMB[40][37] ), 
        .CO(\CARRYB[41][36] ), .S(\SUMB[41][36] ) );
  FA1A S2_40_20 ( .A(\ab[40][20] ), .B(\CARRYB[39][20] ), .CI(\SUMB[39][21] ), 
        .CO(\CARRYB[40][20] ), .S(\SUMB[40][20] ) );
  FA1A S2_41_39 ( .A(\ab[41][39] ), .B(\CARRYB[40][39] ), .CI(\SUMB[40][40] ), 
        .CO(\CARRYB[41][39] ), .S(\SUMB[41][39] ) );
  FA1A S2_41_21 ( .A(\ab[41][21] ), .B(\CARRYB[40][21] ), .CI(\SUMB[40][22] ), 
        .CO(\CARRYB[41][21] ), .S(\SUMB[41][21] ) );
  FA1A S2_2_9 ( .A(n316), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_10_11 ( .A(n575), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), .CO(
        \CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_12_11 ( .A(n602), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), .CO(
        \CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_40_37 ( .A(\ab[40][37] ), .B(\CARRYB[39][37] ), .CI(\SUMB[39][38] ), 
        .CO(\CARRYB[40][37] ), .S(\SUMB[40][37] ) );
  FA1A S2_40_40 ( .A(n1510), .B(\CARRYB[39][40] ), .CI(\SUMB[39][41] ), .CO(
        \CARRYB[40][40] ), .S(\SUMB[40][40] ) );
  FA1A S2_4_10 ( .A(n378), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), .CO(
        \CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_5_11 ( .A(n412), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), .CO(
        \CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_10_12 ( .A(n576), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), .CO(
        \CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_9_12 ( .A(n553), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), .CO(
        \CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_25_13 ( .A(n625), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), .CO(
        \CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA1A S2_39_41 ( .A(\ab[41][39] ), .B(\CARRYB[38][41] ), .CI(\SUMB[38][42] ), 
        .CO(\CARRYB[39][41] ), .S(\SUMB[39][41] ) );
  FA1A S2_38_40 ( .A(\ab[40][38] ), .B(\CARRYB[37][40] ), .CI(\SUMB[37][41] ), 
        .CO(\CARRYB[38][40] ), .S(\SUMB[38][40] ) );
  FA1A S2_37_40 ( .A(\ab[40][37] ), .B(\CARRYB[36][40] ), .CI(\SUMB[36][41] ), 
        .CO(\CARRYB[37][40] ), .S(\SUMB[37][40] ) );
  FA1A S2_37_39 ( .A(\ab[39][37] ), .B(\CARRYB[36][39] ), .CI(\SUMB[36][40] ), 
        .CO(\CARRYB[37][39] ), .S(\SUMB[37][39] ) );
  FA1A S2_4_12 ( .A(n380), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), .CO(
        \CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_16_11 ( .A(n589), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), .CO(
        \CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA1A S2_38_43 ( .A(\ab[43][38] ), .B(\CARRYB[37][43] ), .CI(\SUMB[37][44] ), 
        .CO(\CARRYB[38][43] ), .S(\SUMB[38][43] ) );
  FA1A S2_37_42 ( .A(\ab[42][37] ), .B(\CARRYB[36][42] ), .CI(\SUMB[36][43] ), 
        .CO(\CARRYB[37][42] ), .S(\SUMB[37][42] ) );
  FA1A S2_2_13 ( .A(n317), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), .CO(
        \CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S2_7_13 ( .A(n465), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), .CO(
        \CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_7_14 ( .A(n459), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_36_43 ( .A(\ab[43][36] ), .B(\CARRYB[35][43] ), .CI(\SUMB[35][44] ), 
        .CO(\CARRYB[36][43] ), .S(\SUMB[36][43] ) );
  FA1A S2_37_25 ( .A(\ab[37][25] ), .B(\CARRYB[36][25] ), .CI(\SUMB[36][26] ), 
        .CO(\CARRYB[37][25] ), .S(\SUMB[37][25] ) );
  FA1A S2_4_13 ( .A(n391), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), .CO(
        \CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_6_14 ( .A(n438), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_6_15 ( .A(n442), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), .CO(
        \CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_8_15 ( .A(n492), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), .CO(
        \CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_30_14 ( .A(\CARRYB[29][14] ), .B(\ab[30][14] ), .CI(\SUMB[29][15] ), 
        .CO(\CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FA1A S2_35_24 ( .A(\ab[35][24] ), .B(\CARRYB[34][24] ), .CI(\SUMB[34][25] ), 
        .CO(\CARRYB[35][24] ), .S(\SUMB[35][24] ) );
  FA1A S2_35_44 ( .A(\ab[44][35] ), .B(\CARRYB[34][44] ), .CI(\SUMB[34][45] ), 
        .CO(\CARRYB[35][44] ), .S(\SUMB[35][44] ) );
  FA1A S2_34_42 ( .A(\ab[42][34] ), .B(\CARRYB[33][42] ), .CI(\SUMB[33][43] ), 
        .CO(\CARRYB[34][42] ), .S(\SUMB[34][42] ) );
  FA1A S2_34_43 ( .A(\ab[43][34] ), .B(\CARRYB[33][43] ), .CI(\SUMB[33][44] ), 
        .CO(\CARRYB[34][43] ), .S(\SUMB[34][43] ) );
  FA1A S2_33_37 ( .A(\ab[37][33] ), .B(\CARRYB[32][37] ), .CI(\SUMB[32][38] ), 
        .CO(\CARRYB[33][37] ), .S(\SUMB[33][37] ) );
  FA1A S2_5_15 ( .A(n413), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), .CO(
        \CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_5_16 ( .A(n404), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), .CO(
        \CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA1A S2_7_16 ( .A(n479), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), .CO(
        \CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1A S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA1A S2_31_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FA1A S2_35_45 ( .A(\ab[45][35] ), .B(\CARRYB[34][45] ), .CI(\SUMB[34][46] ), 
        .CO(\CARRYB[35][45] ), .S(\SUMB[35][45] ) );
  FA1A S2_33_44 ( .A(\ab[44][33] ), .B(\CARRYB[32][44] ), .CI(\SUMB[32][45] ), 
        .CO(\CARRYB[33][44] ), .S(\SUMB[33][44] ) );
  FA1A S2_4_16 ( .A(n361), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), .CO(
        \CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA1A S2_32_43 ( .A(\ab[43][32] ), .B(\CARRYB[31][43] ), .CI(\SUMB[31][44] ), 
        .CO(\CARRYB[32][43] ), .S(\SUMB[32][43] ) );
  FA1A S2_32_45 ( .A(\ab[45][32] ), .B(\CARRYB[31][45] ), .CI(\SUMB[31][46] ), 
        .CO(\CARRYB[32][45] ), .S(\SUMB[32][45] ) );
  FA1A S2_3_17 ( .A(n333), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), .CO(
        \CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1A S2_31_45 ( .A(\ab[45][31] ), .B(\CARRYB[30][45] ), .CI(\SUMB[30][46] ), 
        .CO(\CARRYB[31][45] ), .S(\SUMB[31][45] ) );
  FA1A S2_31_44 ( .A(\ab[44][31] ), .B(\CARRYB[30][44] ), .CI(\SUMB[30][45] ), 
        .CO(\CARRYB[31][44] ), .S(\SUMB[31][44] ) );
  FA1A S2_31_43 ( .A(\ab[43][31] ), .B(\CARRYB[30][43] ), .CI(\SUMB[30][44] ), 
        .CO(\CARRYB[31][43] ), .S(\SUMB[31][43] ) );
  FA1A S2_30_43 ( .A(\ab[43][30] ), .B(\CARRYB[29][43] ), .CI(\SUMB[29][44] ), 
        .CO(\CARRYB[30][43] ), .S(\SUMB[30][43] ) );
  FA1A S2_2_18 ( .A(n1339), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), .CO(
        \CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1AP S2_2_19 ( .A(n291), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), .CO(
        \CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA1A S2_16_17 ( .A(\ab[17][16] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA1A S3_30_46 ( .A(\ab[46][30] ), .B(\CARRYB[29][46] ), .CI(\ab[47][29] ), 
        .CO(\CARRYB[30][46] ), .S(\SUMB[30][46] ) );
  FA1A S2_30_44 ( .A(\ab[44][30] ), .B(\CARRYB[29][44] ), .CI(\SUMB[29][45] ), 
        .CO(\CARRYB[30][44] ), .S(\SUMB[30][44] ) );
  FA1A S2_29_44 ( .A(\ab[44][29] ), .B(\CARRYB[28][44] ), .CI(\SUMB[28][45] ), 
        .CO(\CARRYB[29][44] ), .S(\SUMB[29][44] ) );
  FA1A S2_13_21 ( .A(n626), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), .CO(
        \CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA1A S3_29_46 ( .A(\ab[46][29] ), .B(\CARRYB[28][46] ), .CI(\ab[47][28] ), 
        .CO(\CARRYB[29][46] ), .S(\SUMB[29][46] ) );
  FA1A S2_28_45 ( .A(\ab[45][28] ), .B(\CARRYB[27][45] ), .CI(\SUMB[27][46] ), 
        .CO(\CARRYB[28][45] ), .S(\SUMB[28][45] ) );
  FA1A S2_28_44 ( .A(\ab[44][28] ), .B(\CARRYB[27][44] ), .CI(\SUMB[27][45] ), 
        .CO(\CARRYB[28][44] ), .S(\SUMB[28][44] ) );
  FA1A S2_28_42 ( .A(\ab[42][28] ), .B(\CARRYB[27][42] ), .CI(\SUMB[27][43] ), 
        .CO(\CARRYB[28][42] ), .S(\SUMB[28][42] ) );
  FA1A S2_13_24 ( .A(n631), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), .CO(
        \CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA1A S2_26_29 ( .A(\ab[29][26] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA1A S3_28_46 ( .A(\ab[46][28] ), .B(\CARRYB[27][46] ), .CI(\ab[47][27] ), 
        .CO(\CARRYB[28][46] ), .S(\SUMB[28][46] ) );
  FA1A S2_27_45 ( .A(\ab[45][27] ), .B(\CARRYB[26][45] ), .CI(\SUMB[26][46] ), 
        .CO(\CARRYB[27][45] ), .S(\SUMB[27][45] ) );
  FA1A S2_27_44 ( .A(\ab[44][27] ), .B(\CARRYB[26][44] ), .CI(\SUMB[26][45] ), 
        .CO(\CARRYB[27][44] ), .S(\SUMB[27][44] ) );
  FA1A S2_24_32 ( .A(\ab[32][24] ), .B(\CARRYB[23][32] ), .CI(\SUMB[23][33] ), 
        .CO(\CARRYB[24][32] ), .S(\SUMB[24][32] ) );
  FA1A S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA1A S3_26_46 ( .A(\ab[46][26] ), .B(\CARRYB[25][46] ), .CI(\ab[47][25] ), 
        .CO(\CARRYB[26][46] ), .S(\SUMB[26][46] ) );
  FA1A S2_26_45 ( .A(\ab[45][26] ), .B(\CARRYB[25][45] ), .CI(\SUMB[25][46] ), 
        .CO(\CARRYB[26][45] ), .S(\SUMB[26][45] ) );
  FA1A S2_24_30 ( .A(\ab[30][24] ), .B(\CARRYB[23][30] ), .CI(\SUMB[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA1A S3_25_46 ( .A(\ab[46][25] ), .B(\CARRYB[24][46] ), .CI(\ab[47][24] ), 
        .CO(\CARRYB[25][46] ), .S(\SUMB[25][46] ) );
  FA1A S3_24_46 ( .A(\ab[46][24] ), .B(\CARRYB[23][46] ), .CI(\ab[47][23] ), 
        .CO(\CARRYB[24][46] ), .S(\SUMB[24][46] ) );
  FA1A S2_23_24 ( .A(\ab[24][23] ), .B(\CARRYB[22][24] ), .CI(\SUMB[22][25] ), 
        .CO(\CARRYB[23][24] ), .S(\SUMB[23][24] ) );
  FA1A S3_23_46 ( .A(\ab[46][23] ), .B(\CARRYB[22][46] ), .CI(\ab[47][22] ), 
        .CO(\CARRYB[23][46] ), .S(\SUMB[23][46] ) );
  FA1A S2_21_37 ( .A(\ab[37][21] ), .B(\CARRYB[20][37] ), .CI(\SUMB[20][38] ), 
        .CO(\CARRYB[21][37] ), .S(\SUMB[21][37] ) );
  FA1A S2_11_27 ( .A(\CARRYB[10][27] ), .B(n543), .CI(\SUMB[10][28] ), .CO(
        \CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA1A S2_9_28 ( .A(n502), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), .CO(
        \CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA1A S2_18_27 ( .A(\ab[27][18] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA1A S3_22_46 ( .A(\ab[46][22] ), .B(\CARRYB[21][46] ), .CI(\ab[47][21] ), 
        .CO(\CARRYB[22][46] ), .S(\SUMB[22][46] ) );
  FA1A S2_23_41 ( .A(\ab[41][23] ), .B(\CARRYB[22][41] ), .CI(\SUMB[22][42] ), 
        .CO(\CARRYB[23][41] ), .S(\SUMB[23][41] ) );
  FA1A S2_10_28 ( .A(n548), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), .CO(
        \CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA1A S2_21_43 ( .A(\ab[43][21] ), .B(\CARRYB[20][43] ), .CI(\SUMB[20][44] ), 
        .CO(\CARRYB[21][43] ), .S(\SUMB[21][43] ) );
  FA1A S2_22_41 ( .A(\ab[41][22] ), .B(\CARRYB[21][41] ), .CI(\SUMB[21][42] ), 
        .CO(\CARRYB[22][41] ), .S(\SUMB[22][41] ) );
  FA1A S2_9_29 ( .A(n509), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), .CO(
        \CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA1A S2_20_43 ( .A(\ab[43][20] ), .B(\CARRYB[19][43] ), .CI(\SUMB[19][44] ), 
        .CO(\CARRYB[20][43] ), .S(\SUMB[20][43] ) );
  FA1A S2_4_31 ( .A(n365), .B(\CARRYB[3][31] ), .CI(\SUMB[3][32] ), .CO(
        \CARRYB[4][31] ), .S(\SUMB[4][31] ) );
  FA1A S2_14_33 ( .A(\ab[33][14] ), .B(\CARRYB[13][33] ), .CI(\SUMB[13][34] ), 
        .CO(\CARRYB[14][33] ), .S(\SUMB[14][33] ) );
  FA1A S2_2_32 ( .A(n1315), .B(\CARRYB[1][32] ), .CI(\SUMB[1][33] ), .CO(
        \CARRYB[2][32] ), .S(\SUMB[2][32] ) );
  FA1A S2_6_37 ( .A(n1286), .B(\CARRYB[5][37] ), .CI(\SUMB[5][38] ), .CO(
        \CARRYB[6][37] ), .S(\SUMB[6][37] ) );
  FA1A S2_36_1 ( .A(n1404), .B(\CARRYB[35][1] ), .CI(\SUMB[35][2] ), .CO(
        \CARRYB[36][1] ), .S(\SUMB[36][1] ) );
  FA1A S2_23_3 ( .A(n287), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), .CO(
        \CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA1A S2_11_3 ( .A(n331), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(
        \CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_19_5 ( .A(n1283), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), .CO(
        \CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1A S2_19_6 ( .A(n1289), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), .CO(
        \CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1A S2_32_3 ( .A(n321), .B(\CARRYB[31][3] ), .CI(\SUMB[31][4] ), .CO(
        \CARRYB[32][3] ), .S(\SUMB[32][3] ) );
  FA1A S2_38_36 ( .A(\ab[38][36] ), .B(\CARRYB[37][36] ), .CI(\SUMB[37][37] ), 
        .CO(\CARRYB[38][36] ), .S(\SUMB[38][36] ) );
  FA1A S2_27_31 ( .A(\ab[31][27] ), .B(\CARRYB[26][31] ), .CI(\SUMB[26][32] ), 
        .CO(\CARRYB[27][31] ), .S(\SUMB[27][31] ) );
  FA1A S2_26_44 ( .A(\ab[44][26] ), .B(\CARRYB[25][44] ), .CI(\SUMB[25][45] ), 
        .CO(\CARRYB[26][44] ), .S(\SUMB[26][44] ) );
  FA1A S2_22_33 ( .A(\ab[33][22] ), .B(\CARRYB[21][33] ), .CI(\SUMB[21][34] ), 
        .CO(\CARRYB[22][33] ), .S(\SUMB[22][33] ) );
  FA1A S2_4_25 ( .A(n357), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), .CO(
        \CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA1A S2_16_34 ( .A(\ab[34][16] ), .B(\CARRYB[15][34] ), .CI(\SUMB[15][35] ), 
        .CO(\CARRYB[16][34] ), .S(\SUMB[16][34] ) );
  FA1A S2_28_43 ( .A(\ab[43][28] ), .B(\CARRYB[27][43] ), .CI(\SUMB[27][44] ), 
        .CO(\CARRYB[28][43] ), .S(\SUMB[28][43] ) );
  FA1P S2_46_45 ( .A(\ab[46][45] ), .B(\CARRYB[45][45] ), .CI(\SUMB[45][46] ), 
        .CO(\CARRYB[46][45] ), .S(\SUMB[46][45] ) );
  FA1AP S4_45 ( .A(\ab[47][45] ), .B(\CARRYB[46][45] ), .CI(\SUMB[46][46] ), 
        .CO(\CARRYB[47][45] ), .S(\SUMB[47][45] ) );
  FA1AP S2_46_44 ( .A(\ab[46][44] ), .B(\CARRYB[45][44] ), .CI(\SUMB[45][45] ), 
        .CO(\CARRYB[46][44] ), .S(\SUMB[46][44] ) );
  FA1AP S4_44 ( .A(\ab[47][44] ), .B(\CARRYB[46][44] ), .CI(\SUMB[46][45] ), 
        .CO(\CARRYB[47][44] ), .S(\SUMB[47][44] ) );
  FA1P S2_12_45 ( .A(\ab[45][12] ), .B(\CARRYB[11][45] ), .CI(\SUMB[11][46] ), 
        .CO(\CARRYB[12][45] ), .S(\SUMB[12][45] ) );
  FA1 S3_44_46 ( .A(\ab[46][44] ), .B(\CARRYB[43][46] ), .CI(\ab[47][43] ), 
        .CO(\CARRYB[44][46] ), .S(\SUMB[44][46] ) );
  FA1P S3_45_46 ( .A(\ab[46][45] ), .B(\CARRYB[44][46] ), .CI(\ab[47][44] ), 
        .CO(\CARRYB[45][46] ), .S(\SUMB[45][46] ) );
  FA1P S2_39_8 ( .A(n482), .B(\CARRYB[38][8] ), .CI(\SUMB[38][9] ), .CO(
        \CARRYB[39][8] ), .S(\SUMB[39][8] ) );
  FA1P S2_10_45 ( .A(\ab[45][10] ), .B(\CARRYB[9][45] ), .CI(\SUMB[9][46] ), 
        .CO(\CARRYB[10][45] ), .S(\SUMB[10][45] ) );
  FA1P S2_11_45 ( .A(\ab[45][11] ), .B(\CARRYB[10][45] ), .CI(\SUMB[10][46] ), 
        .CO(\CARRYB[11][45] ), .S(\SUMB[11][45] ) );
  FA1P S3_10_46 ( .A(\ab[46][10] ), .B(\CARRYB[9][46] ), .CI(\ab[9][47] ), 
        .CO(\CARRYB[10][46] ), .S(\SUMB[10][46] ) );
  FA1P S3_11_46 ( .A(\ab[46][11] ), .B(\CARRYB[10][46] ), .CI(\ab[47][10] ), 
        .CO(\CARRYB[11][46] ), .S(\SUMB[11][46] ) );
  FA1P S2_33_7 ( .A(n445), .B(\CARRYB[32][7] ), .CI(\SUMB[32][8] ), .CO(
        \CARRYB[33][7] ), .S(\SUMB[33][7] ) );
  FA1P S2_27_9 ( .A(n491), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), .CO(
        \CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA1P S3_8_46 ( .A(\ab[8][46] ), .B(\CARRYB[7][46] ), .CI(\ab[7][47] ), .CO(
        \CARRYB[8][46] ), .S(\SUMB[8][46] ) );
  FA1P S3_9_46 ( .A(\ab[9][46] ), .B(\CARRYB[8][46] ), .CI(\ab[8][47] ), .CO(
        \CARRYB[9][46] ), .S(\SUMB[9][46] ) );
  FA1P S2_32_7 ( .A(n440), .B(\CARRYB[31][7] ), .CI(\SUMB[31][8] ), .CO(
        \CARRYB[32][7] ), .S(\SUMB[32][7] ) );
  FA1P S2_8_45 ( .A(\ab[8][45] ), .B(\CARRYB[7][45] ), .CI(\SUMB[7][46] ), 
        .CO(\CARRYB[8][45] ), .S(\SUMB[8][45] ) );
  FA1P S2_9_45 ( .A(\ab[9][45] ), .B(\CARRYB[8][45] ), .CI(\SUMB[8][46] ), 
        .CO(\CARRYB[9][45] ), .S(\SUMB[9][45] ) );
  FA1P S2_27_8 ( .A(n446), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), .CO(
        \CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA1P S2_24_9 ( .A(n513), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), .CO(
        \CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA1P S2_25_9 ( .A(n483), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), .CO(
        \CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA1AP S2_25_8 ( .A(n468), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), .CO(
        \CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA1P S2_26_8 ( .A(n497), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), .CO(
        \CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA1P S3_6_46 ( .A(n420), .B(\CARRYB[5][46] ), .CI(n274), .CO(\CARRYB[6][46] ), .S(\SUMB[6][46] ) );
  FA1P S3_7_46 ( .A(\ab[7][46] ), .B(\CARRYB[6][46] ), .CI(\ab[6][47] ), .CO(
        \CARRYB[7][46] ), .S(\SUMB[7][46] ) );
  FA1P S2_36_4 ( .A(n367), .B(\CARRYB[35][4] ), .CI(\SUMB[35][5] ), .CO(
        \CARRYB[36][4] ), .S(\SUMB[36][4] ) );
  FA1P S2_6_45 ( .A(n435), .B(\CARRYB[5][45] ), .CI(\SUMB[5][46] ), .CO(
        \CARRYB[6][45] ), .S(\SUMB[6][45] ) );
  FA1P S2_7_45 ( .A(n473), .B(\CARRYB[6][45] ), .CI(\SUMB[6][46] ), .CO(
        \CARRYB[7][45] ), .S(\SUMB[7][45] ) );
  FA1P S2_37_35 ( .A(\ab[37][35] ), .B(\CARRYB[36][35] ), .CI(\SUMB[36][36] ), 
        .CO(\CARRYB[37][35] ), .S(\SUMB[37][35] ) );
  FA1P S2_22_9 ( .A(n280), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), .CO(
        \CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA1P S2_23_9 ( .A(n521), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), .CO(
        \CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA1AP S2_19_9 ( .A(n531), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), .CO(
        \CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA1P S2_35_35 ( .A(n1500), .B(\CARRYB[34][35] ), .CI(\SUMB[34][36] ), .CO(
        \CARRYB[35][35] ), .S(\SUMB[35][35] ) );
  FA1P S2_36_35 ( .A(\ab[36][35] ), .B(\CARRYB[35][35] ), .CI(\SUMB[35][36] ), 
        .CO(\CARRYB[36][35] ), .S(\SUMB[36][35] ) );
  FA1 S2_18_8 ( .A(n506), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), .CO(
        \CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA1P S2_30_7 ( .A(n411), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), .CO(
        \CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA1 S2_20_8 ( .A(n478), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), .CO(
        \CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA1P S3_4_46 ( .A(n334), .B(\CARRYB[3][46] ), .CI(n270), .CO(\CARRYB[4][46] ), .S(\SUMB[4][46] ) );
  FA1P S3_5_46 ( .A(n388), .B(\CARRYB[4][46] ), .CI(n272), .CO(\CARRYB[5][46] ), .S(\SUMB[5][46] ) );
  FA1 S2_46_6 ( .A(n420), .B(\CARRYB[45][6] ), .CI(\SUMB[45][7] ), .CO(
        \CARRYB[46][6] ), .S(\SUMB[46][6] ) );
  FA1AP S4_6 ( .A(\ab[6][47] ), .B(\CARRYB[46][6] ), .CI(\SUMB[46][7] ), .CO(
        \CARRYB[47][6] ), .S(\SUMB[47][6] ) );
  FA1AP S2_39_36 ( .A(\ab[39][36] ), .B(\CARRYB[38][36] ), .CI(\SUMB[38][37] ), 
        .CO(\CARRYB[39][36] ), .S(\SUMB[39][36] ) );
  FA1 S2_40_35 ( .A(\ab[40][35] ), .B(\CARRYB[39][35] ), .CI(\SUMB[39][36] ), 
        .CO(\CARRYB[40][35] ), .S(\SUMB[40][35] ) );
  FA1A S2_39_34 ( .A(\ab[39][34] ), .B(\CARRYB[38][34] ), .CI(\SUMB[38][35] ), 
        .CO(\CARRYB[39][34] ), .S(\SUMB[39][34] ) );
  FA1P S2_33_38 ( .A(\ab[38][33] ), .B(\CARRYB[32][38] ), .CI(\SUMB[32][39] ), 
        .CO(\CARRYB[33][38] ), .S(\SUMB[33][38] ) );
  FA1 S2_27_5 ( .A(n374), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), .CO(
        \CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA1P S2_33_35 ( .A(\ab[35][33] ), .B(\CARRYB[32][35] ), .CI(\SUMB[32][36] ), 
        .CO(\CARRYB[33][35] ), .S(\SUMB[33][35] ) );
  FA1P S2_34_35 ( .A(\ab[35][34] ), .B(\CARRYB[33][35] ), .CI(\SUMB[33][36] ), 
        .CO(\CARRYB[34][35] ), .S(\SUMB[34][35] ) );
  FA1P S2_4_45 ( .A(n344), .B(\CARRYB[3][45] ), .CI(\SUMB[3][46] ), .CO(
        \CARRYB[4][45] ), .S(\SUMB[4][45] ) );
  FA1P S2_5_45 ( .A(n401), .B(\CARRYB[4][45] ), .CI(\SUMB[4][46] ), .CO(
        \CARRYB[5][45] ), .S(\SUMB[5][45] ) );
  FA1P S2_37_8 ( .A(n486), .B(\CARRYB[36][8] ), .CI(\SUMB[36][9] ), .CO(
        \CARRYB[37][8] ), .S(\SUMB[37][8] ) );
  FA1P S2_21_22 ( .A(\SUMB[20][23] ), .B(\CARRYB[20][22] ), .CI(\ab[22][21] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA1AP S2_38_38 ( .A(A[38]), .B(\CARRYB[37][38] ), .CI(\SUMB[37][39] ), .CO(
        \CARRYB[38][38] ), .S(\SUMB[38][38] ) );
  FA1P S2_35_39 ( .A(\ab[39][35] ), .B(\CARRYB[34][39] ), .CI(\SUMB[34][40] ), 
        .CO(\CARRYB[35][39] ), .S(\SUMB[35][39] ) );
  FA1P S2_36_39 ( .A(\ab[39][36] ), .B(\CARRYB[35][39] ), .CI(\SUMB[35][40] ), 
        .CO(\CARRYB[36][39] ), .S(\SUMB[36][39] ) );
  FA1AP S2_26_5 ( .A(n389), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), .CO(
        \CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA1P S2_38_37 ( .A(\ab[38][37] ), .B(\CARRYB[37][37] ), .CI(\SUMB[37][38] ), 
        .CO(\CARRYB[38][37] ), .S(\SUMB[38][37] ) );
  FA1P S2_39_37 ( .A(\ab[39][37] ), .B(\CARRYB[38][37] ), .CI(\SUMB[38][38] ), 
        .CO(\CARRYB[39][37] ), .S(\SUMB[39][37] ) );
  FA1P S2_33_39 ( .A(\ab[39][33] ), .B(\CARRYB[32][39] ), .CI(\SUMB[32][40] ), 
        .CO(\CARRYB[33][39] ), .S(\SUMB[33][39] ) );
  FA1AP S2_24_6 ( .A(n1282), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), .CO(
        \CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA1 S2_25_5 ( .A(n406), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), .CO(
        \CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA1 S2_31_38 ( .A(\ab[38][31] ), .B(\CARRYB[30][38] ), .CI(\SUMB[30][39] ), 
        .CO(\CARRYB[31][38] ), .S(\SUMB[31][38] ) );
  FA1P S2_16_44 ( .A(\ab[44][16] ), .B(\CARRYB[15][44] ), .CI(\SUMB[15][45] ), 
        .CO(\CARRYB[16][44] ), .S(\SUMB[16][44] ) );
  FA1P S2_44_6 ( .A(n273), .B(\CARRYB[43][6] ), .CI(\SUMB[43][7] ), .CO(
        \CARRYB[44][6] ), .S(\SUMB[44][6] ) );
  FA1P S2_45_6 ( .A(n435), .B(\CARRYB[44][6] ), .CI(\SUMB[44][7] ), .CO(
        \CARRYB[45][6] ), .S(\SUMB[45][6] ) );
  FA1P S2_31_6 ( .A(n453), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), .CO(
        \CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FA1A S2_34_36 ( .A(\ab[36][34] ), .B(\CARRYB[33][36] ), .CI(\SUMB[33][37] ), 
        .CO(\CARRYB[34][36] ), .S(\SUMB[34][36] ) );
  FA1P S2_34_34 ( .A(\ab[34][34] ), .B(\CARRYB[33][34] ), .CI(\SUMB[33][35] ), 
        .CO(\CARRYB[34][34] ), .S(\SUMB[34][34] ) );
  FA1P S2_35_34 ( .A(\ab[35][34] ), .B(\CARRYB[34][34] ), .CI(\SUMB[34][35] ), 
        .CO(\CARRYB[35][34] ), .S(\SUMB[35][34] ) );
  FA1P S2_17_6 ( .A(n1292), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), .CO(
        \CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1AP S2_32_37 ( .A(\ab[37][32] ), .B(\CARRYB[31][37] ), .CI(\SUMB[31][38] ), 
        .CO(\CARRYB[32][37] ), .S(\SUMB[32][37] ) );
  FA1 S2_27_6 ( .A(n397), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), .CO(
        \CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA1P S2_31_22 ( .A(\ab[31][22] ), .B(\CARRYB[30][22] ), .CI(\SUMB[30][23] ), 
        .CO(\CARRYB[31][22] ), .S(\SUMB[31][22] ) );
  FA1P S2_15_10 ( .A(n558), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), .CO(
        \CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1P S2_38_8 ( .A(n1293), .B(\CARRYB[37][8] ), .CI(\SUMB[37][9] ), .CO(
        \CARRYB[38][8] ), .S(\SUMB[38][8] ) );
  FA1P S2_35_9 ( .A(n496), .B(\CARRYB[34][9] ), .CI(\SUMB[34][10] ), .CO(
        \CARRYB[35][9] ), .S(\SUMB[35][9] ) );
  FA1P S2_36_9 ( .A(n537), .B(\CARRYB[35][9] ), .CI(\SUMB[35][10] ), .CO(
        \CARRYB[36][9] ), .S(\SUMB[36][9] ) );
  FA1P S2_25_43 ( .A(\ab[43][25] ), .B(\CARRYB[24][43] ), .CI(\SUMB[24][44] ), 
        .CO(\CARRYB[25][43] ), .S(\SUMB[25][43] ) );
  FA1P S2_26_43 ( .A(\ab[43][26] ), .B(\CARRYB[25][43] ), .CI(\SUMB[25][44] ), 
        .CO(\CARRYB[26][43] ), .S(\SUMB[26][43] ) );
  FA1P S2_15_45 ( .A(\ab[45][15] ), .B(\CARRYB[14][45] ), .CI(\SUMB[14][46] ), 
        .CO(\CARRYB[15][45] ), .S(\SUMB[15][45] ) );
  FA1P S2_16_45 ( .A(\ab[45][16] ), .B(\CARRYB[15][45] ), .CI(\SUMB[15][46] ), 
        .CO(\CARRYB[16][45] ), .S(\SUMB[16][45] ) );
  FA1P S2_31_36 ( .A(\ab[36][31] ), .B(\CARRYB[30][36] ), .CI(\SUMB[30][37] ), 
        .CO(\CARRYB[31][36] ), .S(\SUMB[31][36] ) );
  FA1P S2_34_10 ( .A(n564), .B(\CARRYB[33][10] ), .CI(\SUMB[33][11] ), .CO(
        \CARRYB[34][10] ), .S(\SUMB[34][10] ) );
  FA1P S2_14_44 ( .A(\ab[44][14] ), .B(\CARRYB[13][44] ), .CI(\SUMB[13][45] ), 
        .CO(\CARRYB[14][44] ), .S(\SUMB[14][44] ) );
  FA1P S2_15_44 ( .A(\ab[44][15] ), .B(\CARRYB[14][44] ), .CI(\SUMB[14][45] ), 
        .CO(\CARRYB[15][44] ), .S(\SUMB[15][44] ) );
  FA1AP S2_31_24 ( .A(\ab[31][24] ), .B(\CARRYB[30][24] ), .CI(\SUMB[30][25] ), 
        .CO(\CARRYB[31][24] ), .S(\SUMB[31][24] ) );
  FA1P S2_29_37 ( .A(\ab[37][29] ), .B(\CARRYB[28][37] ), .CI(\SUMB[28][38] ), 
        .CO(\CARRYB[29][37] ), .S(\SUMB[29][37] ) );
  FA1P S2_27_38 ( .A(\ab[38][27] ), .B(\CARRYB[26][38] ), .CI(\SUMB[26][39] ), 
        .CO(\CARRYB[27][38] ), .S(\SUMB[27][38] ) );
  FA1P S2_28_38 ( .A(\ab[38][28] ), .B(\CARRYB[27][38] ), .CI(\SUMB[27][39] ), 
        .CO(\CARRYB[28][38] ), .S(\SUMB[28][38] ) );
  FA1P S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA1P S2_30_22 ( .A(\ab[30][22] ), .B(\CARRYB[29][22] ), .CI(\SUMB[29][23] ), 
        .CO(\CARRYB[30][22] ), .S(\SUMB[30][22] ) );
  FA1P S2_32_21 ( .A(\ab[32][21] ), .B(\CARRYB[31][21] ), .CI(\SUMB[31][22] ), 
        .CO(\CARRYB[32][21] ), .S(\SUMB[32][21] ) );
  FA1P S2_31_35 ( .A(\ab[35][31] ), .B(\CARRYB[30][35] ), .CI(\SUMB[30][36] ), 
        .CO(\CARRYB[31][35] ), .S(\SUMB[31][35] ) );
  FA1P S2_32_35 ( .A(\ab[35][32] ), .B(\CARRYB[31][35] ), .CI(\SUMB[31][36] ), 
        .CO(\CARRYB[32][35] ), .S(\SUMB[32][35] ) );
  FA1P S2_26_25 ( .A(\ab[26][25] ), .B(\CARRYB[25][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA1P S2_31_10 ( .A(n545), .B(\CARRYB[30][10] ), .CI(\SUMB[30][11] ), .CO(
        \CARRYB[31][10] ), .S(\SUMB[31][10] ) );
  FA1 S2_22_4 ( .A(n313), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), .CO(
        \CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA1P S2_11_8 ( .A(n533), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(
        \CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1P S2_12_8 ( .A(n538), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), .CO(
        \CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1P S2_13_45 ( .A(\ab[45][13] ), .B(\CARRYB[12][45] ), .CI(\SUMB[12][46] ), 
        .CO(\CARRYB[13][45] ), .S(\SUMB[13][45] ) );
  FA1P S2_14_45 ( .A(\ab[45][14] ), .B(\CARRYB[13][45] ), .CI(\SUMB[13][46] ), 
        .CO(\CARRYB[14][45] ), .S(\SUMB[14][45] ) );
  FA1 S2_18_5 ( .A(n398), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), .CO(
        \CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1P S3_13_46 ( .A(\ab[46][13] ), .B(\CARRYB[12][46] ), .CI(\ab[47][12] ), 
        .CO(\CARRYB[13][46] ), .S(\SUMB[13][46] ) );
  FA1P S3_14_46 ( .A(\ab[46][14] ), .B(\CARRYB[13][46] ), .CI(\ab[47][13] ), 
        .CO(\CARRYB[14][46] ), .S(\SUMB[14][46] ) );
  FA1P S2_16_5 ( .A(n404), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), .CO(
        \CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1P S2_17_5 ( .A(n1284), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), .CO(
        \CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1P S2_31_39 ( .A(\ab[39][31] ), .B(\CARRYB[30][39] ), .CI(\SUMB[30][40] ), 
        .CO(\CARRYB[31][39] ), .S(\SUMB[31][39] ) );
  FA1P S2_32_39 ( .A(\ab[39][32] ), .B(\CARRYB[31][39] ), .CI(\SUMB[31][40] ), 
        .CO(\CARRYB[32][39] ), .S(\SUMB[32][39] ) );
  FA1P S2_30_37 ( .A(\ab[37][30] ), .B(\CARRYB[29][37] ), .CI(\SUMB[29][38] ), 
        .CO(\CARRYB[30][37] ), .S(\SUMB[30][37] ) );
  FA1P S2_8_4 ( .A(n372), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1P S2_9_4 ( .A(n375), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1P S2_37_33 ( .A(\ab[37][33] ), .B(\CARRYB[36][33] ), .CI(\SUMB[36][34] ), 
        .CO(\CARRYB[37][33] ), .S(\SUMB[37][33] ) );
  FA1P S2_38_33 ( .A(\ab[38][33] ), .B(\CARRYB[37][33] ), .CI(\SUMB[37][34] ), 
        .CO(\CARRYB[38][33] ), .S(\SUMB[38][33] ) );
  FA1P S1_35_0 ( .A(n1362), .B(\CARRYB[34][0] ), .CI(\SUMB[34][1] ), .CO(
        \CARRYB[35][0] ), .S(\A1[33] ) );
  FA1P S2_44_45 ( .A(\ab[45][44] ), .B(\CARRYB[43][45] ), .CI(\SUMB[43][46] ), 
        .CO(\CARRYB[44][45] ), .S(\SUMB[44][45] ) );
  FA1AP S2_45_44 ( .A(\ab[45][44] ), .B(\CARRYB[44][44] ), .CI(\SUMB[44][45] ), 
        .CO(\CARRYB[45][44] ), .S(\SUMB[45][44] ) );
  FA1P S2_32_34 ( .A(\ab[34][32] ), .B(\CARRYB[31][34] ), .CI(\SUMB[31][35] ), 
        .CO(\CARRYB[32][34] ), .S(\SUMB[32][34] ) );
  FA1P S2_33_34 ( .A(\ab[34][33] ), .B(\CARRYB[32][34] ), .CI(\SUMB[32][35] ), 
        .CO(\CARRYB[33][34] ), .S(\SUMB[33][34] ) );
  FA1AP S2_39_39 ( .A(n1507), .B(\CARRYB[38][39] ), .CI(\SUMB[38][40] ), .CO(
        \CARRYB[39][39] ), .S(\SUMB[39][39] ) );
  FA1AP S2_40_39 ( .A(\ab[40][39] ), .B(\CARRYB[39][39] ), .CI(\SUMB[39][40] ), 
        .CO(\CARRYB[40][39] ), .S(\SUMB[40][39] ) );
  FA1A S2_28_28 ( .A(n1487), .B(\CARRYB[27][28] ), .CI(\SUMB[27][29] ), .CO(
        \CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA1AP S2_29_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA1P S2_25_29 ( .A(\ab[29][25] ), .B(\CARRYB[24][29] ), .CI(\SUMB[24][30] ), 
        .CO(\CARRYB[25][29] ), .S(\SUMB[25][29] ) );
  FA1 S2_46_43 ( .A(\ab[46][43] ), .B(\CARRYB[45][43] ), .CI(\SUMB[45][44] ), 
        .CO(\CARRYB[46][43] ), .S(\SUMB[46][43] ) );
  FA1AP S4_43 ( .A(\ab[47][43] ), .B(\CARRYB[46][43] ), .CI(\SUMB[46][44] ), 
        .CO(\CARRYB[47][43] ), .S(\SUMB[47][43] ) );
  FA1P S2_27_23 ( .A(\ab[27][23] ), .B(\CARRYB[26][23] ), .CI(\SUMB[26][24] ), 
        .CO(\CARRYB[27][23] ), .S(\SUMB[27][23] ) );
  FA1P S2_41_40 ( .A(\ab[41][40] ), .B(\CARRYB[40][40] ), .CI(\SUMB[40][41] ), 
        .CO(\CARRYB[41][40] ), .S(\SUMB[41][40] ) );
  FA1P S2_42_40 ( .A(\ab[42][40] ), .B(\CARRYB[41][40] ), .CI(\SUMB[41][41] ), 
        .CO(\CARRYB[42][40] ), .S(\SUMB[42][40] ) );
  FA1P S2_44_14 ( .A(\ab[44][14] ), .B(\CARRYB[43][14] ), .CI(\SUMB[43][15] ), 
        .CO(\CARRYB[44][14] ), .S(\SUMB[44][14] ) );
  FA1P S2_29_22 ( .A(\ab[29][22] ), .B(\CARRYB[28][22] ), .CI(\SUMB[28][23] ), 
        .CO(\CARRYB[29][22] ), .S(\SUMB[29][22] ) );
  FA1P S2_13_10 ( .A(n566), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), .CO(
        \CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1P S2_30_10 ( .A(n507), .B(\CARRYB[29][10] ), .CI(\SUMB[29][11] ), .CO(
        \CARRYB[30][10] ), .S(\SUMB[30][10] ) );
  FA1AP S2_32_38 ( .A(\ab[38][32] ), .B(\CARRYB[31][38] ), .CI(\SUMB[31][39] ), 
        .CO(\CARRYB[32][38] ), .S(\SUMB[32][38] ) );
  FA1P S2_33_31 ( .A(\ab[33][31] ), .B(\CARRYB[32][31] ), .CI(\SUMB[32][32] ), 
        .CO(\CARRYB[33][31] ), .S(\SUMB[33][31] ) );
  FA1P S2_42_45 ( .A(\ab[45][42] ), .B(\CARRYB[41][45] ), .CI(\SUMB[41][46] ), 
        .CO(\CARRYB[42][45] ), .S(\SUMB[42][45] ) );
  FA1AP S2_43_45 ( .A(\ab[45][43] ), .B(\CARRYB[42][45] ), .CI(\SUMB[42][46] ), 
        .CO(\CARRYB[43][45] ), .S(\SUMB[43][45] ) );
  FA1 S2_31_41 ( .A(\ab[41][31] ), .B(\CARRYB[30][41] ), .CI(\SUMB[30][42] ), 
        .CO(\CARRYB[31][41] ), .S(\SUMB[31][41] ) );
  FA1AP S2_32_41 ( .A(\ab[41][32] ), .B(\CARRYB[31][41] ), .CI(\SUMB[31][42] ), 
        .CO(\CARRYB[32][41] ), .S(\SUMB[32][41] ) );
  FA1 S2_29_39 ( .A(\ab[39][29] ), .B(\CARRYB[28][39] ), .CI(\SUMB[28][40] ), 
        .CO(\CARRYB[29][39] ), .S(\SUMB[29][39] ) );
  FA1P S2_13_12 ( .A(n604), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), .CO(
        \CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1P S2_41_44 ( .A(\ab[44][41] ), .B(\CARRYB[40][44] ), .CI(\SUMB[40][45] ), 
        .CO(\CARRYB[41][44] ), .S(\SUMB[41][44] ) );
  FA1P S2_41_45 ( .A(\ab[45][41] ), .B(\CARRYB[40][45] ), .CI(\SUMB[40][46] ), 
        .CO(\CARRYB[41][45] ), .S(\SUMB[41][45] ) );
  FA1P S2_17_22 ( .A(\ab[22][17] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA1P S2_18_22 ( .A(\ab[22][18] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA1P S2_30_36 ( .A(\ab[36][30] ), .B(\CARRYB[29][36] ), .CI(\SUMB[29][37] ), 
        .CO(\CARRYB[30][36] ), .S(\SUMB[30][36] ) );
  FA1P S2_26_37 ( .A(\ab[37][26] ), .B(\CARRYB[25][37] ), .CI(\SUMB[25][38] ), 
        .CO(\CARRYB[26][37] ), .S(\SUMB[26][37] ) );
  FA1P S2_27_37 ( .A(\ab[37][27] ), .B(\CARRYB[26][37] ), .CI(\SUMB[26][38] ), 
        .CO(\CARRYB[27][37] ), .S(\SUMB[27][37] ) );
  FA1P S2_25_38 ( .A(\ab[38][25] ), .B(\CARRYB[24][38] ), .CI(\SUMB[24][39] ), 
        .CO(\CARRYB[25][38] ), .S(\SUMB[25][38] ) );
  FA1P S2_26_38 ( .A(\ab[38][26] ), .B(\CARRYB[25][38] ), .CI(\SUMB[25][39] ), 
        .CO(\CARRYB[26][38] ), .S(\SUMB[26][38] ) );
  FA1P S3_40_46 ( .A(\ab[46][40] ), .B(\CARRYB[39][46] ), .CI(\ab[47][39] ), 
        .CO(\CARRYB[40][46] ), .S(\SUMB[40][46] ) );
  FA1P S2_12_23 ( .A(n600), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), .CO(
        \CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA1P S2_42_14 ( .A(\ab[42][14] ), .B(\CARRYB[41][14] ), .CI(\SUMB[41][15] ), 
        .CO(\CARRYB[42][14] ), .S(\SUMB[42][14] ) );
  FA1P S2_43_14 ( .A(\ab[43][14] ), .B(\CARRYB[42][14] ), .CI(\SUMB[42][15] ), 
        .CO(\CARRYB[43][14] ), .S(\SUMB[43][14] ) );
  FA1P S2_10_9 ( .A(n552), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1P S2_7_6 ( .A(n480), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1P S2_7_7 ( .A(n1453), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1AP S2_8_6 ( .A(n456), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1P S1_34_0 ( .A(n1349), .B(\CARRYB[33][0] ), .CI(\SUMB[33][1] ), .CO(
        \CARRYB[34][0] ), .S(\A1[32] ) );
  FA1P S2_14_5 ( .A(n414), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(
        \CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1P S2_15_5 ( .A(n413), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1 S2_23_23 ( .A(A[23]), .B(\CARRYB[22][23] ), .CI(\SUMB[22][24] ), .CO(
        \CARRYB[23][23] ), .S(\SUMB[23][23] ) );
  FA1P S2_27_39 ( .A(\ab[39][27] ), .B(\CARRYB[26][39] ), .CI(\SUMB[26][40] ), 
        .CO(\CARRYB[27][39] ), .S(\SUMB[27][39] ) );
  FA1P S2_28_39 ( .A(\ab[39][28] ), .B(\CARRYB[27][39] ), .CI(\SUMB[27][40] ), 
        .CO(\CARRYB[28][39] ), .S(\SUMB[28][39] ) );
  FA1P S2_25_25 ( .A(A[25]), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), .CO(
        \CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA1P S2_12_14 ( .A(n611), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), .CO(
        \CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1P S2_13_14 ( .A(n622), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), .CO(
        \CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1P S2_29_35 ( .A(\ab[35][29] ), .B(\CARRYB[28][35] ), .CI(\SUMB[28][36] ), 
        .CO(\CARRYB[29][35] ), .S(\SUMB[29][35] ) );
  FA1P S2_30_35 ( .A(\ab[35][30] ), .B(\CARRYB[29][35] ), .CI(\SUMB[29][36] ), 
        .CO(\CARRYB[30][35] ), .S(\SUMB[30][35] ) );
  FA1AP S2_9_5 ( .A(n427), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1 S2_10_4 ( .A(n378), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1AP S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), 
        .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA1 S2_44_43 ( .A(\ab[44][43] ), .B(\CARRYB[43][43] ), .CI(\SUMB[43][44] ), 
        .CO(\CARRYB[44][43] ), .S(\SUMB[44][43] ) );
  FA1P S2_20_28 ( .A(\ab[28][20] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA1P S2_21_28 ( .A(\ab[28][21] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA1P S2_5_6 ( .A(n410), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1 S2_5_7 ( .A(n426), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1AP S2_6_6 ( .A(n1449), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1P S2_25_39 ( .A(\ab[39][25] ), .B(\CARRYB[24][39] ), .CI(\SUMB[24][40] ), 
        .CO(\CARRYB[25][39] ), .S(\SUMB[25][39] ) );
  FA1A S2_25_40 ( .A(\ab[40][25] ), .B(\CARRYB[24][40] ), .CI(\SUMB[24][41] ), 
        .CO(\CARRYB[25][40] ), .S(\SUMB[25][40] ) );
  FA1P S2_26_39 ( .A(\ab[39][26] ), .B(\CARRYB[25][39] ), .CI(\SUMB[25][40] ), 
        .CO(\CARRYB[26][39] ), .S(\SUMB[26][39] ) );
  FA1P S2_32_31 ( .A(\ab[32][31] ), .B(\CARRYB[31][31] ), .CI(\SUMB[31][32] ), 
        .CO(\CARRYB[32][31] ), .S(\SUMB[32][31] ) );
  FA1P S2_3_6 ( .A(n314), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1P S2_40_32 ( .A(\ab[40][32] ), .B(\CARRYB[39][32] ), .CI(\SUMB[39][33] ), 
        .CO(\CARRYB[40][32] ), .S(\SUMB[40][32] ) );
  FA1P S2_41_32 ( .A(\ab[41][32] ), .B(\CARRYB[40][32] ), .CI(\SUMB[40][33] ), 
        .CO(\CARRYB[41][32] ), .S(\SUMB[41][32] ) );
  FA1P S2_31_40 ( .A(\ab[40][31] ), .B(\CARRYB[30][40] ), .CI(\SUMB[30][41] ), 
        .CO(\CARRYB[31][40] ), .S(\SUMB[31][40] ) );
  FA1P S2_13_8 ( .A(n487), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), .CO(
        \CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1 S2_11_11 ( .A(A[11]), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), .CO(
        \CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1 S2_11_12 ( .A(n602), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), .CO(
        \CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1AP S2_40_44 ( .A(\ab[44][40] ), .B(\CARRYB[39][44] ), .CI(\SUMB[39][45] ), 
        .CO(\CARRYB[40][44] ), .S(\SUMB[40][44] ) );
  FA1P S2_17_31 ( .A(\ab[31][17] ), .B(\CARRYB[16][31] ), .CI(\SUMB[16][32] ), 
        .CO(\CARRYB[17][31] ), .S(\SUMB[17][31] ) );
  FA1 S2_44_44 ( .A(A[44]), .B(\CARRYB[43][44] ), .CI(\SUMB[43][45] ), .CO(
        \CARRYB[44][44] ), .S(\SUMB[44][44] ) );
  FA1P S2_26_24 ( .A(\ab[26][24] ), .B(\CARRYB[25][24] ), .CI(\SUMB[25][25] ), 
        .CO(\CARRYB[26][24] ), .S(\SUMB[26][24] ) );
  FA1P S2_29_8 ( .A(\SUMB[28][9] ), .B(\CARRYB[28][8] ), .CI(n1290), .CO(
        \CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA1P S2_30_8 ( .A(n275), .B(\CARRYB[29][8] ), .CI(\SUMB[29][9] ), .CO(
        \CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA1P S2_32_5 ( .A(n390), .B(\CARRYB[31][5] ), .CI(\SUMB[31][6] ), .CO(
        \CARRYB[32][5] ), .S(\SUMB[32][5] ) );
  FA1P S2_19_27 ( .A(\ab[27][19] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA1P S2_20_27 ( .A(\ab[27][20] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA1P S2_26_41 ( .A(\ab[41][26] ), .B(\CARRYB[25][41] ), .CI(\SUMB[25][42] ), 
        .CO(\CARRYB[26][41] ), .S(\SUMB[26][41] ) );
  FA1P S3_12_46 ( .A(\ab[46][12] ), .B(\CARRYB[11][46] ), .CI(\ab[47][11] ), 
        .CO(\CARRYB[12][46] ), .S(\SUMB[12][46] ) );
  FA1AP S2_42_31 ( .A(\ab[42][31] ), .B(\CARRYB[41][31] ), .CI(\SUMB[41][32] ), 
        .CO(\CARRYB[42][31] ), .S(\SUMB[42][31] ) );
  FA1P S2_43_31 ( .A(\ab[43][31] ), .B(\CARRYB[42][31] ), .CI(\SUMB[42][32] ), 
        .CO(\CARRYB[43][31] ), .S(\SUMB[43][31] ) );
  FA1AP S2_22_38 ( .A(\ab[38][22] ), .B(\CARRYB[21][38] ), .CI(\SUMB[21][39] ), 
        .CO(\CARRYB[22][38] ), .S(\SUMB[22][38] ) );
  FA1P S2_23_38 ( .A(\ab[38][23] ), .B(\CARRYB[22][38] ), .CI(\SUMB[22][39] ), 
        .CO(\CARRYB[23][38] ), .S(\SUMB[23][38] ) );
  FA1 S3_39_46 ( .A(\ab[46][39] ), .B(\CARRYB[38][46] ), .CI(\ab[47][38] ), 
        .CO(\CARRYB[39][46] ), .S(\SUMB[39][46] ) );
  FA1A S2_11_9 ( .A(n568), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), .CO(
        \CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1AP S2_12_9 ( .A(n553), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), .CO(
        \CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1 S2_21_25 ( .A(\ab[25][21] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA1 S2_2_44 ( .A(n308), .B(\CARRYB[1][44] ), .CI(\SUMB[1][45] ), .CO(
        \CARRYB[2][44] ), .S(\SUMB[2][44] ) );
  FA1P S2_3_44 ( .A(n341), .B(\CARRYB[2][44] ), .CI(\SUMB[2][45] ), .CO(
        \CARRYB[3][44] ), .S(\SUMB[3][44] ) );
  FA1P S2_23_25 ( .A(\ab[25][23] ), .B(\CARRYB[22][25] ), .CI(\SUMB[22][26] ), 
        .CO(\CARRYB[23][25] ), .S(\SUMB[23][25] ) );
  FA1P S2_24_25 ( .A(\ab[25][24] ), .B(\CARRYB[23][25] ), .CI(\SUMB[23][26] ), 
        .CO(\CARRYB[24][25] ), .S(\SUMB[24][25] ) );
  FA1 S2_35_3 ( .A(n298), .B(\CARRYB[34][3] ), .CI(\SUMB[34][4] ), .CO(
        \CARRYB[35][3] ), .S(\SUMB[35][3] ) );
  FA1AP S3_38_46 ( .A(\ab[46][38] ), .B(\CARRYB[37][46] ), .CI(\ab[47][37] ), 
        .CO(\CARRYB[38][46] ), .S(\SUMB[38][46] ) );
  FA1P S2_21_41 ( .A(\ab[41][21] ), .B(\CARRYB[20][41] ), .CI(\SUMB[20][42] ), 
        .CO(\CARRYB[21][41] ), .S(\SUMB[21][41] ) );
  FA1AP S2_31_5 ( .A(n403), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), .CO(
        \CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FA1AP S2_34_31 ( .A(\ab[34][31] ), .B(\CARRYB[33][31] ), .CI(\SUMB[33][32] ), 
        .CO(\CARRYB[34][31] ), .S(\SUMB[34][31] ) );
  FA1P S2_27_36 ( .A(\ab[36][27] ), .B(\CARRYB[26][36] ), .CI(\SUMB[26][37] ), 
        .CO(\CARRYB[27][36] ), .S(\SUMB[27][36] ) );
  FA1P S2_28_36 ( .A(\ab[36][28] ), .B(\CARRYB[27][36] ), .CI(\SUMB[27][37] ), 
        .CO(\CARRYB[28][36] ), .S(\SUMB[28][36] ) );
  FA1AP S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA1 S2_6_28 ( .A(\CARRYB[5][28] ), .B(n396), .CI(\SUMB[5][29] ), .CO(
        \CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA1 S2_35_33 ( .A(\ab[35][33] ), .B(\CARRYB[34][33] ), .CI(\SUMB[34][34] ), 
        .CO(\CARRYB[35][33] ), .S(\SUMB[35][33] ) );
  FA1P S2_33_2 ( .A(n1306), .B(\CARRYB[32][2] ), .CI(\SUMB[32][3] ), .CO(
        \CARRYB[33][2] ), .S(\SUMB[33][2] ) );
  FA1P S2_30_34 ( .A(\ab[34][30] ), .B(\CARRYB[29][34] ), .CI(\SUMB[29][35] ), 
        .CO(\CARRYB[30][34] ), .S(\SUMB[30][34] ) );
  FA1P S2_31_34 ( .A(\ab[34][31] ), .B(\CARRYB[30][34] ), .CI(\SUMB[30][35] ), 
        .CO(\CARRYB[31][34] ), .S(\SUMB[31][34] ) );
  FA1P S2_8_10 ( .A(n508), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), .CO(
        \CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1P S1_32_0 ( .A(n871), .B(\CARRYB[31][0] ), .CI(\SUMB[31][1] ), .CO(
        \CARRYB[32][0] ), .S(\A1[30] ) );
  FA1P S1_33_0 ( .A(n1326), .B(\CARRYB[32][0] ), .CI(\SUMB[32][1] ), .CO(
        \CARRYB[33][0] ), .S(\A1[31] ) );
  FA1P S2_19_28 ( .A(\ab[28][19] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA1P S2_15_24 ( .A(\ab[24][15] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA1P S2_16_24 ( .A(\ab[24][16] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA1 S2_32_4 ( .A(n376), .B(\CARRYB[31][4] ), .CI(\SUMB[31][5] ), .CO(
        \CARRYB[32][4] ), .S(\SUMB[32][4] ) );
  FA1P S2_32_30 ( .A(\ab[32][30] ), .B(\CARRYB[31][30] ), .CI(\SUMB[31][31] ), 
        .CO(\CARRYB[32][30] ), .S(\SUMB[32][30] ) );
  FA1P S2_33_30 ( .A(\ab[33][30] ), .B(\CARRYB[32][30] ), .CI(\SUMB[32][31] ), 
        .CO(\CARRYB[33][30] ), .S(\SUMB[33][30] ) );
  FA1P S2_24_43 ( .A(\ab[43][24] ), .B(\CARRYB[23][43] ), .CI(\SUMB[23][44] ), 
        .CO(\CARRYB[24][43] ), .S(\SUMB[24][43] ) );
  FA1AP S2_35_14 ( .A(\ab[35][14] ), .B(\CARRYB[34][14] ), .CI(\SUMB[34][15] ), 
        .CO(\CARRYB[35][14] ), .S(\SUMB[35][14] ) );
  FA1P S2_30_31 ( .A(\ab[31][30] ), .B(\CARRYB[29][31] ), .CI(\SUMB[29][32] ), 
        .CO(\CARRYB[30][31] ), .S(\SUMB[30][31] ) );
  FA1P S2_31_31 ( .A(n1493), .B(\CARRYB[30][31] ), .CI(\SUMB[30][32] ), .CO(
        \CARRYB[31][31] ), .S(\SUMB[31][31] ) );
  FA1 S2_32_14 ( .A(\ab[32][14] ), .B(\CARRYB[31][14] ), .CI(\SUMB[31][15] ), 
        .CO(\CARRYB[32][14] ), .S(\SUMB[32][14] ) );
  FA1AP S2_33_14 ( .A(\ab[33][14] ), .B(\CARRYB[32][14] ), .CI(\SUMB[32][15] ), 
        .CO(\CARRYB[33][14] ), .S(\SUMB[33][14] ) );
  FA1 S2_16_8 ( .A(n518), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), .CO(
        \CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1P S2_32_1 ( .A(n1323), .B(\CARRYB[31][1] ), .CI(\SUMB[31][2] ), .CO(
        \CARRYB[32][1] ), .S(\SUMB[32][1] ) );
  FA1P S2_16_23 ( .A(\ab[23][16] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA1P S2_17_23 ( .A(\ab[23][17] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA1AP S2_26_14 ( .A(n645), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), .CO(
        \CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA1A S2_41_42 ( .A(\ab[42][41] ), .B(\CARRYB[40][42] ), .CI(\SUMB[40][43] ), 
        .CO(\CARRYB[41][42] ), .S(\SUMB[41][42] ) );
  FA1P S2_39_42 ( .A(\ab[42][39] ), .B(\CARRYB[38][42] ), .CI(\SUMB[38][43] ), 
        .CO(\CARRYB[39][42] ), .S(\SUMB[39][42] ) );
  FA1P S4_7 ( .A(\ab[7][47] ), .B(\CARRYB[46][7] ), .CI(\SUMB[46][8] ), .CO(
        \CARRYB[47][7] ), .S(\SUMB[47][7] ) );
  FA1AP S2_20_44 ( .A(\ab[44][20] ), .B(\CARRYB[19][44] ), .CI(\SUMB[19][45] ), 
        .CO(\CARRYB[20][44] ), .S(\SUMB[20][44] ) );
  FA1P S2_29_32 ( .A(\ab[32][29] ), .B(\CARRYB[28][32] ), .CI(\SUMB[28][33] ), 
        .CO(\CARRYB[29][32] ), .S(\SUMB[29][32] ) );
  FA1P S2_9_9 ( .A(A[9]), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1AP S2_9_8 ( .A(n526), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1P S2_12_40 ( .A(\ab[40][12] ), .B(\CARRYB[11][40] ), .CI(\SUMB[11][41] ), 
        .CO(\CARRYB[12][40] ), .S(\SUMB[12][40] ) );
  FA1AP S2_6_42 ( .A(n455), .B(\CARRYB[5][42] ), .CI(\SUMB[5][43] ), .CO(
        \CARRYB[6][42] ), .S(\SUMB[6][42] ) );
  FA1P S2_29_42 ( .A(\ab[42][29] ), .B(\CARRYB[28][42] ), .CI(\SUMB[28][43] ), 
        .CO(\CARRYB[29][42] ), .S(\SUMB[29][42] ) );
  FA1A S2_20_45 ( .A(\ab[45][20] ), .B(\CARRYB[19][45] ), .CI(\SUMB[19][46] ), 
        .CO(\CARRYB[20][45] ), .S(\SUMB[20][45] ) );
  FA1P S3_18_46 ( .A(\ab[46][18] ), .B(\CARRYB[17][46] ), .CI(\ab[47][17] ), 
        .CO(\CARRYB[18][46] ), .S(\SUMB[18][46] ) );
  FA1P S2_7_10 ( .A(n503), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), .CO(
        \CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1 S2_7_9 ( .A(n514), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1P S2_19_41 ( .A(\ab[41][19] ), .B(\CARRYB[18][41] ), .CI(\SUMB[18][42] ), 
        .CO(\CARRYB[19][41] ), .S(\SUMB[19][41] ) );
  FA1P S2_38_22 ( .A(\ab[38][22] ), .B(\CARRYB[37][22] ), .CI(\SUMB[37][23] ), 
        .CO(\CARRYB[38][22] ), .S(\SUMB[38][22] ) );
  FA1P S2_38_21 ( .A(\ab[38][21] ), .B(\CARRYB[37][21] ), .CI(\SUMB[37][22] ), 
        .CO(\CARRYB[38][21] ), .S(\SUMB[38][21] ) );
  FA1AP S2_7_41 ( .A(n463), .B(\CARRYB[6][41] ), .CI(\SUMB[6][42] ), .CO(
        \CARRYB[7][41] ), .S(\SUMB[7][41] ) );
  FA1AP S2_5_42 ( .A(n402), .B(\CARRYB[4][42] ), .CI(\SUMB[4][43] ), .CO(
        \CARRYB[5][42] ), .S(\SUMB[5][42] ) );
  FA1P S2_5_41 ( .A(n385), .B(\CARRYB[4][41] ), .CI(\SUMB[4][42] ), .CO(
        \CARRYB[5][41] ), .S(\SUMB[5][41] ) );
  FA1AP S2_15_23 ( .A(\ab[23][15] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA1P S2_14_15 ( .A(n641), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), .CO(
        \CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1P S2_24_10 ( .A(n554), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), .CO(
        \CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA1P S3_16_46 ( .A(\ab[46][16] ), .B(\CARRYB[15][46] ), .CI(\ab[47][15] ), 
        .CO(\CARRYB[16][46] ), .S(\SUMB[16][46] ) );
  FA1AP S2_6_21 ( .A(n439), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), .CO(
        \CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA1P S2_4_21 ( .A(n363), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), .CO(
        \CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA1AP S2_14_10 ( .A(n569), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), .CO(
        \CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1P S2_12_12 ( .A(A[12]), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), .CO(
        \CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1 S2_5_43 ( .A(n399), .B(\CARRYB[4][43] ), .CI(\SUMB[4][44] ), .CO(
        \CARRYB[5][43] ), .S(\SUMB[5][43] ) );
  FA1 S2_3_43 ( .A(\CARRYB[2][43] ), .B(n1320), .CI(\SUMB[2][44] ), .CO(
        \CARRYB[3][43] ), .S(\SUMB[3][43] ) );
  FA1A S2_29_6 ( .A(n1279), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), .CO(
        \CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA1P S2_26_6 ( .A(n433), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), .CO(
        \CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA1P S2_30_5 ( .A(n319), .B(\CARRYB[29][5] ), .CI(\SUMB[29][6] ), .CO(
        \CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA1P S2_30_4 ( .A(n339), .B(\CARRYB[29][4] ), .CI(\SUMB[29][5] ), .CO(
        \CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA1AP S2_15_31 ( .A(\ab[31][15] ), .B(\CARRYB[14][31] ), .CI(\SUMB[14][32] ), 
        .CO(\CARRYB[15][31] ), .S(\SUMB[15][31] ) );
  FA1AP S2_7_11 ( .A(n494), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), .CO(
        \CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1P S2_19_35 ( .A(\ab[35][19] ), .B(\CARRYB[18][35] ), .CI(\SUMB[18][36] ), 
        .CO(\CARRYB[19][35] ), .S(\SUMB[19][35] ) );
  FA1P S2_4_11 ( .A(n381), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), .CO(
        \CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1P S2_2_11 ( .A(n312), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), .CO(
        \CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1P S2_45_30 ( .A(\ab[45][30] ), .B(\CARRYB[44][30] ), .CI(\SUMB[44][31] ), 
        .CO(\CARRYB[45][30] ), .S(\SUMB[45][30] ) );
  FA1AP S2_45_29 ( .A(\ab[45][29] ), .B(\CARRYB[44][29] ), .CI(\SUMB[44][30] ), 
        .CO(\CARRYB[45][29] ), .S(\SUMB[45][29] ) );
  FA1AP S2_12_17 ( .A(n608), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), .CO(
        \CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA1P S2_10_17 ( .A(n556), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), .CO(
        \CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1AP S2_19_44 ( .A(\ab[44][19] ), .B(\CARRYB[18][44] ), .CI(\SUMB[18][45] ), 
        .CO(\CARRYB[19][44] ), .S(\SUMB[19][44] ) );
  FA1 S2_17_44 ( .A(\ab[44][17] ), .B(\CARRYB[16][44] ), .CI(\SUMB[16][45] ), 
        .CO(\CARRYB[17][44] ), .S(\SUMB[17][44] ) );
  FA1P S2_14_6 ( .A(n438), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), .CO(
        \CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1P S1_31_0 ( .A(n1342), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), .CO(
        \CARRYB[31][0] ), .S(\A1[29] ) );
  FA1P S1_26_0 ( .A(n1337), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), .CO(
        \CARRYB[26][0] ), .S(\A1[24] ) );
  FA1 S1_39_0 ( .A(n1365), .B(\CARRYB[38][0] ), .CI(\SUMB[38][1] ), .CO(
        \CARRYB[39][0] ), .S(\A1[37] ) );
  FA1 S4_0 ( .A(n1327), .B(\CARRYB[46][0] ), .CI(\SUMB[46][1] ), .CO(
        \CARRYB[47][0] ), .S(\SUMB[47][0] ) );
  FA1A S4_1 ( .A(n1343), .B(\CARRYB[46][1] ), .CI(\SUMB[46][2] ), .CO(
        \CARRYB[47][1] ), .S(\SUMB[47][1] ) );
  FA1 S1_13_0 ( .A(n1358), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), .CO(
        \CARRYB[13][0] ), .S(\A1[11] ) );
  FA1 S2_11_1 ( .A(n1382), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(
        \CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1P S2_40_1 ( .A(n1348), .B(\CARRYB[39][1] ), .CI(\SUMB[39][2] ), .CO(
        \CARRYB[40][1] ), .S(\SUMB[40][1] ) );
  FA1P S2_9_32 ( .A(n501), .B(\CARRYB[8][32] ), .CI(\SUMB[8][33] ), .CO(
        \CARRYB[9][32] ), .S(\SUMB[9][32] ) );
  FA1 S2_10_32 ( .A(n551), .B(\CARRYB[9][32] ), .CI(\SUMB[9][33] ), .CO(
        \CARRYB[10][32] ), .S(\SUMB[10][32] ) );
  FA1P S2_46_23 ( .A(\ab[46][23] ), .B(\CARRYB[45][23] ), .CI(\SUMB[45][24] ), 
        .CO(\CARRYB[46][23] ), .S(\SUMB[46][23] ) );
  FA1 S2_27_29 ( .A(\ab[29][27] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA1P S2_37_26 ( .A(\ab[37][26] ), .B(\CARRYB[36][26] ), .CI(\SUMB[36][27] ), 
        .CO(\CARRYB[37][26] ), .S(\SUMB[37][26] ) );
  FA1P S2_5_10 ( .A(n437), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), .CO(
        \CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1 S2_11_10 ( .A(n575), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), .CO(
        \CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1AP S2_12_10 ( .A(n576), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), .CO(
        \CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1P S2_6_10 ( .A(n464), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), .CO(
        \CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1P S2_42_3 ( .A(n1380), .B(\CARRYB[41][3] ), .CI(\SUMB[41][4] ), .CO(
        \CARRYB[42][3] ), .S(\SUMB[42][3] ) );
  FA1P S2_43_3 ( .A(n1320), .B(\CARRYB[42][3] ), .CI(\SUMB[42][4] ), .CO(
        \CARRYB[43][3] ), .S(\SUMB[43][3] ) );
  FA1AP S2_2_43 ( .A(n1302), .B(\CARRYB[1][43] ), .CI(\SUMB[1][44] ), .CO(
        \CARRYB[2][43] ), .S(\SUMB[2][43] ) );
  FA1AP S2_10_39 ( .A(\CARRYB[9][39] ), .B(\ab[39][10] ), .CI(\SUMB[9][40] ), 
        .CO(\CARRYB[10][39] ), .S(\SUMB[10][39] ) );
  FA1P S2_23_34 ( .A(\ab[34][23] ), .B(\CARRYB[22][34] ), .CI(\SUMB[22][35] ), 
        .CO(\CARRYB[23][34] ), .S(\SUMB[23][34] ) );
  FA1AP S2_27_34 ( .A(\ab[34][27] ), .B(\CARRYB[26][34] ), .CI(\SUMB[26][35] ), 
        .CO(\CARRYB[27][34] ), .S(\SUMB[27][34] ) );
  FA1P S2_38_32 ( .A(\ab[38][32] ), .B(\CARRYB[37][32] ), .CI(\SUMB[37][33] ), 
        .CO(\CARRYB[38][32] ), .S(\SUMB[38][32] ) );
  FA1P S2_39_32 ( .A(\ab[39][32] ), .B(\CARRYB[38][32] ), .CI(\SUMB[38][33] ), 
        .CO(\CARRYB[39][32] ), .S(\SUMB[39][32] ) );
  FA1 S2_33_32 ( .A(\ab[33][32] ), .B(\CARRYB[32][32] ), .CI(\SUMB[32][33] ), 
        .CO(\CARRYB[33][32] ), .S(\SUMB[33][32] ) );
  FA1AP S2_34_32 ( .A(\ab[34][32] ), .B(\CARRYB[33][32] ), .CI(\SUMB[33][33] ), 
        .CO(\CARRYB[34][32] ), .S(\SUMB[34][32] ) );
  FA1P S2_13_22 ( .A(n620), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), .CO(
        \CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA1P S2_14_22 ( .A(n646), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), .CO(
        \CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA1P S2_45_19 ( .A(\ab[45][19] ), .B(\CARRYB[44][19] ), .CI(\SUMB[44][20] ), 
        .CO(\CARRYB[45][19] ), .S(\SUMB[45][19] ) );
  FA1 S2_7_23 ( .A(n466), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), .CO(
        \CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA1P S2_16_21 ( .A(\ab[21][16] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA1P S2_34_21 ( .A(\ab[34][21] ), .B(\CARRYB[33][21] ), .CI(\SUMB[33][22] ), 
        .CO(\CARRYB[34][21] ), .S(\SUMB[34][21] ) );
  FA1P S2_35_21 ( .A(\ab[35][21] ), .B(\CARRYB[34][21] ), .CI(\SUMB[34][22] ), 
        .CO(\CARRYB[35][21] ), .S(\SUMB[35][21] ) );
  FA1P S2_14_40 ( .A(\ab[40][14] ), .B(\CARRYB[13][40] ), .CI(\SUMB[13][41] ), 
        .CO(\CARRYB[14][40] ), .S(\SUMB[14][40] ) );
  FA1P S2_9_41 ( .A(\CARRYB[8][41] ), .B(\ab[9][41] ), .CI(\SUMB[8][42] ), 
        .CO(\CARRYB[9][41] ), .S(\SUMB[9][41] ) );
  FA1P S2_36_36 ( .A(\ab[36][36] ), .B(\CARRYB[35][36] ), .CI(\SUMB[35][37] ), 
        .CO(\CARRYB[36][36] ), .S(\SUMB[36][36] ) );
  FA1P S2_46_35 ( .A(\ab[46][35] ), .B(\CARRYB[45][35] ), .CI(\SUMB[45][36] ), 
        .CO(\CARRYB[46][35] ), .S(\SUMB[46][35] ) );
  FA1P S4_35 ( .A(\ab[47][35] ), .B(\CARRYB[46][35] ), .CI(\SUMB[46][36] ), 
        .CO(\CARRYB[47][35] ), .S(\SUMB[47][35] ) );
  FA1P S4_34 ( .A(\ab[47][34] ), .B(\CARRYB[46][34] ), .CI(\SUMB[46][35] ), 
        .CO(\CARRYB[47][34] ), .S(\SUMB[47][34] ) );
  FA1P S2_18_39 ( .A(\ab[39][18] ), .B(\CARRYB[17][39] ), .CI(\SUMB[17][40] ), 
        .CO(\CARRYB[18][39] ), .S(\SUMB[18][39] ) );
  FA1 S2_10_26 ( .A(\SUMB[9][27] ), .B(\CARRYB[9][26] ), .CI(n544), .CO(
        \CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA1P S2_24_24 ( .A(n1479), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), .CO(
        \CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA1P S2_25_24 ( .A(\ab[25][24] ), .B(\CARRYB[24][24] ), .CI(\SUMB[24][25] ), 
        .CO(\CARRYB[25][24] ), .S(\SUMB[25][24] ) );
  FA1P S2_33_22 ( .A(\ab[33][22] ), .B(\CARRYB[32][22] ), .CI(\SUMB[32][23] ), 
        .CO(\CARRYB[33][22] ), .S(\SUMB[33][22] ) );
  FA1P S2_34_22 ( .A(\ab[34][22] ), .B(\CARRYB[33][22] ), .CI(\SUMB[33][23] ), 
        .CO(\CARRYB[34][22] ), .S(\SUMB[34][22] ) );
  FA1AP S2_5_29 ( .A(n1276), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), .CO(
        \CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA1P S2_43_21 ( .A(\ab[43][21] ), .B(\CARRYB[42][21] ), .CI(\SUMB[42][22] ), 
        .CO(\CARRYB[43][21] ), .S(\SUMB[43][21] ) );
  FA1P S2_44_21 ( .A(\ab[44][21] ), .B(\CARRYB[43][21] ), .CI(\SUMB[43][22] ), 
        .CO(\CARRYB[44][21] ), .S(\SUMB[44][21] ) );
  FA1P S2_26_2 ( .A(n299), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), .CO(
        \CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA1P S2_27_2 ( .A(n1310), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), .CO(
        \CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA1AP S2_38_2 ( .A(n1312), .B(\CARRYB[37][2] ), .CI(\SUMB[37][3] ), .CO(
        \CARRYB[38][2] ), .S(\SUMB[38][2] ) );
  FA1P S2_39_2 ( .A(n1313), .B(\CARRYB[38][2] ), .CI(\SUMB[38][3] ), .CO(
        \CARRYB[39][2] ), .S(\SUMB[39][2] ) );
  FA1 S2_2_2 ( .A(A[2]), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1 S2_16_2 ( .A(n1299), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), .CO(
        \CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1 S2_12_2 ( .A(n332), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), .CO(
        \CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1 S2_21_2 ( .A(n1305), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), .CO(
        \CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1 S2_37_45 ( .A(\ab[45][37] ), .B(\CARRYB[36][45] ), .CI(\SUMB[36][46] ), 
        .CO(\CARRYB[37][45] ), .S(\SUMB[37][45] ) );
  FA1P S3_37_46 ( .A(\ab[46][37] ), .B(\CARRYB[36][46] ), .CI(\ab[47][36] ), 
        .CO(\CARRYB[37][46] ), .S(\SUMB[37][46] ) );
  FA1 S2_38_45 ( .A(\ab[45][38] ), .B(\CARRYB[37][45] ), .CI(\SUMB[37][46] ), 
        .CO(\CARRYB[38][45] ), .S(\SUMB[38][45] ) );
  FA1 S2_42_44 ( .A(\ab[44][42] ), .B(\CARRYB[41][44] ), .CI(\SUMB[41][45] ), 
        .CO(\CARRYB[42][44] ), .S(\SUMB[42][44] ) );
  FA1P S2_43_44 ( .A(\ab[44][43] ), .B(\CARRYB[42][44] ), .CI(\SUMB[42][45] ), 
        .CO(\CARRYB[43][44] ), .S(\SUMB[43][44] ) );
  FA1 S2_18_45 ( .A(\ab[45][18] ), .B(\CARRYB[17][45] ), .CI(\SUMB[17][46] ), 
        .CO(\CARRYB[18][45] ), .S(\SUMB[18][45] ) );
  FA1P S2_29_45 ( .A(\ab[45][29] ), .B(\CARRYB[28][45] ), .CI(\SUMB[28][46] ), 
        .CO(\CARRYB[29][45] ), .S(\SUMB[29][45] ) );
  FA1 S2_30_45 ( .A(\ab[45][30] ), .B(\CARRYB[29][45] ), .CI(\SUMB[29][46] ), 
        .CO(\CARRYB[30][45] ), .S(\SUMB[30][45] ) );
  FA1 S2_39_45 ( .A(\ab[45][39] ), .B(\CARRYB[38][45] ), .CI(\SUMB[38][46] ), 
        .CO(\CARRYB[39][45] ), .S(\SUMB[39][45] ) );
  FA1A S2_40_45 ( .A(\ab[45][40] ), .B(\CARRYB[39][45] ), .CI(\SUMB[39][46] ), 
        .CO(\CARRYB[40][45] ), .S(\SUMB[40][45] ) );
  FA1P S2_23_44 ( .A(\ab[44][23] ), .B(\CARRYB[22][44] ), .CI(\SUMB[22][45] ), 
        .CO(\CARRYB[23][44] ), .S(\SUMB[23][44] ) );
  FA1A S2_42_42 ( .A(n1515), .B(\CARRYB[41][42] ), .CI(\SUMB[41][43] ), .CO(
        \CARRYB[42][42] ), .S(\SUMB[42][42] ) );
  FA1P S2_6_16 ( .A(n431), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), .CO(
        \CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1P S2_12_15 ( .A(n617), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), .CO(
        \CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1P S2_13_15 ( .A(n628), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), .CO(
        \CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1P S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA1P S2_19_15 ( .A(\CARRYB[18][15] ), .B(\ab[19][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA1P S2_45_8 ( .A(\ab[8][45] ), .B(\CARRYB[44][8] ), .CI(\SUMB[44][9] ), 
        .CO(\CARRYB[45][8] ), .S(\SUMB[45][8] ) );
  FA1P S2_41_25 ( .A(\ab[41][25] ), .B(\CARRYB[40][25] ), .CI(\SUMB[40][26] ), 
        .CO(\CARRYB[41][25] ), .S(\SUMB[41][25] ) );
  FA1P S2_43_25 ( .A(\ab[43][25] ), .B(\CARRYB[42][25] ), .CI(\SUMB[42][26] ), 
        .CO(\CARRYB[43][25] ), .S(\SUMB[43][25] ) );
  FA1 S2_28_7 ( .A(n424), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), .CO(
        \CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA1P S2_2_14 ( .A(n342), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1P S2_18_13 ( .A(n623), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), .CO(
        \CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA1P S2_29_12 ( .A(n609), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), .CO(
        \CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA1A S2_27_12 ( .A(n603), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), .CO(
        \CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA1P S2_39_10 ( .A(\ab[39][10] ), .B(\CARRYB[38][10] ), .CI(\SUMB[38][11] ), 
        .CO(\CARRYB[39][10] ), .S(\SUMB[39][10] ) );
  FA1P S2_40_10 ( .A(\ab[40][10] ), .B(\CARRYB[39][10] ), .CI(\SUMB[39][11] ), 
        .CO(\CARRYB[40][10] ), .S(\SUMB[40][10] ) );
  FA1P S2_33_11 ( .A(n573), .B(\CARRYB[32][11] ), .CI(\SUMB[32][12] ), .CO(
        \CARRYB[33][11] ), .S(\SUMB[33][11] ) );
  FA1P S2_46_9 ( .A(\ab[9][46] ), .B(\CARRYB[45][9] ), .CI(\SUMB[45][10] ), 
        .CO(\CARRYB[46][9] ), .S(\SUMB[46][9] ) );
  FA1P S4_9 ( .A(\ab[9][47] ), .B(\CARRYB[46][9] ), .CI(\SUMB[46][10] ), .CO(
        \CARRYB[47][9] ), .S(\SUMB[47][9] ) );
  FA1 S2_25_36 ( .A(\ab[36][25] ), .B(\CARRYB[24][36] ), .CI(\SUMB[24][37] ), 
        .CO(\CARRYB[25][36] ), .S(\SUMB[25][36] ) );
  FA1AP S2_26_36 ( .A(\ab[36][26] ), .B(\CARRYB[25][36] ), .CI(\SUMB[25][37] ), 
        .CO(\CARRYB[26][36] ), .S(\SUMB[26][36] ) );
  FA1P S2_45_34 ( .A(\ab[45][34] ), .B(\CARRYB[44][34] ), .CI(\SUMB[44][35] ), 
        .CO(\CARRYB[45][34] ), .S(\SUMB[45][34] ) );
  FA1P S2_45_35 ( .A(\ab[45][35] ), .B(\CARRYB[44][35] ), .CI(\SUMB[44][36] ), 
        .CO(\CARRYB[45][35] ), .S(\SUMB[45][35] ) );
  FA1AP S2_46_34 ( .A(\ab[46][34] ), .B(\CARRYB[45][34] ), .CI(\SUMB[45][35] ), 
        .CO(\CARRYB[46][34] ), .S(\SUMB[46][34] ) );
  FA1P S2_41_34 ( .A(\ab[41][34] ), .B(\CARRYB[40][34] ), .CI(\SUMB[40][35] ), 
        .CO(\CARRYB[41][34] ), .S(\SUMB[41][34] ) );
  FA1AP S2_18_34 ( .A(\ab[34][18] ), .B(\CARRYB[17][34] ), .CI(\SUMB[17][35] ), 
        .CO(\CARRYB[18][34] ), .S(\SUMB[18][34] ) );
  FA1 S2_32_28 ( .A(\CARRYB[31][28] ), .B(\ab[32][28] ), .CI(\SUMB[31][29] ), 
        .CO(\CARRYB[32][28] ), .S(\SUMB[32][28] ) );
  FA1AP S2_33_28 ( .A(\ab[33][28] ), .B(\CARRYB[32][28] ), .CI(\SUMB[32][29] ), 
        .CO(\CARRYB[33][28] ), .S(\SUMB[33][28] ) );
  FA1AP S2_2_41 ( .A(n1311), .B(\CARRYB[1][41] ), .CI(\SUMB[1][42] ), .CO(
        \CARRYB[2][41] ), .S(\SUMB[2][41] ) );
  FA1 S2_14_36 ( .A(\ab[36][14] ), .B(\CARRYB[13][36] ), .CI(\SUMB[13][37] ), 
        .CO(\CARRYB[14][36] ), .S(\SUMB[14][36] ) );
  FA1P S2_19_32 ( .A(\CARRYB[18][32] ), .B(\ab[32][19] ), .CI(\SUMB[18][33] ), 
        .CO(\CARRYB[19][32] ), .S(\SUMB[19][32] ) );
  FA1AP S2_20_32 ( .A(\ab[32][20] ), .B(\CARRYB[19][32] ), .CI(\SUMB[19][33] ), 
        .CO(\CARRYB[20][32] ), .S(\SUMB[20][32] ) );
  FA1P S2_37_28 ( .A(\ab[37][28] ), .B(\CARRYB[36][28] ), .CI(\SUMB[36][29] ), 
        .CO(\CARRYB[37][28] ), .S(\SUMB[37][28] ) );
  FA1P S2_38_28 ( .A(\ab[38][28] ), .B(\CARRYB[37][28] ), .CI(\SUMB[37][29] ), 
        .CO(\CARRYB[38][28] ), .S(\SUMB[38][28] ) );
  FA1P S2_46_28 ( .A(\ab[46][28] ), .B(\CARRYB[45][28] ), .CI(\SUMB[45][29] ), 
        .CO(\CARRYB[46][28] ), .S(\SUMB[46][28] ) );
  FA1AP S4_28 ( .A(\ab[47][28] ), .B(\CARRYB[46][28] ), .CI(\SUMB[46][29] ), 
        .CO(\CARRYB[47][28] ), .S(\SUMB[47][28] ) );
  FA1P S2_21_36 ( .A(\SUMB[20][37] ), .B(\CARRYB[20][36] ), .CI(\ab[36][21] ), 
        .CO(\CARRYB[21][36] ), .S(\SUMB[21][36] ) );
  FA1P S2_42_33 ( .A(\ab[42][33] ), .B(\CARRYB[41][33] ), .CI(\SUMB[41][34] ), 
        .CO(\CARRYB[42][33] ), .S(\SUMB[42][33] ) );
  FA1P S2_43_33 ( .A(\ab[43][33] ), .B(\CARRYB[42][33] ), .CI(\SUMB[42][34] ), 
        .CO(\CARRYB[43][33] ), .S(\SUMB[43][33] ) );
  FA1A S2_22_42 ( .A(\ab[42][22] ), .B(\CARRYB[21][42] ), .CI(\SUMB[21][43] ), 
        .CO(\CARRYB[22][42] ), .S(\SUMB[22][42] ) );
  FA1 S2_14_38 ( .A(\ab[38][14] ), .B(\CARRYB[13][38] ), .CI(\SUMB[13][39] ), 
        .CO(\CARRYB[14][38] ), .S(\SUMB[14][38] ) );
  FA1P S2_37_32 ( .A(\ab[37][32] ), .B(\CARRYB[36][32] ), .CI(\SUMB[36][33] ), 
        .CO(\CARRYB[37][32] ), .S(\SUMB[37][32] ) );
  FA1AP S2_15_38 ( .A(\ab[38][15] ), .B(\CARRYB[14][38] ), .CI(\SUMB[14][39] ), 
        .CO(\CARRYB[15][38] ), .S(\SUMB[15][38] ) );
  FA1P S2_35_32 ( .A(\ab[35][32] ), .B(\CARRYB[34][32] ), .CI(\SUMB[34][33] ), 
        .CO(\CARRYB[35][32] ), .S(\SUMB[35][32] ) );
  FA1 S2_5_12 ( .A(n441), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), .CO(
        \CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1P S2_6_12 ( .A(n476), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), .CO(
        \CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_16_9 ( .A(n535), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), .CO(
        \CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1P S2_14_9 ( .A(n536), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), .CO(
        \CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1P S2_44_7 ( .A(n467), .B(\CARRYB[43][7] ), .CI(\SUMB[43][8] ), .CO(
        \CARRYB[44][7] ), .S(\SUMB[44][7] ) );
  FA1P S2_45_7 ( .A(n473), .B(\CARRYB[44][7] ), .CI(\SUMB[44][8] ), .CO(
        \CARRYB[45][7] ), .S(\SUMB[45][7] ) );
  FA1P S2_28_9 ( .A(n502), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), .CO(
        \CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA1 S2_42_7 ( .A(n498), .B(\CARRYB[41][7] ), .CI(\SUMB[41][8] ), .CO(
        \CARRYB[42][7] ), .S(\SUMB[42][7] ) );
  FA1 S2_17_4 ( .A(n1278), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), .CO(
        \CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1 S2_25_4 ( .A(n357), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), .CO(
        \CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA1P S2_33_3 ( .A(n318), .B(\CARRYB[32][3] ), .CI(\SUMB[32][4] ), .CO(
        \CARRYB[33][3] ), .S(\SUMB[33][3] ) );
  FA1P S2_3_30 ( .A(n300), .B(\CARRYB[2][30] ), .CI(\SUMB[2][31] ), .CO(
        \CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA1P S2_4_30 ( .A(n339), .B(\CARRYB[3][30] ), .CI(\SUMB[3][31] ), .CO(
        \CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA1P S2_5_30 ( .A(n319), .B(\CARRYB[4][30] ), .CI(\SUMB[4][31] ), .CO(
        \CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA1AP S2_22_24 ( .A(\ab[24][22] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA1P S2_19_29 ( .A(\ab[29][19] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA1 S2_34_27 ( .A(\ab[34][27] ), .B(\CARRYB[33][27] ), .CI(\SUMB[33][28] ), 
        .CO(\CARRYB[34][27] ), .S(\SUMB[34][27] ) );
  FA1AP S2_35_27 ( .A(\ab[35][27] ), .B(\CARRYB[34][27] ), .CI(\SUMB[34][28] ), 
        .CO(\CARRYB[35][27] ), .S(\SUMB[35][27] ) );
  FA1P S2_45_24 ( .A(\ab[45][24] ), .B(\CARRYB[44][24] ), .CI(\SUMB[44][25] ), 
        .CO(\CARRYB[45][24] ), .S(\SUMB[45][24] ) );
  FA1 S2_21_45 ( .A(\ab[45][21] ), .B(\CARRYB[20][45] ), .CI(\SUMB[20][46] ), 
        .CO(\CARRYB[21][45] ), .S(\SUMB[21][45] ) );
  FA1 S2_22_45 ( .A(\ab[45][22] ), .B(\CARRYB[21][45] ), .CI(\SUMB[21][46] ), 
        .CO(\CARRYB[22][45] ), .S(\SUMB[22][45] ) );
  FA1AP S2_38_44 ( .A(\ab[44][38] ), .B(\CARRYB[37][44] ), .CI(\SUMB[37][45] ), 
        .CO(\CARRYB[38][44] ), .S(\SUMB[38][44] ) );
  FA1P S2_41_43 ( .A(\ab[43][41] ), .B(\CARRYB[40][43] ), .CI(\SUMB[40][44] ), 
        .CO(\CARRYB[41][43] ), .S(\SUMB[41][43] ) );
  FA1P S2_17_37 ( .A(\ab[37][17] ), .B(\CARRYB[16][37] ), .CI(\SUMB[16][38] ), 
        .CO(\CARRYB[17][37] ), .S(\SUMB[17][37] ) );
  FA1P S3_35_46 ( .A(\ab[46][35] ), .B(\CARRYB[34][46] ), .CI(\ab[47][34] ), 
        .CO(\CARRYB[35][46] ), .S(\SUMB[35][46] ) );
  FA1P S3_36_46 ( .A(\ab[46][36] ), .B(\CARRYB[35][46] ), .CI(\ab[47][35] ), 
        .CO(\CARRYB[36][46] ), .S(\SUMB[36][46] ) );
  FA1 S2_46_42 ( .A(\ab[46][42] ), .B(\CARRYB[45][42] ), .CI(\SUMB[45][43] ), 
        .CO(\CARRYB[46][42] ), .S(\SUMB[46][42] ) );
  FA1AP S2_42_43 ( .A(\ab[43][42] ), .B(\CARRYB[41][43] ), .CI(\SUMB[41][44] ), 
        .CO(\CARRYB[42][43] ), .S(\SUMB[42][43] ) );
  FA1 S2_43_43 ( .A(n1520), .B(\CARRYB[42][43] ), .CI(\SUMB[42][44] ), .CO(
        \CARRYB[43][43] ), .S(\SUMB[43][43] ) );
  FA1AP S4_42 ( .A(\ab[47][42] ), .B(\CARRYB[46][42] ), .CI(\SUMB[46][43] ), 
        .CO(\CARRYB[47][42] ), .S(\SUMB[47][42] ) );
  FA1P S3_15_46 ( .A(\ab[46][15] ), .B(\CARRYB[14][46] ), .CI(\ab[47][14] ), 
        .CO(\CARRYB[15][46] ), .S(\SUMB[15][46] ) );
  FA1P S3_20_46 ( .A(\ab[46][20] ), .B(\CARRYB[19][46] ), .CI(\ab[47][19] ), 
        .CO(\CARRYB[20][46] ), .S(\SUMB[20][46] ) );
  FA1P S3_19_46 ( .A(\ab[46][19] ), .B(\CARRYB[18][46] ), .CI(\ab[47][18] ), 
        .CO(\CARRYB[19][46] ), .S(\SUMB[19][46] ) );
  FA1AP S2_4_22 ( .A(n313), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), .CO(
        \CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA1AP S2_31_16 ( .A(\ab[31][16] ), .B(\CARRYB[30][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FA1AP S2_16_37 ( .A(\ab[37][16] ), .B(\CARRYB[15][37] ), .CI(\SUMB[15][38] ), 
        .CO(\CARRYB[16][37] ), .S(\SUMB[16][37] ) );
  FA1AP S2_25_35 ( .A(\ab[35][25] ), .B(\CARRYB[24][35] ), .CI(\SUMB[24][36] ), 
        .CO(\CARRYB[25][35] ), .S(\SUMB[25][35] ) );
  FA1P S4_29 ( .A(\ab[47][29] ), .B(\CARRYB[46][29] ), .CI(\SUMB[46][30] ), 
        .CO(\CARRYB[47][29] ), .S(\SUMB[47][29] ) );
  FA1 S2_28_34 ( .A(\ab[34][28] ), .B(\CARRYB[27][34] ), .CI(\SUMB[27][35] ), 
        .CO(\CARRYB[28][34] ), .S(\SUMB[28][34] ) );
  FA1AP S2_29_33 ( .A(\ab[33][29] ), .B(\CARRYB[28][33] ), .CI(\SUMB[28][34] ), 
        .CO(\CARRYB[29][33] ), .S(\SUMB[29][33] ) );
  FA1P S2_43_29 ( .A(\ab[43][29] ), .B(\CARRYB[42][29] ), .CI(\SUMB[42][30] ), 
        .CO(\CARRYB[43][29] ), .S(\SUMB[43][29] ) );
  FA1 S2_44_29 ( .A(\ab[44][29] ), .B(\CARRYB[43][29] ), .CI(\SUMB[43][30] ), 
        .CO(\CARRYB[44][29] ), .S(\SUMB[44][29] ) );
  FA1 S2_30_33 ( .A(\ab[33][30] ), .B(\CARRYB[29][33] ), .CI(\SUMB[29][34] ), 
        .CO(\CARRYB[30][33] ), .S(\SUMB[30][33] ) );
  FA1 S2_6_3 ( .A(n314), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1 S2_2_3 ( .A(n301), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1P S2_14_3 ( .A(n338), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), .CO(
        \CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1P S2_31_3 ( .A(n296), .B(\CARRYB[30][3] ), .CI(\SUMB[30][4] ), .CO(
        \CARRYB[31][3] ), .S(\SUMB[31][3] ) );
  FA1 S2_43_2 ( .A(n1302), .B(\CARRYB[42][2] ), .CI(\SUMB[42][3] ), .CO(
        \CARRYB[43][2] ), .S(\SUMB[43][2] ) );
  FA1AP S2_38_25 ( .A(\ab[38][25] ), .B(\CARRYB[37][25] ), .CI(\SUMB[37][26] ), 
        .CO(\CARRYB[38][25] ), .S(\SUMB[38][25] ) );
  FA1AP S2_31_27 ( .A(\ab[31][27] ), .B(\CARRYB[30][27] ), .CI(\SUMB[30][28] ), 
        .CO(\CARRYB[31][27] ), .S(\SUMB[31][27] ) );
  FA1P S4_24 ( .A(\ab[47][24] ), .B(\CARRYB[46][24] ), .CI(\SUMB[46][25] ), 
        .CO(\CARRYB[47][24] ), .S(\SUMB[47][24] ) );
  FA1P S4_23 ( .A(\ab[47][23] ), .B(\CARRYB[46][23] ), .CI(\SUMB[46][24] ), 
        .CO(\CARRYB[47][23] ), .S(\SUMB[47][23] ) );
  FA1 S2_37_16 ( .A(\ab[37][16] ), .B(\CARRYB[36][16] ), .CI(\SUMB[36][17] ), 
        .CO(\CARRYB[37][16] ), .S(\SUMB[37][16] ) );
  FA1P S2_35_16 ( .A(\ab[35][16] ), .B(\CARRYB[34][16] ), .CI(\SUMB[34][17] ), 
        .CO(\CARRYB[35][16] ), .S(\SUMB[35][16] ) );
  FA1P S2_36_16 ( .A(\ab[36][16] ), .B(\CARRYB[35][16] ), .CI(\SUMB[35][17] ), 
        .CO(\CARRYB[36][16] ), .S(\SUMB[36][16] ) );
  FA1P S2_15_21 ( .A(\ab[21][15] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA1P S2_2_15 ( .A(n1304), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1P S2_13_13 ( .A(\CARRYB[12][13] ), .B(A[13]), .CI(\SUMB[12][14] ), .CO(
        \CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1P S2_14_13 ( .A(n622), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), .CO(
        \CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1 S2_9_14 ( .A(n536), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1 S2_20_11 ( .A(n1322), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), .CO(
        \CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA1P S2_4_15 ( .A(n362), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), .CO(
        \CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1 S2_25_12 ( .A(n610), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), .CO(
        \CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA1P S2_27_7 ( .A(n423), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), .CO(
        \CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA1P S2_15_7 ( .A(n471), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1 S2_24_8 ( .A(n1291), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), .CO(
        \CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA1AP S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA1 S2_2_25 ( .A(n327), .B(\CARRYB[1][25] ), .CI(\SUMB[1][26] ), .CO(
        \CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA1 S2_27_16 ( .A(\SUMB[26][17] ), .B(\CARRYB[26][16] ), .CI(\ab[27][16] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA1AP S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA1A S2_41_12 ( .A(\ab[41][12] ), .B(\CARRYB[40][12] ), .CI(\SUMB[40][13] ), 
        .CO(\CARRYB[41][12] ), .S(\SUMB[41][12] ) );
  FA1AP S2_44_11 ( .A(\CARRYB[43][11] ), .B(\ab[44][11] ), .CI(\SUMB[43][12] ), 
        .CO(\CARRYB[44][11] ), .S(\SUMB[44][11] ) );
  FA1P S2_45_11 ( .A(\ab[45][11] ), .B(\CARRYB[44][11] ), .CI(\SUMB[44][12] ), 
        .CO(\CARRYB[45][11] ), .S(\SUMB[45][11] ) );
  FA1P S2_14_42 ( .A(\ab[42][14] ), .B(\CARRYB[13][42] ), .CI(\SUMB[13][43] ), 
        .CO(\CARRYB[14][42] ), .S(\SUMB[14][42] ) );
  FA1AP S2_30_41 ( .A(\ab[41][30] ), .B(\CARRYB[29][41] ), .CI(\SUMB[29][42] ), 
        .CO(\CARRYB[30][41] ), .S(\SUMB[30][41] ) );
  FA1P S2_43_39 ( .A(\ab[43][39] ), .B(\CARRYB[42][39] ), .CI(\SUMB[42][40] ), 
        .CO(\CARRYB[43][39] ), .S(\SUMB[43][39] ) );
  FA1P S2_44_39 ( .A(\ab[44][39] ), .B(\CARRYB[43][39] ), .CI(\SUMB[43][40] ), 
        .CO(\CARRYB[44][39] ), .S(\SUMB[44][39] ) );
  FA1P S2_46_39 ( .A(\ab[46][39] ), .B(\CARRYB[45][39] ), .CI(\SUMB[45][40] ), 
        .CO(\CARRYB[46][39] ), .S(\SUMB[46][39] ) );
  FA1AP S4_39 ( .A(\ab[47][39] ), .B(\CARRYB[46][39] ), .CI(\SUMB[46][40] ), 
        .CO(\CARRYB[47][39] ), .S(\SUMB[47][39] ) );
  FA1 S2_21_42 ( .A(\ab[42][21] ), .B(\CARRYB[20][42] ), .CI(\SUMB[20][43] ), 
        .CO(\CARRYB[21][42] ), .S(\SUMB[21][42] ) );
  FA1P S2_20_42 ( .A(\ab[42][20] ), .B(\CARRYB[19][42] ), .CI(\SUMB[19][43] ), 
        .CO(\CARRYB[20][42] ), .S(\SUMB[20][42] ) );
  FA1P S4_38 ( .A(\ab[47][38] ), .B(\CARRYB[46][38] ), .CI(\SUMB[46][39] ), 
        .CO(\CARRYB[47][38] ), .S(\SUMB[47][38] ) );
  FA1 S2_19_26 ( .A(\ab[26][19] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA1A S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), 
        .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FA1AP S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA1AP S2_20_25 ( .A(\ab[25][20] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA1 S2_41_19 ( .A(\ab[41][19] ), .B(\CARRYB[40][19] ), .CI(\SUMB[40][20] ), 
        .CO(\CARRYB[41][19] ), .S(\SUMB[41][19] ) );
  FA1P S2_41_20 ( .A(\ab[41][20] ), .B(\CARRYB[40][20] ), .CI(\SUMB[40][21] ), 
        .CO(\CARRYB[41][20] ), .S(\SUMB[41][20] ) );
  FA1P S2_21_40 ( .A(\ab[40][21] ), .B(\CARRYB[20][40] ), .CI(\SUMB[20][41] ), 
        .CO(\CARRYB[21][40] ), .S(\SUMB[21][40] ) );
  FA1P S2_17_40 ( .A(\ab[40][17] ), .B(\CARRYB[16][40] ), .CI(\SUMB[16][41] ), 
        .CO(\CARRYB[17][40] ), .S(\SUMB[17][40] ) );
  FA1P S2_18_40 ( .A(\ab[40][18] ), .B(\CARRYB[17][40] ), .CI(\SUMB[17][41] ), 
        .CO(\CARRYB[18][40] ), .S(\SUMB[18][40] ) );
  FA1P S2_28_40 ( .A(\ab[40][28] ), .B(\CARRYB[27][40] ), .CI(\SUMB[27][41] ), 
        .CO(\CARRYB[28][40] ), .S(\SUMB[28][40] ) );
  FA1P S2_24_40 ( .A(\ab[40][24] ), .B(\CARRYB[23][40] ), .CI(\SUMB[23][41] ), 
        .CO(\CARRYB[24][40] ), .S(\SUMB[24][40] ) );
  FA1AP S2_8_41 ( .A(n519), .B(\CARRYB[7][41] ), .CI(\SUMB[7][42] ), .CO(
        \CARRYB[8][41] ), .S(\SUMB[8][41] ) );
  FA1A S2_10_40 ( .A(\ab[40][10] ), .B(\CARRYB[9][40] ), .CI(\SUMB[9][41] ), 
        .CO(\CARRYB[10][40] ), .S(\SUMB[10][40] ) );
  FA1P S2_35_40 ( .A(\ab[40][35] ), .B(\CARRYB[34][40] ), .CI(\SUMB[34][41] ), 
        .CO(\CARRYB[35][40] ), .S(\SUMB[35][40] ) );
  FA1 S2_36_40 ( .A(\ab[40][36] ), .B(\CARRYB[35][40] ), .CI(\SUMB[35][41] ), 
        .CO(\CARRYB[36][40] ), .S(\SUMB[36][40] ) );
  FA1P S2_36_11 ( .A(\ab[36][11] ), .B(\CARRYB[35][11] ), .CI(\SUMB[35][12] ), 
        .CO(\CARRYB[36][11] ), .S(\SUMB[36][11] ) );
  FA1P S2_44_9 ( .A(\ab[9][44] ), .B(\CARRYB[43][9] ), .CI(\SUMB[43][10] ), 
        .CO(\CARRYB[44][9] ), .S(\SUMB[44][9] ) );
  FA1P S2_45_9 ( .A(\ab[9][45] ), .B(\CARRYB[44][9] ), .CI(\SUMB[44][10] ), 
        .CO(\CARRYB[45][9] ), .S(\SUMB[45][9] ) );
  FA1AP S2_37_11 ( .A(\ab[37][11] ), .B(\CARRYB[36][11] ), .CI(\SUMB[36][12] ), 
        .CO(\CARRYB[37][11] ), .S(\SUMB[37][11] ) );
  FA1P S2_38_11 ( .A(\ab[38][11] ), .B(\CARRYB[37][11] ), .CI(\SUMB[37][12] ), 
        .CO(\CARRYB[38][11] ), .S(\SUMB[38][11] ) );
  FA1P S4_8 ( .A(\ab[8][47] ), .B(\CARRYB[46][8] ), .CI(\SUMB[46][9] ), .CO(
        \CARRYB[47][8] ), .S(\SUMB[47][8] ) );
  FA1P S2_23_32 ( .A(\ab[32][23] ), .B(\CARRYB[22][32] ), .CI(\SUMB[22][33] ), 
        .CO(\CARRYB[23][32] ), .S(\SUMB[23][32] ) );
  FA1P S2_42_27 ( .A(\ab[42][27] ), .B(\CARRYB[41][27] ), .CI(\SUMB[41][28] ), 
        .CO(\CARRYB[42][27] ), .S(\SUMB[42][27] ) );
  FA1 S2_40_27 ( .A(\ab[40][27] ), .B(\CARRYB[39][27] ), .CI(\SUMB[39][28] ), 
        .CO(\CARRYB[40][27] ), .S(\SUMB[40][27] ) );
  FA1P S2_41_27 ( .A(\ab[41][27] ), .B(\CARRYB[40][27] ), .CI(\SUMB[40][28] ), 
        .CO(\CARRYB[41][27] ), .S(\SUMB[41][27] ) );
  FA1P S2_3_21 ( .A(n330), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), .CO(
        \CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA1P S2_19_13 ( .A(n630), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), .CO(
        \CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA1AP S2_5_20 ( .A(\CARRYB[4][20] ), .B(n383), .CI(\SUMB[4][21] ), .CO(
        \CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1P S2_39_7 ( .A(n475), .B(\CARRYB[38][7] ), .CI(\SUMB[38][8] ), .CO(
        \CARRYB[39][7] ), .S(\SUMB[39][7] ) );
  FA1AP S2_13_4 ( .A(n391), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), .CO(
        \CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1P S2_24_2 ( .A(n1300), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), .CO(
        \CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA1P S2_25_2 ( .A(n327), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), .CO(
        \CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA1P S2_19_3 ( .A(n329), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), .CO(
        \CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1P S2_20_3 ( .A(n1379), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), .CO(
        \CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1P S2_29_1 ( .A(n1324), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), .CO(
        \CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA1P S2_2_5 ( .A(n359), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1P S2_3_5 ( .A(n324), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1AP S2_29_34 ( .A(\ab[34][29] ), .B(\CARRYB[28][34] ), .CI(\SUMB[28][35] ), 
        .CO(\CARRYB[29][34] ), .S(\SUMB[29][34] ) );
  FA1P S2_34_33 ( .A(\ab[34][33] ), .B(\CARRYB[33][33] ), .CI(\SUMB[33][34] ), 
        .CO(\CARRYB[34][33] ), .S(\SUMB[34][33] ) );
  FA1P S2_36_33 ( .A(\ab[36][33] ), .B(\CARRYB[35][33] ), .CI(\SUMB[35][34] ), 
        .CO(\CARRYB[36][33] ), .S(\SUMB[36][33] ) );
  FA1P S2_33_33 ( .A(A[33]), .B(\CARRYB[32][33] ), .CI(\SUMB[32][34] ), .CO(
        \CARRYB[33][33] ), .S(\SUMB[33][33] ) );
  FA1AP S2_14_30 ( .A(\ab[30][14] ), .B(\CARRYB[13][30] ), .CI(\SUMB[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA1P S2_42_21 ( .A(\ab[42][21] ), .B(\CARRYB[41][21] ), .CI(\SUMB[41][22] ), 
        .CO(\CARRYB[42][21] ), .S(\SUMB[42][21] ) );
  FA1P S4_18 ( .A(\ab[47][18] ), .B(\CARRYB[46][18] ), .CI(\SUMB[46][19] ), 
        .CO(\CARRYB[47][18] ), .S(\SUMB[47][18] ) );
  FA1 S2_14_24 ( .A(n640), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), .CO(
        \CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA1 S2_23_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA1AP S2_32_33 ( .A(\ab[33][32] ), .B(\CARRYB[31][33] ), .CI(\SUMB[31][34] ), 
        .CO(\CARRYB[32][33] ), .S(\SUMB[32][33] ) );
  FA1P S2_45_28 ( .A(\ab[45][28] ), .B(\CARRYB[44][28] ), .CI(\SUMB[44][29] ), 
        .CO(\CARRYB[45][28] ), .S(\SUMB[45][28] ) );
  FA1 S2_21_23 ( .A(\ab[23][21] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA1AP S2_22_23 ( .A(\CARRYB[21][23] ), .B(\ab[23][22] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA1P S2_42_17 ( .A(\ab[42][17] ), .B(\CARRYB[41][17] ), .CI(\SUMB[41][18] ), 
        .CO(\CARRYB[42][17] ), .S(\SUMB[42][17] ) );
  FA1P S2_19_20 ( .A(\ab[20][19] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA1A S1_25_0 ( .A(n1399), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), .CO(
        \CARRYB[25][0] ), .S(\A1[23] ) );
  FA1 S2_46_21 ( .A(\ab[46][21] ), .B(\CARRYB[45][21] ), .CI(\SUMB[45][22] ), 
        .CO(\CARRYB[46][21] ), .S(\SUMB[46][21] ) );
  FA1AP S2_11_22 ( .A(n565), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), .CO(
        \CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA1P S2_43_8 ( .A(n511), .B(\CARRYB[42][8] ), .CI(\SUMB[42][9] ), .CO(
        \CARRYB[43][8] ), .S(\SUMB[43][8] ) );
  FA1P S2_44_8 ( .A(\ab[8][44] ), .B(\CARRYB[43][8] ), .CI(\SUMB[43][9] ), 
        .CO(\CARRYB[44][8] ), .S(\SUMB[44][8] ) );
  FA1P S2_38_10 ( .A(\ab[38][10] ), .B(\CARRYB[37][10] ), .CI(\SUMB[37][11] ), 
        .CO(\CARRYB[38][10] ), .S(\SUMB[38][10] ) );
  FA1AP S2_8_23 ( .A(n499), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), .CO(
        \CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA1P S2_12_22 ( .A(\CARRYB[11][22] ), .B(n594), .CI(\SUMB[11][23] ), .CO(
        \CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA1A S1_42_0 ( .A(n1350), .B(\CARRYB[41][0] ), .CI(\SUMB[41][1] ), .CO(
        \CARRYB[42][0] ), .S(\A1[40] ) );
  FA1 S1_11_0 ( .A(n1371), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(
        \CARRYB[11][0] ), .S(\A1[9] ) );
  FA1P S1_29_0 ( .A(n1366), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), .CO(
        \CARRYB[29][0] ), .S(\A1[27] ) );
  FA1 S1_24_0 ( .A(n1325), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), .CO(
        \CARRYB[24][0] ), .S(\A1[22] ) );
  FA1 S1_41_0 ( .A(n1373), .B(\CARRYB[40][0] ), .CI(\SUMB[40][1] ), .CO(
        \CARRYB[41][0] ), .S(\A1[39] ) );
  FA1 S2_38_1 ( .A(n1369), .B(\CARRYB[37][1] ), .CI(\SUMB[37][2] ), .CO(
        \CARRYB[38][1] ), .S(\SUMB[38][1] ) );
  FA1 S1_3_0 ( .A(n1531), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1P S2_5_13 ( .A(n421), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), .CO(
        \CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1 S2_6_13 ( .A(n450), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), .CO(
        \CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1 S2_15_9 ( .A(n527), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), .CO(
        \CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1P S2_34_4 ( .A(n352), .B(\CARRYB[33][4] ), .CI(\SUMB[33][5] ), .CO(
        \CARRYB[34][4] ), .S(\SUMB[34][4] ) );
  FA1P S2_7_12 ( .A(n510), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), .CO(
        \CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1 S2_8_12 ( .A(n538), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), .CO(
        \CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1AP S2_26_7 ( .A(n472), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), .CO(
        \CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA1A S2_10_31 ( .A(\CARRYB[9][31] ), .B(n545), .CI(\SUMB[9][32] ), .CO(
        \CARRYB[10][31] ), .S(\SUMB[10][31] ) );
  FA1P S2_2_33 ( .A(n1306), .B(\CARRYB[1][33] ), .CI(\SUMB[1][34] ), .CO(
        \CARRYB[2][33] ), .S(\SUMB[2][33] ) );
  FA1AP S2_24_34 ( .A(\ab[34][24] ), .B(\CARRYB[23][34] ), .CI(\SUMB[23][35] ), 
        .CO(\CARRYB[24][34] ), .S(\SUMB[24][34] ) );
  FA1AP S2_41_24 ( .A(\CARRYB[40][24] ), .B(\ab[41][24] ), .CI(\SUMB[40][25] ), 
        .CO(\CARRYB[41][24] ), .S(\SUMB[41][24] ) );
  FA1AP S2_22_34 ( .A(\ab[34][22] ), .B(\CARRYB[21][34] ), .CI(\SUMB[21][35] ), 
        .CO(\CARRYB[22][34] ), .S(\SUMB[22][34] ) );
  FA1P S2_38_31 ( .A(\ab[38][31] ), .B(\CARRYB[37][31] ), .CI(\SUMB[37][32] ), 
        .CO(\CARRYB[38][31] ), .S(\SUMB[38][31] ) );
  FA1P S2_36_32 ( .A(\ab[36][32] ), .B(\CARRYB[35][32] ), .CI(\SUMB[35][33] ), 
        .CO(\CARRYB[36][32] ), .S(\SUMB[36][32] ) );
  FA1P S2_44_31 ( .A(\ab[44][31] ), .B(\CARRYB[43][31] ), .CI(\SUMB[43][32] ), 
        .CO(\CARRYB[44][31] ), .S(\SUMB[44][31] ) );
  FA1AP S2_7_26 ( .A(n472), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), .CO(
        \CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA1P S2_12_24 ( .A(n593), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), .CO(
        \CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA1AP S2_20_20 ( .A(A[20]), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), .CO(
        \CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA1P S2_24_44 ( .A(\ab[44][24] ), .B(\CARRYB[23][44] ), .CI(\SUMB[23][45] ), 
        .CO(\CARRYB[24][44] ), .S(\SUMB[24][44] ) );
  FA1P S2_25_44 ( .A(\ab[44][25] ), .B(\CARRYB[24][44] ), .CI(\SUMB[24][45] ), 
        .CO(\CARRYB[25][44] ), .S(\SUMB[25][44] ) );
  FA1 S2_37_44 ( .A(\ab[44][37] ), .B(\CARRYB[36][44] ), .CI(\SUMB[36][45] ), 
        .CO(\CARRYB[37][44] ), .S(\SUMB[37][44] ) );
  FA1P S2_45_42 ( .A(\ab[45][42] ), .B(\CARRYB[44][42] ), .CI(\SUMB[44][43] ), 
        .CO(\CARRYB[45][42] ), .S(\SUMB[45][42] ) );
  FA1P S2_45_43 ( .A(\ab[45][43] ), .B(\CARRYB[44][43] ), .CI(\SUMB[44][44] ), 
        .CO(\CARRYB[45][43] ), .S(\SUMB[45][43] ) );
  FA1P S2_22_44 ( .A(\ab[44][22] ), .B(\CARRYB[21][44] ), .CI(\SUMB[21][45] ), 
        .CO(\CARRYB[22][44] ), .S(\SUMB[22][44] ) );
  FA1P S2_39_44 ( .A(\ab[44][39] ), .B(\CARRYB[38][44] ), .CI(\SUMB[38][45] ), 
        .CO(\CARRYB[39][44] ), .S(\SUMB[39][44] ) );
  FA1P S2_40_43 ( .A(\ab[43][40] ), .B(\CARRYB[39][43] ), .CI(\SUMB[39][44] ), 
        .CO(\CARRYB[40][43] ), .S(\SUMB[40][43] ) );
  FA1 S2_24_33 ( .A(\ab[33][24] ), .B(\CARRYB[23][33] ), .CI(\SUMB[23][34] ), 
        .CO(\CARRYB[24][33] ), .S(\SUMB[24][33] ) );
  FA1AP S2_28_32 ( .A(\ab[32][28] ), .B(\CARRYB[27][32] ), .CI(\SUMB[27][33] ), 
        .CO(\CARRYB[28][32] ), .S(\SUMB[28][32] ) );
  FA1 S2_28_33 ( .A(\ab[33][28] ), .B(\CARRYB[27][33] ), .CI(\SUMB[27][34] ), 
        .CO(\CARRYB[28][33] ), .S(\SUMB[28][33] ) );
  FA1 S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA1AP S2_35_15 ( .A(\ab[35][15] ), .B(\CARRYB[34][15] ), .CI(\SUMB[34][16] ), 
        .CO(\CARRYB[35][15] ), .S(\SUMB[35][15] ) );
  FA1P S2_13_23 ( .A(n619), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), .CO(
        \CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA1P S2_14_23 ( .A(n642), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), .CO(
        \CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA1 S2_46_11 ( .A(\ab[46][11] ), .B(\CARRYB[45][11] ), .CI(\SUMB[45][12] ), 
        .CO(\CARRYB[46][11] ), .S(\SUMB[46][11] ) );
  FA1AP S4_11 ( .A(\ab[47][11] ), .B(\CARRYB[46][11] ), .CI(\SUMB[46][12] ), 
        .CO(\CARRYB[47][11] ), .S(\SUMB[47][11] ) );
  FA1 S2_6_26 ( .A(n433), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), .CO(
        \CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA1A S2_7_25 ( .A(n419), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), .CO(
        \CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA1AP S2_18_33 ( .A(\ab[33][18] ), .B(\CARRYB[17][33] ), .CI(\SUMB[17][34] ), 
        .CO(\CARRYB[18][33] ), .S(\SUMB[18][33] ) );
  FA1 S2_39_24 ( .A(\ab[39][24] ), .B(\CARRYB[38][24] ), .CI(\SUMB[38][25] ), 
        .CO(\CARRYB[39][24] ), .S(\SUMB[39][24] ) );
  FA1A S2_42_28 ( .A(\ab[42][28] ), .B(\CARRYB[41][28] ), .CI(\SUMB[41][29] ), 
        .CO(\CARRYB[42][28] ), .S(\SUMB[42][28] ) );
  FA1P S2_42_29 ( .A(\ab[42][29] ), .B(\CARRYB[41][29] ), .CI(\SUMB[41][30] ), 
        .CO(\CARRYB[42][29] ), .S(\SUMB[42][29] ) );
  FA1P S2_44_28 ( .A(\ab[44][28] ), .B(\CARRYB[43][28] ), .CI(\SUMB[43][29] ), 
        .CO(\CARRYB[44][28] ), .S(\SUMB[44][28] ) );
  FA1P S2_41_23 ( .A(\ab[41][23] ), .B(\CARRYB[40][23] ), .CI(\SUMB[40][24] ), 
        .CO(\CARRYB[41][23] ), .S(\SUMB[41][23] ) );
  FA1 S2_42_23 ( .A(\ab[42][23] ), .B(\CARRYB[41][23] ), .CI(\SUMB[41][24] ), 
        .CO(\CARRYB[42][23] ), .S(\SUMB[42][23] ) );
  FA1A S2_16_32 ( .A(\ab[32][16] ), .B(\CARRYB[15][32] ), .CI(\SUMB[15][33] ), 
        .CO(\CARRYB[16][32] ), .S(\SUMB[16][32] ) );
  FA1P S2_23_12 ( .A(n600), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), .CO(
        \CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA1 S2_33_9 ( .A(n516), .B(\CARRYB[32][9] ), .CI(\SUMB[32][10] ), .CO(
        \CARRYB[33][9] ), .S(\SUMB[33][9] ) );
  FA1P S2_41_6 ( .A(n443), .B(\CARRYB[40][6] ), .CI(\SUMB[40][7] ), .CO(
        \CARRYB[41][6] ), .S(\SUMB[41][6] ) );
  FA1 S2_16_7 ( .A(n479), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), .CO(
        \CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1 S2_3_9 ( .A(n347), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_24_7 ( .A(n1285), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), .CO(
        \CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA1 S2_44_3 ( .A(n341), .B(\CARRYB[43][3] ), .CI(\SUMB[43][4] ), .CO(
        \CARRYB[44][3] ), .S(\SUMB[44][3] ) );
  FA1 S2_13_33 ( .A(\ab[33][13] ), .B(\CARRYB[12][33] ), .CI(\SUMB[12][34] ), 
        .CO(\CARRYB[13][33] ), .S(\SUMB[13][33] ) );
  FA1P S2_15_33 ( .A(\ab[33][15] ), .B(\CARRYB[14][33] ), .CI(\SUMB[14][34] ), 
        .CO(\CARRYB[15][33] ), .S(\SUMB[15][33] ) );
  FA1 S2_6_36 ( .A(n436), .B(\CARRYB[5][36] ), .CI(\SUMB[5][37] ), .CO(
        \CARRYB[6][36] ), .S(\SUMB[6][36] ) );
  FA1 S2_32_27 ( .A(\ab[32][27] ), .B(\CARRYB[31][27] ), .CI(\SUMB[31][28] ), 
        .CO(\CARRYB[32][27] ), .S(\SUMB[32][27] ) );
  FA1AP S2_33_27 ( .A(\ab[33][27] ), .B(\CARRYB[32][27] ), .CI(\SUMB[32][28] ), 
        .CO(\CARRYB[33][27] ), .S(\SUMB[33][27] ) );
  FA1 S2_13_36 ( .A(\CARRYB[12][36] ), .B(\ab[36][13] ), .CI(\SUMB[12][37] ), 
        .CO(\CARRYB[13][36] ), .S(\SUMB[13][36] ) );
  FA1A S2_35_25 ( .A(\ab[35][25] ), .B(\CARRYB[34][25] ), .CI(\SUMB[34][26] ), 
        .CO(\CARRYB[35][25] ), .S(\SUMB[35][25] ) );
  FA1P S2_3_31 ( .A(n296), .B(\CARRYB[2][31] ), .CI(\SUMB[2][32] ), .CO(
        \CARRYB[3][31] ), .S(\SUMB[3][31] ) );
  FA1 S2_17_28 ( .A(\ab[28][17] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA1P S2_46_18 ( .A(\ab[46][18] ), .B(\CARRYB[45][18] ), .CI(\SUMB[45][19] ), 
        .CO(\CARRYB[46][18] ), .S(\SUMB[46][18] ) );
  FA1AP S2_39_22 ( .A(\CARRYB[38][22] ), .B(\ab[39][22] ), .CI(\SUMB[38][23] ), 
        .CO(\CARRYB[39][22] ), .S(\SUMB[39][22] ) );
  FA1AP S2_5_28 ( .A(n393), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), .CO(
        \CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA1AP S2_38_18 ( .A(\ab[38][18] ), .B(\CARRYB[37][18] ), .CI(\SUMB[37][19] ), 
        .CO(\CARRYB[38][18] ), .S(\SUMB[38][18] ) );
  FA1P S2_39_18 ( .A(\ab[39][18] ), .B(\CARRYB[38][18] ), .CI(\SUMB[38][19] ), 
        .CO(\CARRYB[39][18] ), .S(\SUMB[39][18] ) );
  FA1 S2_34_26 ( .A(\ab[34][26] ), .B(\CARRYB[33][26] ), .CI(\SUMB[33][27] ), 
        .CO(\CARRYB[34][26] ), .S(\SUMB[34][26] ) );
  FA1 S2_32_26 ( .A(\ab[32][26] ), .B(\CARRYB[31][26] ), .CI(\SUMB[31][27] ), 
        .CO(\CARRYB[32][26] ), .S(\SUMB[32][26] ) );
  FA1AP S2_33_26 ( .A(\ab[33][26] ), .B(\CARRYB[32][26] ), .CI(\SUMB[32][27] ), 
        .CO(\CARRYB[33][26] ), .S(\SUMB[33][26] ) );
  FA1AP S2_30_21 ( .A(\ab[30][21] ), .B(\CARRYB[29][21] ), .CI(\SUMB[29][22] ), 
        .CO(\CARRYB[30][21] ), .S(\SUMB[30][21] ) );
  FA1P S2_31_21 ( .A(\ab[31][21] ), .B(\CARRYB[30][21] ), .CI(\SUMB[30][22] ), 
        .CO(\CARRYB[31][21] ), .S(\SUMB[31][21] ) );
  FA1P S2_33_21 ( .A(\ab[33][21] ), .B(\CARRYB[32][21] ), .CI(\SUMB[32][22] ), 
        .CO(\CARRYB[33][21] ), .S(\SUMB[33][21] ) );
  FA1AP S2_26_22 ( .A(\CARRYB[25][22] ), .B(\ab[26][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA1A S2_7_28 ( .A(n424), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), .CO(
        \CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA1P S2_13_32 ( .A(\ab[32][13] ), .B(\CARRYB[12][32] ), .CI(\SUMB[12][33] ), 
        .CO(\CARRYB[13][32] ), .S(\SUMB[13][32] ) );
  FA1AP S2_35_26 ( .A(\ab[35][26] ), .B(\CARRYB[34][26] ), .CI(\SUMB[34][27] ), 
        .CO(\CARRYB[35][26] ), .S(\SUMB[35][26] ) );
  FA1 S2_30_28 ( .A(\CARRYB[29][28] ), .B(\ab[30][28] ), .CI(\SUMB[29][29] ), 
        .CO(\CARRYB[30][28] ), .S(\SUMB[30][28] ) );
  FA1P S2_3_7 ( .A(\CARRYB[2][7] ), .B(n345), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_34_2 ( .A(n1307), .B(\CARRYB[33][2] ), .CI(\SUMB[33][3] ), .CO(
        \CARRYB[34][2] ), .S(\SUMB[34][2] ) );
  FA1P S2_35_2 ( .A(n1316), .B(\CARRYB[34][2] ), .CI(\SUMB[34][3] ), .CO(
        \CARRYB[35][2] ), .S(\SUMB[35][2] ) );
  FA1P S2_16_4 ( .A(n361), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), .CO(
        \CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1P S2_26_4 ( .A(n364), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), .CO(
        \CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA1P S2_7_5 ( .A(n426), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1AP S2_28_4 ( .A(n351), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), .CO(
        \CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA1P S2_45_2 ( .A(n1314), .B(\CARRYB[44][2] ), .CI(\SUMB[44][3] ), .CO(
        \CARRYB[45][2] ), .S(\SUMB[45][2] ) );
  FA1P S2_38_35 ( .A(\ab[38][35] ), .B(\CARRYB[37][35] ), .CI(\SUMB[37][36] ), 
        .CO(\CARRYB[38][35] ), .S(\SUMB[38][35] ) );
  FA1P S2_29_38 ( .A(\ab[38][29] ), .B(\CARRYB[28][38] ), .CI(\SUMB[28][39] ), 
        .CO(\CARRYB[29][38] ), .S(\SUMB[29][38] ) );
  FA1P S4_33 ( .A(\ab[47][33] ), .B(\CARRYB[46][33] ), .CI(\SUMB[46][34] ), 
        .CO(\CARRYB[47][33] ), .S(\SUMB[47][33] ) );
  FA1P S2_21_38 ( .A(\ab[38][21] ), .B(\CARRYB[20][38] ), .CI(\SUMB[20][39] ), 
        .CO(\CARRYB[21][38] ), .S(\SUMB[21][38] ) );
  FA1P S2_19_38 ( .A(\ab[38][19] ), .B(\SUMB[18][39] ), .CI(\CARRYB[18][38] ), 
        .CO(\CARRYB[19][38] ), .S(\SUMB[19][38] ) );
  FA1P S2_20_38 ( .A(\ab[38][20] ), .B(\CARRYB[19][38] ), .CI(\SUMB[19][39] ), 
        .CO(\CARRYB[20][38] ), .S(\SUMB[20][38] ) );
  FA1P S2_40_6 ( .A(n387), .B(\CARRYB[39][6] ), .CI(\SUMB[39][7] ), .CO(
        \CARRYB[40][6] ), .S(\SUMB[40][6] ) );
  FA1 S2_2_20 ( .A(n1341), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), .CO(
        \CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1AP S2_8_19 ( .A(n484), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), .CO(
        \CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA1AP S2_31_28 ( .A(\ab[31][28] ), .B(\CARRYB[30][28] ), .CI(\SUMB[30][29] ), 
        .CO(\CARRYB[31][28] ), .S(\SUMB[31][28] ) );
  FA1P S2_22_25 ( .A(\ab[25][22] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA1 S2_11_28 ( .A(n562), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), .CO(
        \CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA1AP S2_12_27 ( .A(n603), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), .CO(
        \CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA1A S2_12_34 ( .A(\ab[34][12] ), .B(\CARRYB[11][34] ), .CI(\SUMB[11][35] ), 
        .CO(\CARRYB[12][34] ), .S(\SUMB[12][34] ) );
  FA1 S2_17_18 ( .A(\ab[18][17] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA1AP S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA1AP S2_9_22 ( .A(n280), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), .CO(
        \CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA1AP S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA1 S2_31_14 ( .A(\ab[31][14] ), .B(\CARRYB[30][14] ), .CI(\SUMB[30][15] ), 
        .CO(\CARRYB[31][14] ), .S(\SUMB[31][14] ) );
  FA1P S2_40_11 ( .A(\CARRYB[39][11] ), .B(\ab[40][11] ), .CI(\SUMB[39][12] ), 
        .CO(\CARRYB[40][11] ), .S(\SUMB[40][11] ) );
  FA1 S2_29_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA1A S2_6_23 ( .A(n422), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), .CO(
        \CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA1 S2_10_16 ( .A(n559), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), .CO(
        \CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1P S2_4_17 ( .A(n1278), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), .CO(
        \CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1AP S2_5_17 ( .A(n1284), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), .CO(
        \CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1P S2_38_7 ( .A(n1288), .B(\CARRYB[37][7] ), .CI(\SUMB[37][8] ), .CO(
        \CARRYB[38][7] ), .S(\SUMB[38][7] ) );
  FA1P S2_13_34 ( .A(\ab[34][13] ), .B(\CARRYB[12][34] ), .CI(\SUMB[12][35] ), 
        .CO(\CARRYB[13][34] ), .S(\SUMB[13][34] ) );
  FA1P S2_45_23 ( .A(\ab[45][23] ), .B(\CARRYB[44][23] ), .CI(\SUMB[44][24] ), 
        .CO(\CARRYB[45][23] ), .S(\SUMB[45][23] ) );
  FA1A S2_46_22 ( .A(\CARRYB[45][22] ), .B(\ab[46][22] ), .CI(\SUMB[45][23] ), 
        .CO(\CARRYB[46][22] ), .S(\SUMB[46][22] ) );
  FA1A S2_17_21 ( .A(\ab[21][17] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA1AP S2_18_21 ( .A(\ab[21][18] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA1AP S2_40_14 ( .A(\ab[40][14] ), .B(\CARRYB[39][14] ), .CI(\SUMB[39][15] ), 
        .CO(\CARRYB[40][14] ), .S(\SUMB[40][14] ) );
  FA1 S2_41_14 ( .A(\ab[41][14] ), .B(\CARRYB[40][14] ), .CI(\SUMB[40][15] ), 
        .CO(\CARRYB[41][14] ), .S(\SUMB[41][14] ) );
  FA1A S2_11_25 ( .A(n563), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), .CO(
        \CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA1P S2_19_43 ( .A(\ab[43][19] ), .B(\CARRYB[18][43] ), .CI(\SUMB[18][44] ), 
        .CO(\CARRYB[19][43] ), .S(\SUMB[19][43] ) );
  FA1 S2_43_37 ( .A(\ab[43][37] ), .B(\CARRYB[42][37] ), .CI(\SUMB[42][38] ), 
        .CO(\CARRYB[43][37] ), .S(\SUMB[43][37] ) );
  FA1A S2_34_39 ( .A(\ab[39][34] ), .B(\CARRYB[33][39] ), .CI(\SUMB[33][40] ), 
        .CO(\CARRYB[34][39] ), .S(\SUMB[34][39] ) );
  FA1 S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA1AP S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA1A S2_44_19 ( .A(\ab[44][19] ), .B(\CARRYB[43][19] ), .CI(\SUMB[43][20] ), 
        .CO(\CARRYB[44][19] ), .S(\SUMB[44][19] ) );
  FA1AP S2_5_33 ( .A(n386), .B(\CARRYB[4][33] ), .CI(\SUMB[4][34] ), .CO(
        \CARRYB[5][33] ), .S(\SUMB[5][33] ) );
  FA1P S2_39_30 ( .A(\ab[39][30] ), .B(\CARRYB[38][30] ), .CI(\SUMB[38][31] ), 
        .CO(\CARRYB[39][30] ), .S(\SUMB[39][30] ) );
  FA1AP S2_31_33 ( .A(\ab[33][31] ), .B(\CARRYB[30][33] ), .CI(\SUMB[30][34] ), 
        .CO(\CARRYB[31][33] ), .S(\SUMB[31][33] ) );
  FA1 S2_26_35 ( .A(\ab[35][26] ), .B(\CARRYB[25][35] ), .CI(\SUMB[25][36] ), 
        .CO(\CARRYB[26][35] ), .S(\SUMB[26][35] ) );
  FA1A S2_27_35 ( .A(\ab[35][27] ), .B(\CARRYB[26][35] ), .CI(\SUMB[26][36] ), 
        .CO(\CARRYB[27][35] ), .S(\SUMB[27][35] ) );
  FA1P S2_41_17 ( .A(\ab[41][17] ), .B(\CARRYB[40][17] ), .CI(\SUMB[40][18] ), 
        .CO(\CARRYB[41][17] ), .S(\SUMB[41][17] ) );
  FA1A S2_34_19 ( .A(\ab[34][19] ), .B(\CARRYB[33][19] ), .CI(\SUMB[33][20] ), 
        .CO(\CARRYB[34][19] ), .S(\SUMB[34][19] ) );
  FA1P S2_22_12 ( .A(n594), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), .CO(
        \CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA1A S2_34_9 ( .A(n539), .B(\CARRYB[33][9] ), .CI(\SUMB[33][10] ), .CO(
        \CARRYB[34][9] ), .S(\SUMB[34][9] ) );
  FA1P S2_10_29 ( .A(n555), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), .CO(
        \CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA1 S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA1A S2_42_18 ( .A(\ab[42][18] ), .B(\CARRYB[41][18] ), .CI(\SUMB[41][19] ), 
        .CO(\CARRYB[42][18] ), .S(\SUMB[42][18] ) );
  FA1P S2_40_26 ( .A(\ab[40][26] ), .B(\CARRYB[39][26] ), .CI(\SUMB[39][27] ), 
        .CO(\CARRYB[40][26] ), .S(\SUMB[40][26] ) );
  FA1P S2_41_26 ( .A(\ab[41][26] ), .B(\CARRYB[40][26] ), .CI(\SUMB[40][27] ), 
        .CO(\CARRYB[41][26] ), .S(\SUMB[41][26] ) );
  FA1AP S2_26_33 ( .A(\ab[33][26] ), .B(\CARRYB[25][33] ), .CI(\SUMB[25][34] ), 
        .CO(\CARRYB[26][33] ), .S(\SUMB[26][33] ) );
  FA1A S2_31_29 ( .A(\ab[31][29] ), .B(\CARRYB[30][29] ), .CI(\SUMB[30][30] ), 
        .CO(\CARRYB[31][29] ), .S(\SUMB[31][29] ) );
  FA1 S2_12_16 ( .A(n612), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), .CO(
        \CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA1P S2_2_21 ( .A(n1305), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), .CO(
        \CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA1 S2_42_9 ( .A(\ab[9][42] ), .B(\CARRYB[41][9] ), .CI(\SUMB[41][10] ), 
        .CO(\CARRYB[42][9] ), .S(\SUMB[42][9] ) );
  FA1P S2_46_8 ( .A(\ab[8][46] ), .B(\CARRYB[45][8] ), .CI(\SUMB[45][9] ), 
        .CO(\CARRYB[46][8] ), .S(\SUMB[46][8] ) );
  FA1P S2_16_19 ( .A(\ab[19][16] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA1AP S2_24_15 ( .A(\CARRYB[23][15] ), .B(\ab[24][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA1P S2_16_41 ( .A(\ab[41][16] ), .B(\CARRYB[15][41] ), .CI(\SUMB[15][42] ), 
        .CO(\CARRYB[16][41] ), .S(\SUMB[16][41] ) );
  FA1P S2_34_38 ( .A(\ab[38][34] ), .B(\CARRYB[33][38] ), .CI(\SUMB[33][39] ), 
        .CO(\CARRYB[34][38] ), .S(\SUMB[34][38] ) );
  FA1 S2_41_37 ( .A(\ab[41][37] ), .B(\CARRYB[40][37] ), .CI(\SUMB[40][38] ), 
        .CO(\CARRYB[41][37] ), .S(\SUMB[41][37] ) );
  FA1 S2_23_39 ( .A(\ab[39][23] ), .B(\CARRYB[22][39] ), .CI(\SUMB[22][40] ), 
        .CO(\CARRYB[23][39] ), .S(\SUMB[23][39] ) );
  FA1P S2_30_38 ( .A(\ab[38][30] ), .B(\CARRYB[29][38] ), .CI(\SUMB[29][39] ), 
        .CO(\CARRYB[30][38] ), .S(\SUMB[30][38] ) );
  FA1A S2_30_39 ( .A(\ab[39][30] ), .B(\CARRYB[29][39] ), .CI(\SUMB[29][40] ), 
        .CO(\CARRYB[30][39] ), .S(\SUMB[30][39] ) );
  FA1P S2_44_37 ( .A(\ab[44][37] ), .B(\CARRYB[43][37] ), .CI(\SUMB[43][38] ), 
        .CO(\CARRYB[44][37] ), .S(\SUMB[44][37] ) );
  FA1 S2_45_37 ( .A(\ab[45][37] ), .B(\CARRYB[44][37] ), .CI(\SUMB[44][38] ), 
        .CO(\CARRYB[45][37] ), .S(\SUMB[45][37] ) );
  FA1P S2_19_7 ( .A(n451), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), .CO(
        \CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA1P S2_20_7 ( .A(n458), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), .CO(
        \CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1P S2_37_3 ( .A(n283), .B(\CARRYB[36][3] ), .CI(\SUMB[36][4] ), .CO(
        \CARRYB[37][3] ), .S(\SUMB[37][3] ) );
  FA1P S2_4_8 ( .A(n372), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1P S2_5_8 ( .A(n425), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1P S2_10_7 ( .A(n503), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_6_8 ( .A(n456), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1 S2_7_8 ( .A(n493), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1P S2_2_37 ( .A(n309), .B(\CARRYB[1][37] ), .CI(\SUMB[1][38] ), .CO(
        \CARRYB[2][37] ), .S(\SUMB[2][37] ) );
  FA1 S2_36_25 ( .A(\ab[36][25] ), .B(\CARRYB[35][25] ), .CI(\SUMB[35][26] ), 
        .CO(\CARRYB[36][25] ), .S(\SUMB[36][25] ) );
  FA1 S2_20_9 ( .A(n525), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), .CO(
        \CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1P S2_21_9 ( .A(n512), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), .CO(
        \CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1AP S2_10_13 ( .A(n566), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), .CO(
        \CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1P S2_23_8 ( .A(n499), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), .CO(
        \CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA1P S2_3_18 ( .A(n1391), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), .CO(
        \CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1P S2_4_18 ( .A(n350), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), .CO(
        \CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1AP S2_6_39 ( .A(n432), .B(\CARRYB[5][39] ), .CI(\SUMB[5][40] ), .CO(
        \CARRYB[6][39] ), .S(\SUMB[6][39] ) );
  FA1P S2_13_27 ( .A(n613), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), .CO(
        \CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA1 S2_37_20 ( .A(\ab[37][20] ), .B(\CARRYB[36][20] ), .CI(\SUMB[36][21] ), 
        .CO(\CARRYB[37][20] ), .S(\SUMB[37][20] ) );
  FA1 S2_37_19 ( .A(\ab[37][19] ), .B(\CARRYB[36][19] ), .CI(\SUMB[36][20] ), 
        .CO(\CARRYB[37][19] ), .S(\SUMB[37][19] ) );
  FA1AP S2_3_27 ( .A(n292), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), .CO(
        \CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA1 S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA1AP S2_33_15 ( .A(\ab[33][15] ), .B(\CARRYB[32][15] ), .CI(\SUMB[32][16] ), 
        .CO(\CARRYB[33][15] ), .S(\SUMB[33][15] ) );
  FA1A S1_30_0 ( .A(n1396), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), .CO(
        \CARRYB[30][0] ), .S(\A1[28] ) );
  FA1P S2_42_11 ( .A(\ab[42][11] ), .B(\CARRYB[41][11] ), .CI(\SUMB[41][12] ), 
        .CO(\CARRYB[42][11] ), .S(\SUMB[42][11] ) );
  FA1 S2_43_11 ( .A(\ab[43][11] ), .B(\CARRYB[42][11] ), .CI(\SUMB[42][12] ), 
        .CO(\CARRYB[43][11] ), .S(\SUMB[43][11] ) );
  FA1A S2_20_24 ( .A(\ab[24][20] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA1P S2_44_17 ( .A(\ab[44][17] ), .B(\CARRYB[43][17] ), .CI(\SUMB[43][18] ), 
        .CO(\CARRYB[44][17] ), .S(\SUMB[44][17] ) );
  FA1AP S2_39_17 ( .A(\ab[39][17] ), .B(\CARRYB[38][17] ), .CI(\SUMB[38][18] ), 
        .CO(\CARRYB[39][17] ), .S(\SUMB[39][17] ) );
  FA1AP S2_16_29 ( .A(\ab[29][16] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA1A S2_23_27 ( .A(\ab[27][23] ), .B(\CARRYB[22][27] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA1AP S2_3_29 ( .A(\CARRYB[2][29] ), .B(n297), .CI(\SUMB[2][30] ), .CO(
        \CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA1AP S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA1P S2_25_21 ( .A(\ab[25][21] ), .B(\CARRYB[24][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA1P S2_8_27 ( .A(\CARRYB[7][27] ), .B(n446), .CI(\SUMB[7][28] ), .CO(
        \CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA1 S2_17_24 ( .A(\CARRYB[16][24] ), .B(\ab[24][17] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA1A S2_18_24 ( .A(\CARRYB[17][24] ), .B(\ab[24][18] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA1AP S2_40_29 ( .A(\ab[40][29] ), .B(\CARRYB[39][29] ), .CI(\SUMB[39][30] ), 
        .CO(\CARRYB[40][29] ), .S(\SUMB[40][29] ) );
  FA1 S2_41_29 ( .A(\ab[41][29] ), .B(\CARRYB[40][29] ), .CI(\SUMB[40][30] ), 
        .CO(\CARRYB[41][29] ), .S(\SUMB[41][29] ) );
  FA1A S2_31_32 ( .A(\ab[32][31] ), .B(\CARRYB[30][32] ), .CI(\SUMB[30][33] ), 
        .CO(\CARRYB[31][32] ), .S(\SUMB[31][32] ) );
  FA1P S2_46_27 ( .A(\ab[46][27] ), .B(\CARRYB[45][27] ), .CI(\SUMB[45][28] ), 
        .CO(\CARRYB[46][27] ), .S(\SUMB[46][27] ) );
  FA1AP S2_10_14 ( .A(n569), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), .CO(
        \CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1 S2_11_14 ( .A(n586), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), .CO(
        \CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_40_17 ( .A(\ab[40][17] ), .B(\CARRYB[39][17] ), .CI(\SUMB[39][18] ), 
        .CO(\CARRYB[40][17] ), .S(\SUMB[40][17] ) );
  FA1A S2_7_29 ( .A(n1287), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), .CO(
        \CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA1A S2_42_16 ( .A(\ab[42][16] ), .B(\CARRYB[41][16] ), .CI(\SUMB[41][17] ), 
        .CO(\CARRYB[42][16] ), .S(\SUMB[42][16] ) );
  FA1P S2_11_29 ( .A(n571), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), .CO(
        \CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA1P S2_10_10 ( .A(A[10]), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), .CO(
        \CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1 S2_2_12 ( .A(n332), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1P S2_19_8 ( .A(n484), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), .CO(
        \CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1A S2_33_4 ( .A(n353), .B(\CARRYB[32][4] ), .CI(\SUMB[32][5] ), .CO(
        \CARRYB[33][4] ), .S(\SUMB[33][4] ) );
  FA1 S2_41_28 ( .A(\ab[41][28] ), .B(\CARRYB[40][28] ), .CI(\SUMB[40][29] ), 
        .CO(\CARRYB[41][28] ), .S(\SUMB[41][28] ) );
  FA1AP S2_39_38 ( .A(\ab[39][38] ), .B(\CARRYB[38][38] ), .CI(\SUMB[38][39] ), 
        .CO(\CARRYB[39][38] ), .S(\SUMB[39][38] ) );
  FA1P S2_17_43 ( .A(\ab[43][17] ), .B(\CARRYB[16][43] ), .CI(\SUMB[16][44] ), 
        .CO(\CARRYB[17][43] ), .S(\SUMB[17][43] ) );
  FA1P S2_18_43 ( .A(\ab[43][18] ), .B(\CARRYB[17][43] ), .CI(\SUMB[17][44] ), 
        .CO(\CARRYB[18][43] ), .S(\SUMB[18][43] ) );
  FA1P S2_16_43 ( .A(\ab[43][16] ), .B(\CARRYB[15][43] ), .CI(\SUMB[15][44] ), 
        .CO(\CARRYB[16][43] ), .S(\SUMB[16][43] ) );
  FA1P S2_26_42 ( .A(\ab[42][26] ), .B(\CARRYB[25][42] ), .CI(\SUMB[25][43] ), 
        .CO(\CARRYB[26][42] ), .S(\SUMB[26][42] ) );
  FA1AP S2_27_42 ( .A(\ab[42][27] ), .B(\CARRYB[26][42] ), .CI(\SUMB[26][43] ), 
        .CO(\CARRYB[27][42] ), .S(\SUMB[27][42] ) );
  FA1P S2_46_36 ( .A(\ab[46][36] ), .B(\CARRYB[45][36] ), .CI(\SUMB[45][37] ), 
        .CO(\CARRYB[46][36] ), .S(\SUMB[46][36] ) );
  FA1P S2_13_16 ( .A(n624), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), .CO(
        \CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA1AP S2_10_18 ( .A(n557), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), .CO(
        \CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1 S2_8_17 ( .A(n500), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), .CO(
        \CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1P S2_9_17 ( .A(n515), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), .CO(
        \CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1P S2_26_11 ( .A(n578), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), .CO(
        \CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA1P S2_44_23 ( .A(\ab[44][23] ), .B(\CARRYB[43][23] ), .CI(\SUMB[43][24] ), 
        .CO(\CARRYB[44][23] ), .S(\SUMB[44][23] ) );
  FA1AP S2_43_23 ( .A(\ab[43][23] ), .B(\CARRYB[42][23] ), .CI(\SUMB[42][24] ), 
        .CO(\CARRYB[43][23] ), .S(\SUMB[43][23] ) );
  FA1P S2_45_21 ( .A(\ab[45][21] ), .B(\CARRYB[44][21] ), .CI(\SUMB[44][22] ), 
        .CO(\CARRYB[45][21] ), .S(\SUMB[45][21] ) );
  FA1AP S4_21 ( .A(\ab[47][21] ), .B(\CARRYB[46][21] ), .CI(\SUMB[46][22] ), 
        .CO(\CARRYB[47][21] ), .S(\SUMB[47][21] ) );
  FA1A S2_11_31 ( .A(n579), .B(\CARRYB[10][31] ), .CI(\SUMB[10][32] ), .CO(
        \CARRYB[11][31] ), .S(\SUMB[11][31] ) );
  FA1 S2_24_26 ( .A(\ab[26][24] ), .B(\CARRYB[23][26] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA1P S2_36_22 ( .A(\ab[36][22] ), .B(\CARRYB[35][22] ), .CI(\SUMB[35][23] ), 
        .CO(\CARRYB[36][22] ), .S(\SUMB[36][22] ) );
  FA1P S2_37_22 ( .A(\CARRYB[36][22] ), .B(\ab[37][22] ), .CI(\SUMB[36][23] ), 
        .CO(\CARRYB[37][22] ), .S(\SUMB[37][22] ) );
  FA1AP S2_7_30 ( .A(n411), .B(\CARRYB[6][30] ), .CI(\SUMB[6][31] ), .CO(
        \CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA1P S2_43_17 ( .A(\ab[43][17] ), .B(\CARRYB[42][17] ), .CI(\SUMB[42][18] ), 
        .CO(\CARRYB[43][17] ), .S(\SUMB[43][17] ) );
  FA1 S2_33_20 ( .A(\ab[33][20] ), .B(\CARRYB[32][20] ), .CI(\SUMB[32][21] ), 
        .CO(\CARRYB[33][20] ), .S(\SUMB[33][20] ) );
  FA1 S2_25_28 ( .A(\ab[28][25] ), .B(\CARRYB[24][28] ), .CI(\SUMB[24][29] ), 
        .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FA1AP S2_42_12 ( .A(\ab[42][12] ), .B(\CARRYB[41][12] ), .CI(\SUMB[41][13] ), 
        .CO(\CARRYB[42][12] ), .S(\SUMB[42][12] ) );
  FA1 S2_8_24 ( .A(n1291), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), .CO(
        \CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA1AP S2_9_24 ( .A(n513), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), .CO(
        \CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA1AP S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA1P S2_17_45 ( .A(\ab[45][17] ), .B(\CARRYB[16][45] ), .CI(\SUMB[16][46] ), 
        .CO(\CARRYB[17][45] ), .S(\SUMB[17][45] ) );
  FA1P S2_36_44 ( .A(\ab[44][36] ), .B(\CARRYB[35][44] ), .CI(\SUMB[35][45] ), 
        .CO(\CARRYB[36][44] ), .S(\SUMB[36][44] ) );
  FA1P S2_42_41 ( .A(\ab[42][41] ), .B(\CARRYB[41][41] ), .CI(\SUMB[41][42] ), 
        .CO(\CARRYB[42][41] ), .S(\SUMB[42][41] ) );
  FA1AP S2_39_43 ( .A(\ab[43][39] ), .B(\CARRYB[38][43] ), .CI(\SUMB[38][44] ), 
        .CO(\CARRYB[39][43] ), .S(\SUMB[39][43] ) );
  FA1P S2_23_45 ( .A(\ab[45][23] ), .B(\CARRYB[22][45] ), .CI(\SUMB[22][46] ), 
        .CO(\CARRYB[23][45] ), .S(\SUMB[23][45] ) );
  FA1 S2_5_14 ( .A(n414), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1AP S2_8_14 ( .A(n495), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), .CO(
        \CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1 S2_17_10 ( .A(n556), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), .CO(
        \CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA1A S2_18_9 ( .A(n528), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), .CO(
        \CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA1P S2_46_3 ( .A(n295), .B(\CARRYB[45][3] ), .CI(\SUMB[45][4] ), .CO(
        \CARRYB[46][3] ), .S(\SUMB[46][3] ) );
  FA1AP S2_29_29 ( .A(A[29]), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), .CO(
        \CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA1P S2_21_32 ( .A(\ab[32][21] ), .B(\CARRYB[20][32] ), .CI(\SUMB[20][33] ), 
        .CO(\CARRYB[21][32] ), .S(\SUMB[21][32] ) );
  FA1P S2_22_32 ( .A(\ab[32][22] ), .B(\CARRYB[21][32] ), .CI(\SUMB[21][33] ), 
        .CO(\CARRYB[22][32] ), .S(\SUMB[22][32] ) );
  FA1A S2_43_28 ( .A(\CARRYB[42][28] ), .B(\ab[43][28] ), .CI(\SUMB[42][29] ), 
        .CO(\CARRYB[43][28] ), .S(\SUMB[43][28] ) );
  FA1AP S4_13 ( .A(\ab[47][13] ), .B(\CARRYB[46][13] ), .CI(\SUMB[46][14] ), 
        .CO(\CARRYB[47][13] ), .S(\SUMB[47][13] ) );
  FA1A S2_46_25 ( .A(\ab[46][25] ), .B(\CARRYB[45][25] ), .CI(\SUMB[45][26] ), 
        .CO(\CARRYB[46][25] ), .S(\SUMB[46][25] ) );
  FA1P S2_38_30 ( .A(\CARRYB[37][30] ), .B(\ab[38][30] ), .CI(\SUMB[37][31] ), 
        .CO(\CARRYB[38][30] ), .S(\SUMB[38][30] ) );
  FA1 S2_26_34 ( .A(\ab[34][26] ), .B(\CARRYB[25][34] ), .CI(\SUMB[25][35] ), 
        .CO(\CARRYB[26][34] ), .S(\SUMB[26][34] ) );
  FA1P S2_12_32 ( .A(n601), .B(\CARRYB[11][32] ), .CI(\SUMB[11][33] ), .CO(
        \CARRYB[12][32] ), .S(\SUMB[12][32] ) );
  FA1 S2_21_29 ( .A(\ab[29][21] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA1AP S2_45_18 ( .A(\ab[45][18] ), .B(\CARRYB[44][18] ), .CI(\SUMB[44][19] ), 
        .CO(\CARRYB[45][18] ), .S(\SUMB[45][18] ) );
  FA1AP S2_23_36 ( .A(\ab[36][23] ), .B(\CARRYB[22][36] ), .CI(\SUMB[22][37] ), 
        .CO(\CARRYB[23][36] ), .S(\SUMB[23][36] ) );
  FA1 S2_23_35 ( .A(\ab[35][23] ), .B(\CARRYB[22][35] ), .CI(\SUMB[22][36] ), 
        .CO(\CARRYB[23][35] ), .S(\SUMB[23][35] ) );
  FA1AP S2_39_29 ( .A(\ab[39][29] ), .B(\CARRYB[38][29] ), .CI(\SUMB[38][30] ), 
        .CO(\CARRYB[39][29] ), .S(\SUMB[39][29] ) );
  FA1P S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA1P S2_42_8 ( .A(n534), .B(\CARRYB[41][8] ), .CI(\SUMB[41][9] ), .CO(
        \CARRYB[42][8] ), .S(\SUMB[42][8] ) );
  FA1 S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA1P S2_7_18 ( .A(n474), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), .CO(
        \CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1AP S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA1AP S2_18_20 ( .A(\ab[20][18] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA1P S2_4_41 ( .A(n320), .B(\CARRYB[3][41] ), .CI(\SUMB[3][42] ), .CO(
        \CARRYB[4][41] ), .S(\SUMB[4][41] ) );
  FA1AP S2_13_38 ( .A(\ab[38][13] ), .B(\CARRYB[12][38] ), .CI(\SUMB[12][39] ), 
        .CO(\CARRYB[13][38] ), .S(\SUMB[13][38] ) );
  FA1P S2_42_24 ( .A(\ab[42][24] ), .B(\CARRYB[41][24] ), .CI(\SUMB[41][25] ), 
        .CO(\CARRYB[42][24] ), .S(\SUMB[42][24] ) );
  FA1 S2_4_19 ( .A(n1277), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), .CO(
        \CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA1AP S2_5_19 ( .A(n1283), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), .CO(
        \CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1P S2_21_12 ( .A(n596), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), .CO(
        \CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA1P S2_15_14 ( .A(n641), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), .CO(
        \CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA1P S2_16_14 ( .A(n638), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), .CO(
        \CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA1A S2_19_12 ( .A(n605), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), .CO(
        \CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA1P S2_20_12 ( .A(n597), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), .CO(
        \CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA1A S2_32_10 ( .A(\CARRYB[31][10] ), .B(n551), .CI(\SUMB[31][11] ), .CO(
        \CARRYB[32][10] ), .S(\SUMB[32][10] ) );
  FA1A S2_42_6 ( .A(n455), .B(\CARRYB[41][6] ), .CI(\SUMB[41][7] ), .CO(
        \CARRYB[42][6] ), .S(\SUMB[42][6] ) );
  FA1A S2_30_1 ( .A(n1405), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), .CO(
        \CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA1AP S2_28_12 ( .A(\CARRYB[27][12] ), .B(n592), .CI(\SUMB[27][13] ), .CO(
        \CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA1AP S2_36_8 ( .A(n517), .B(\CARRYB[35][8] ), .CI(\SUMB[35][9] ), .CO(
        \CARRYB[36][8] ), .S(\SUMB[36][8] ) );
  FA1P S2_40_34 ( .A(\ab[40][34] ), .B(\CARRYB[39][34] ), .CI(\SUMB[39][35] ), 
        .CO(\CARRYB[40][34] ), .S(\SUMB[40][34] ) );
  FA1P S2_42_34 ( .A(\ab[42][34] ), .B(\CARRYB[41][34] ), .CI(\SUMB[41][35] ), 
        .CO(\CARRYB[42][34] ), .S(\SUMB[42][34] ) );
  FA1A S2_13_39 ( .A(\ab[39][13] ), .B(\CARRYB[12][39] ), .CI(\SUMB[12][40] ), 
        .CO(\CARRYB[13][39] ), .S(\SUMB[13][39] ) );
  FA1P S2_43_7 ( .A(n279), .B(\CARRYB[42][7] ), .CI(\SUMB[42][8] ), .CO(
        \CARRYB[43][7] ), .S(\SUMB[43][7] ) );
  FA1A S2_28_13 ( .A(n627), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), .CO(
        \CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA1 S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA1P S2_17_29 ( .A(\CARRYB[16][29] ), .B(\ab[29][17] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA1 S2_43_19 ( .A(\ab[43][19] ), .B(\CARRYB[42][19] ), .CI(\SUMB[42][20] ), 
        .CO(\CARRYB[43][19] ), .S(\SUMB[43][19] ) );
  FA1P S2_4_33 ( .A(n353), .B(\CARRYB[3][33] ), .CI(\SUMB[3][34] ), .CO(
        \CARRYB[4][33] ), .S(\SUMB[4][33] ) );
  FA1AP S2_36_21 ( .A(\ab[36][21] ), .B(\CARRYB[35][21] ), .CI(\SUMB[35][22] ), 
        .CO(\CARRYB[36][21] ), .S(\SUMB[36][21] ) );
  FA1A S2_7_32 ( .A(n440), .B(\CARRYB[6][32] ), .CI(\SUMB[6][33] ), .CO(
        \CARRYB[7][32] ), .S(\SUMB[7][32] ) );
  FA1 S2_2_27 ( .A(n1310), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), .CO(
        \CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA1P S2_9_25 ( .A(n483), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), .CO(
        \CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA1AP S2_22_35 ( .A(\ab[35][22] ), .B(\CARRYB[21][35] ), .CI(\SUMB[21][36] ), 
        .CO(\CARRYB[22][35] ), .S(\SUMB[22][35] ) );
  FA1P S2_35_30 ( .A(\ab[35][30] ), .B(\CARRYB[34][30] ), .CI(\SUMB[34][31] ), 
        .CO(\CARRYB[35][30] ), .S(\SUMB[35][30] ) );
  FA1AP S2_44_26 ( .A(\ab[44][26] ), .B(\CARRYB[43][26] ), .CI(\SUMB[43][27] ), 
        .CO(\CARRYB[44][26] ), .S(\SUMB[44][26] ) );
  FA1P S2_37_29 ( .A(\ab[37][29] ), .B(\CARRYB[36][29] ), .CI(\SUMB[36][30] ), 
        .CO(\CARRYB[37][29] ), .S(\SUMB[37][29] ) );
  FA1 S2_27_28 ( .A(\ab[28][27] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), 
        .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FA1P S2_36_26 ( .A(\ab[36][26] ), .B(\CARRYB[35][26] ), .CI(\SUMB[35][27] ), 
        .CO(\CARRYB[36][26] ), .S(\SUMB[36][26] ) );
  FA1P S2_13_9 ( .A(n530), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), .CO(
        \CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1AP S2_37_1 ( .A(n1345), .B(\CARRYB[36][1] ), .CI(\SUMB[36][2] ), .CO(
        \CARRYB[37][1] ), .S(\SUMB[37][1] ) );
  FA1A S2_15_27 ( .A(\CARRYB[14][27] ), .B(\ab[27][15] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA1AP S2_13_28 ( .A(n627), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), .CO(
        \CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA1A S2_16_25 ( .A(\ab[25][16] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA1A S2_13_29 ( .A(\CARRYB[12][29] ), .B(n621), .CI(\SUMB[12][30] ), .CO(
        \CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA1 S2_2_36 ( .A(n293), .B(\CARRYB[1][36] ), .CI(\SUMB[1][37] ), .CO(
        \CARRYB[2][36] ), .S(\SUMB[2][36] ) );
  FA1P S2_16_30 ( .A(\ab[30][16] ), .B(\CARRYB[15][30] ), .CI(\SUMB[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA1 S2_29_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), 
        .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FA1A S2_38_20 ( .A(\ab[38][20] ), .B(\CARRYB[37][20] ), .CI(\SUMB[37][21] ), 
        .CO(\CARRYB[38][20] ), .S(\SUMB[38][20] ) );
  FA1AP S4_16 ( .A(\ab[47][16] ), .B(\CARRYB[46][16] ), .CI(\SUMB[46][17] ), 
        .CO(\CARRYB[47][16] ), .S(\SUMB[47][16] ) );
  FA1A S2_22_22 ( .A(n1474), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), .CO(
        \CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA1 S2_36_19 ( .A(\ab[36][19] ), .B(\CARRYB[35][19] ), .CI(\SUMB[35][20] ), 
        .CO(\CARRYB[36][19] ), .S(\SUMB[36][19] ) );
  FA1 S2_27_32 ( .A(\SUMB[26][33] ), .B(\CARRYB[26][32] ), .CI(\ab[32][27] ), 
        .CO(\CARRYB[27][32] ), .S(\SUMB[27][32] ) );
  FA1A S2_34_29 ( .A(\ab[34][29] ), .B(\CARRYB[33][29] ), .CI(\SUMB[33][30] ), 
        .CO(\CARRYB[34][29] ), .S(\SUMB[34][29] ) );
  FA1 S2_3_14 ( .A(n338), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), .CO(
        \CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1P S2_4_14 ( .A(n366), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), .CO(
        \CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1AP S2_14_12 ( .A(n611), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), .CO(
        \CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1P S2_15_12 ( .A(n617), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), .CO(
        \CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA1P S2_21_11 ( .A(n580), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), .CO(
        \CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA1AP S2_32_32 ( .A(A[32]), .B(\CARRYB[31][32] ), .CI(\SUMB[31][33] ), .CO(
        \CARRYB[32][32] ), .S(\SUMB[32][32] ) );
  FA1P S2_16_38 ( .A(\ab[38][16] ), .B(\CARRYB[15][38] ), .CI(\SUMB[15][39] ), 
        .CO(\CARRYB[16][38] ), .S(\SUMB[16][38] ) );
  FA1A S2_19_37 ( .A(\CARRYB[18][37] ), .B(\ab[37][19] ), .CI(\SUMB[18][38] ), 
        .CO(\CARRYB[19][37] ), .S(\SUMB[19][37] ) );
  FA1P S2_20_37 ( .A(\ab[37][20] ), .B(\CARRYB[19][37] ), .CI(\SUMB[19][38] ), 
        .CO(\CARRYB[20][37] ), .S(\SUMB[20][37] ) );
  FA1A S2_44_18 ( .A(\ab[44][18] ), .B(\CARRYB[43][18] ), .CI(\SUMB[43][19] ), 
        .CO(\CARRYB[44][18] ), .S(\SUMB[44][18] ) );
  FA1A S2_18_28 ( .A(\ab[28][18] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA1AP S2_4_37 ( .A(n1274), .B(\CARRYB[3][37] ), .CI(\SUMB[3][38] ), .CO(
        \CARRYB[4][37] ), .S(\SUMB[4][37] ) );
  FA1P S2_39_25 ( .A(\ab[39][25] ), .B(\CARRYB[38][25] ), .CI(\SUMB[38][26] ), 
        .CO(\CARRYB[39][25] ), .S(\SUMB[39][25] ) );
  FA1 S2_40_25 ( .A(\ab[40][25] ), .B(\CARRYB[39][25] ), .CI(\SUMB[39][26] ), 
        .CO(\CARRYB[40][25] ), .S(\SUMB[40][25] ) );
  FA1 S2_4_24 ( .A(n1272), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), .CO(
        \CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA1A S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA1 S2_34_14 ( .A(\ab[34][14] ), .B(\CARRYB[33][14] ), .CI(\SUMB[33][15] ), 
        .CO(\CARRYB[34][14] ), .S(\SUMB[34][14] ) );
  FA1AP S2_18_36 ( .A(\ab[36][18] ), .B(\CARRYB[17][36] ), .CI(\SUMB[17][37] ), 
        .CO(\CARRYB[18][36] ), .S(\SUMB[18][36] ) );
  FA1AP S2_42_20 ( .A(\ab[42][20] ), .B(\CARRYB[41][20] ), .CI(\SUMB[41][21] ), 
        .CO(\CARRYB[42][20] ), .S(\SUMB[42][20] ) );
  FA1P S2_10_36 ( .A(n574), .B(\CARRYB[9][36] ), .CI(\SUMB[9][37] ), .CO(
        \CARRYB[10][36] ), .S(\SUMB[10][36] ) );
  FA1P S2_9_11 ( .A(n568), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), .CO(
        \CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1AP S2_3_12 ( .A(n346), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), .CO(
        \CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_16_10 ( .A(n559), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), .CO(
        \CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1A S2_36_3 ( .A(n289), .B(\CARRYB[35][3] ), .CI(\SUMB[35][4] ), .CO(
        \CARRYB[36][3] ), .S(\SUMB[36][3] ) );
  FA1 S2_17_9 ( .A(n515), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), .CO(
        \CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1A S2_6_24 ( .A(n1282), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), .CO(
        \CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA1 S2_17_20 ( .A(\ab[20][17] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA1P S2_14_39 ( .A(\ab[39][14] ), .B(\CARRYB[13][39] ), .CI(\SUMB[13][40] ), 
        .CO(\CARRYB[14][39] ), .S(\SUMB[14][39] ) );
  FA1P S2_40_28 ( .A(\ab[40][28] ), .B(\CARRYB[39][28] ), .CI(\SUMB[39][29] ), 
        .CO(\CARRYB[40][28] ), .S(\SUMB[40][28] ) );
  FA1 S2_30_29 ( .A(\ab[30][29] ), .B(\CARRYB[29][29] ), .CI(\SUMB[29][30] ), 
        .CO(\CARRYB[30][29] ), .S(\SUMB[30][29] ) );
  FA1P S2_43_24 ( .A(\ab[43][24] ), .B(\CARRYB[42][24] ), .CI(\SUMB[42][25] ), 
        .CO(\CARRYB[43][24] ), .S(\SUMB[43][24] ) );
  FA1P S2_14_37 ( .A(\SUMB[13][38] ), .B(\CARRYB[13][37] ), .CI(\ab[37][14] ), 
        .CO(\CARRYB[14][37] ), .S(\SUMB[14][37] ) );
  FA1P S2_28_29 ( .A(\ab[29][28] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA1AP S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA1A S2_35_12 ( .A(\ab[35][12] ), .B(\CARRYB[34][12] ), .CI(\SUMB[34][13] ), 
        .CO(\CARRYB[35][12] ), .S(\SUMB[35][12] ) );
  FA1A S2_35_13 ( .A(\ab[35][13] ), .B(\CARRYB[34][13] ), .CI(\SUMB[34][14] ), 
        .CO(\CARRYB[35][13] ), .S(\SUMB[35][13] ) );
  FA1A S2_46_16 ( .A(\ab[46][16] ), .B(\CARRYB[45][16] ), .CI(\SUMB[45][17] ), 
        .CO(\CARRYB[46][16] ), .S(\SUMB[46][16] ) );
  FA1 S2_30_27 ( .A(\ab[30][27] ), .B(\CARRYB[29][27] ), .CI(\SUMB[29][28] ), 
        .CO(\CARRYB[30][27] ), .S(\SUMB[30][27] ) );
  FA1A S2_42_19 ( .A(\ab[42][19] ), .B(\CARRYB[41][19] ), .CI(\SUMB[41][20] ), 
        .CO(\CARRYB[42][19] ), .S(\SUMB[42][19] ) );
  FA1 S2_17_26 ( .A(\ab[26][17] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA1P S2_19_23 ( .A(\ab[23][19] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA1A S2_40_19 ( .A(\ab[40][19] ), .B(\CARRYB[39][19] ), .CI(\SUMB[39][20] ), 
        .CO(\CARRYB[40][19] ), .S(\SUMB[40][19] ) );
  FA1 S2_39_19 ( .A(\ab[39][19] ), .B(\CARRYB[38][19] ), .CI(\SUMB[38][20] ), 
        .CO(\CARRYB[39][19] ), .S(\SUMB[39][19] ) );
  FA1AP S2_9_10 ( .A(n552), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), .CO(
        \CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1AP S2_15_8 ( .A(n492), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1P S2_28_5 ( .A(n393), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), .CO(
        \CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA1P S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA1 S2_12_26 ( .A(n595), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), .CO(
        \CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA1A S2_37_13 ( .A(\ab[37][13] ), .B(\CARRYB[36][13] ), .CI(\SUMB[36][14] ), 
        .CO(\CARRYB[37][13] ), .S(\SUMB[37][13] ) );
  FA1 S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA1P S2_32_22 ( .A(\ab[32][22] ), .B(\CARRYB[31][22] ), .CI(\SUMB[31][23] ), 
        .CO(\CARRYB[32][22] ), .S(\SUMB[32][22] ) );
  FA1A S2_18_31 ( .A(\ab[31][18] ), .B(\CARRYB[17][31] ), .CI(\SUMB[17][32] ), 
        .CO(\CARRYB[18][31] ), .S(\SUMB[18][31] ) );
  FA1AP S2_8_32 ( .A(n278), .B(\CARRYB[7][32] ), .CI(\SUMB[7][33] ), .CO(
        \CARRYB[8][32] ), .S(\SUMB[8][32] ) );
  FA1 S2_39_20 ( .A(\ab[39][20] ), .B(\CARRYB[38][20] ), .CI(\SUMB[38][21] ), 
        .CO(\CARRYB[39][20] ), .S(\SUMB[39][20] ) );
  FA1AP S2_11_23 ( .A(n582), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), .CO(
        \CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA1P S2_8_25 ( .A(n468), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), .CO(
        \CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA1A S2_15_22 ( .A(\ab[22][15] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA1AP S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA1 S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  AN2P U2 ( .A(n726), .B(n871), .Z(\CARRYB[1][31] ) );
  EO3P U3 ( .A(\CARRYB[19][31] ), .B(\ab[31][20] ), .C(\SUMB[19][32] ), .Z(
        \SUMB[20][31] ) );
  ND2 U4 ( .A(\CARRYB[19][31] ), .B(\SUMB[19][32] ), .Z(n3) );
  ND2 U5 ( .A(\CARRYB[19][31] ), .B(\ab[31][20] ), .Z(n4) );
  ND2 U6 ( .A(\SUMB[19][32] ), .B(\ab[31][20] ), .Z(n5) );
  ND3 U7 ( .A(n3), .B(n4), .C(n5), .Z(\CARRYB[20][31] ) );
  EO U8 ( .A(\CARRYB[18][31] ), .B(\ab[31][19] ), .Z(n6) );
  EO U9 ( .A(\SUMB[18][32] ), .B(n6), .Z(\SUMB[19][31] ) );
  ND2 U10 ( .A(\SUMB[18][32] ), .B(\CARRYB[18][31] ), .Z(n7) );
  ND2 U11 ( .A(\SUMB[18][32] ), .B(\ab[31][19] ), .Z(n8) );
  ND2 U12 ( .A(\CARRYB[18][31] ), .B(\ab[31][19] ), .Z(n9) );
  ND3 U13 ( .A(n7), .B(n8), .C(n9), .Z(\CARRYB[19][31] ) );
  ND2P U14 ( .A(\SUMB[2][38] ), .B(n283), .Z(n1015) );
  EOP U15 ( .A(\SUMB[22][16] ), .B(\ab[23][15] ), .Z(n967) );
  ND2P U16 ( .A(n692), .B(n693), .Z(\SUMB[3][23] ) );
  ND3 U17 ( .A(n919), .B(n920), .C(n921), .Z(\CARRYB[27][13] ) );
  EOP U18 ( .A(\CARRYB[2][22] ), .B(n1317), .Z(n10) );
  EOP U19 ( .A(\SUMB[2][23] ), .B(n10), .Z(\SUMB[3][22] ) );
  ND2 U20 ( .A(\SUMB[2][23] ), .B(\CARRYB[2][22] ), .Z(n11) );
  ND2 U21 ( .A(\SUMB[2][23] ), .B(n1317), .Z(n12) );
  ND2 U22 ( .A(\CARRYB[2][22] ), .B(n1317), .Z(n13) );
  ND3 U23 ( .A(n11), .B(n12), .C(n13), .Z(\CARRYB[3][22] ) );
  NR2P U24 ( .A(n1514), .B(n1400), .Z(n1143) );
  B4I U25 ( .A(\ab[41][41] ), .Z(n1514) );
  B4IP U26 ( .A(\ab[1][1] ), .Z(n1400) );
  ND2P U27 ( .A(\CARRYB[5][32] ), .B(\SUMB[5][33] ), .Z(n867) );
  EO U28 ( .A(\CARRYB[16][36] ), .B(\ab[36][17] ), .Z(n14) );
  EO U29 ( .A(\SUMB[16][37] ), .B(n14), .Z(\SUMB[17][36] ) );
  ND2P U30 ( .A(\SUMB[16][37] ), .B(\CARRYB[16][36] ), .Z(n15) );
  ND2P U31 ( .A(\SUMB[16][37] ), .B(\ab[36][17] ), .Z(n16) );
  ND2 U32 ( .A(\CARRYB[16][36] ), .B(\ab[36][17] ), .Z(n17) );
  ND3P U33 ( .A(n15), .B(n16), .C(n17), .Z(\CARRYB[17][36] ) );
  EO U34 ( .A(n608), .B(\CARRYB[16][12] ), .Z(n1070) );
  ND3P U35 ( .A(n1093), .B(n1094), .C(n1095), .Z(\CARRYB[36][28] ) );
  EOP U36 ( .A(\CARRYB[11][33] ), .B(\ab[33][12] ), .Z(n18) );
  EOP U37 ( .A(\SUMB[11][34] ), .B(n18), .Z(\SUMB[12][33] ) );
  ND2P U38 ( .A(\SUMB[11][34] ), .B(\CARRYB[11][33] ), .Z(n19) );
  ND2P U39 ( .A(\SUMB[11][34] ), .B(\ab[33][12] ), .Z(n20) );
  ND2 U40 ( .A(\CARRYB[11][33] ), .B(\ab[33][12] ), .Z(n21) );
  ND3P U41 ( .A(n19), .B(n20), .C(n21), .Z(\CARRYB[12][33] ) );
  EOP U42 ( .A(\CARRYB[2][36] ), .B(n289), .Z(n22) );
  EOP U43 ( .A(\SUMB[2][37] ), .B(n22), .Z(\SUMB[3][36] ) );
  ND2 U44 ( .A(\SUMB[2][37] ), .B(\CARRYB[2][36] ), .Z(n23) );
  ND2 U45 ( .A(\SUMB[2][37] ), .B(n289), .Z(n24) );
  ND2 U46 ( .A(\CARRYB[2][36] ), .B(n289), .Z(n25) );
  ND3P U47 ( .A(n23), .B(n24), .C(n25), .Z(\CARRYB[3][36] ) );
  EO3 U48 ( .A(\ab[33][25] ), .B(\CARRYB[32][25] ), .C(\SUMB[32][26] ), .Z(
        \SUMB[33][25] ) );
  ND2 U49 ( .A(\ab[33][25] ), .B(\CARRYB[32][25] ), .Z(n26) );
  ND2 U50 ( .A(\ab[33][25] ), .B(\SUMB[32][26] ), .Z(n27) );
  ND2 U51 ( .A(\CARRYB[32][25] ), .B(\SUMB[32][26] ), .Z(n28) );
  ND3P U52 ( .A(n26), .B(n27), .C(n28), .Z(\CARRYB[33][25] ) );
  EO U53 ( .A(\ab[34][25] ), .B(\SUMB[33][26] ), .Z(n29) );
  EO U54 ( .A(n29), .B(\CARRYB[33][25] ), .Z(\SUMB[34][25] ) );
  ND2P U55 ( .A(\ab[34][25] ), .B(\SUMB[33][26] ), .Z(n30) );
  ND2 U56 ( .A(\ab[34][25] ), .B(\CARRYB[33][25] ), .Z(n31) );
  ND2P U57 ( .A(\SUMB[33][26] ), .B(\CARRYB[33][25] ), .Z(n32) );
  ND3P U58 ( .A(n30), .B(n31), .C(n32), .Z(\CARRYB[34][25] ) );
  EO U59 ( .A(\CARRYB[45][14] ), .B(\ab[46][14] ), .Z(n33) );
  EO U60 ( .A(\SUMB[45][15] ), .B(n33), .Z(\SUMB[46][14] ) );
  ND2 U61 ( .A(\SUMB[45][15] ), .B(\CARRYB[45][14] ), .Z(n34) );
  ND2 U62 ( .A(\SUMB[45][15] ), .B(\ab[46][14] ), .Z(n35) );
  ND2 U63 ( .A(\CARRYB[45][14] ), .B(\ab[46][14] ), .Z(n36) );
  ND3 U64 ( .A(n34), .B(n35), .C(n36), .Z(\CARRYB[46][14] ) );
  EOP U65 ( .A(\CARRYB[16][25] ), .B(\ab[25][17] ), .Z(n37) );
  EOP U66 ( .A(\SUMB[16][26] ), .B(n37), .Z(\SUMB[17][25] ) );
  ND2 U67 ( .A(\SUMB[16][26] ), .B(\CARRYB[16][25] ), .Z(n38) );
  ND2 U68 ( .A(\SUMB[16][26] ), .B(\ab[25][17] ), .Z(n39) );
  ND2 U69 ( .A(\CARRYB[16][25] ), .B(\ab[25][17] ), .Z(n40) );
  ND3P U70 ( .A(n38), .B(n39), .C(n40), .Z(\CARRYB[17][25] ) );
  EO3 U71 ( .A(\CARRYB[13][27] ), .B(\ab[27][14] ), .C(\SUMB[13][28] ), .Z(
        \SUMB[14][27] ) );
  ND2 U72 ( .A(\CARRYB[13][27] ), .B(\SUMB[13][28] ), .Z(n41) );
  ND2 U73 ( .A(\CARRYB[13][27] ), .B(\ab[27][14] ), .Z(n42) );
  ND2 U74 ( .A(\SUMB[13][28] ), .B(\ab[27][14] ), .Z(n43) );
  ND3 U75 ( .A(n41), .B(n42), .C(n43), .Z(\CARRYB[14][27] ) );
  EO U76 ( .A(\CARRYB[44][26] ), .B(n1131), .Z(\SUMB[45][26] ) );
  EOP U77 ( .A(\SUMB[20][15] ), .B(n717), .Z(\SUMB[21][14] ) );
  IV U78 ( .A(n1325), .Z(n1002) );
  ND2P U79 ( .A(\SUMB[21][14] ), .B(n620), .Z(n729) );
  ND2P U80 ( .A(\SUMB[21][14] ), .B(\CARRYB[21][13] ), .Z(n728) );
  ND3P U81 ( .A(n911), .B(n912), .C(n913), .Z(\CARRYB[10][38] ) );
  ND3P U82 ( .A(n777), .B(n778), .C(n779), .Z(\CARRYB[3][41] ) );
  IVA U83 ( .A(\SUMB[7][41] ), .Z(n44) );
  IVP U84 ( .A(n44), .Z(n45) );
  EOP U85 ( .A(\CARRYB[37][29] ), .B(\ab[38][29] ), .Z(n46) );
  EOP U86 ( .A(\SUMB[37][30] ), .B(n46), .Z(\SUMB[38][29] ) );
  ND2 U87 ( .A(\SUMB[37][30] ), .B(\CARRYB[37][29] ), .Z(n47) );
  ND2 U88 ( .A(\SUMB[37][30] ), .B(\ab[38][29] ), .Z(n48) );
  ND2 U89 ( .A(\CARRYB[37][29] ), .B(\ab[38][29] ), .Z(n49) );
  ND3 U90 ( .A(n47), .B(n48), .C(n49), .Z(\CARRYB[38][29] ) );
  EOP U91 ( .A(\SUMB[23][36] ), .B(\ab[35][24] ), .Z(n50) );
  EOP U92 ( .A(\CARRYB[23][35] ), .B(n50), .Z(\SUMB[24][35] ) );
  ND2 U93 ( .A(\CARRYB[23][35] ), .B(\SUMB[23][36] ), .Z(n51) );
  ND2 U94 ( .A(\CARRYB[23][35] ), .B(\ab[35][24] ), .Z(n52) );
  ND2 U95 ( .A(\SUMB[23][36] ), .B(\ab[35][24] ), .Z(n53) );
  ND3 U96 ( .A(n51), .B(n52), .C(n53), .Z(\CARRYB[24][35] ) );
  ND2P U97 ( .A(\SUMB[24][35] ), .B(\ab[34][25] ), .Z(n854) );
  EOP U98 ( .A(\SUMB[42][17] ), .B(n1077), .Z(\SUMB[43][16] ) );
  EO3P U99 ( .A(\SUMB[23][30] ), .B(\ab[29][24] ), .C(\CARRYB[23][29] ), .Z(
        \SUMB[24][29] ) );
  ND2 U100 ( .A(\SUMB[23][30] ), .B(\CARRYB[23][29] ), .Z(n54) );
  ND2 U101 ( .A(\SUMB[23][30] ), .B(\ab[29][24] ), .Z(n55) );
  ND2 U102 ( .A(\CARRYB[23][29] ), .B(\ab[29][24] ), .Z(n56) );
  ND3P U103 ( .A(n54), .B(n55), .C(n56), .Z(\CARRYB[24][29] ) );
  EO3P U104 ( .A(\CARRYB[25][28] ), .B(\ab[28][26] ), .C(\SUMB[25][29] ), .Z(
        \SUMB[26][28] ) );
  ND2 U105 ( .A(\CARRYB[25][28] ), .B(\SUMB[25][29] ), .Z(n57) );
  ND2 U106 ( .A(\CARRYB[25][28] ), .B(\ab[28][26] ), .Z(n58) );
  ND2 U107 ( .A(\SUMB[25][29] ), .B(\ab[28][26] ), .Z(n59) );
  ND3P U108 ( .A(n57), .B(n58), .C(n59), .Z(\CARRYB[26][28] ) );
  ND3 U109 ( .A(n1243), .B(n1244), .C(n1245), .Z(\CARRYB[45][3] ) );
  EO U110 ( .A(\SUMB[37][40] ), .B(\ab[39][38] ), .Z(n975) );
  EO3P U111 ( .A(\ab[40][38] ), .B(\CARRYB[39][38] ), .C(\SUMB[39][39] ), .Z(
        \SUMB[40][38] ) );
  IVP U112 ( .A(n694), .Z(n249) );
  ND2P U113 ( .A(\SUMB[11][29] ), .B(n61), .Z(n62) );
  ND2 U114 ( .A(n60), .B(n764), .Z(n63) );
  ND2P U115 ( .A(n62), .B(n63), .Z(\SUMB[12][28] ) );
  IVDA U116 ( .A(\SUMB[11][29] ), .Y(n60) );
  IVP U117 ( .A(n764), .Z(n61) );
  EOP U118 ( .A(\CARRYB[42][15] ), .B(\ab[43][15] ), .Z(n64) );
  EOP U119 ( .A(\SUMB[42][16] ), .B(n64), .Z(\SUMB[43][15] ) );
  ND2 U120 ( .A(\SUMB[42][16] ), .B(\CARRYB[42][15] ), .Z(n65) );
  ND2 U121 ( .A(\SUMB[42][16] ), .B(\ab[43][15] ), .Z(n66) );
  ND2 U122 ( .A(\CARRYB[42][15] ), .B(\ab[43][15] ), .Z(n67) );
  ND3 U123 ( .A(n65), .B(n66), .C(n67), .Z(\CARRYB[43][15] ) );
  EOP U124 ( .A(\CARRYB[42][18] ), .B(n1088), .Z(\SUMB[43][18] ) );
  EOP U125 ( .A(\SUMB[42][19] ), .B(\ab[43][18] ), .Z(n1088) );
  ND3 U126 ( .A(n878), .B(n879), .C(n880), .Z(\CARRYB[19][24] ) );
  EOP U127 ( .A(\SUMB[22][19] ), .B(n860), .Z(\SUMB[23][18] ) );
  B4IP U128 ( .A(\ab[32][32] ), .Z(n1498) );
  ND2P U129 ( .A(\CARRYB[14][34] ), .B(n69), .Z(n70) );
  ND2 U130 ( .A(n68), .B(n1164), .Z(n71) );
  ND2P U131 ( .A(n70), .B(n71), .Z(\SUMB[15][34] ) );
  IVDA U132 ( .A(\CARRYB[14][34] ), .Y(n68) );
  IVP U133 ( .A(n1164), .Z(n69) );
  EOP U134 ( .A(\SUMB[6][39] ), .B(n1288), .Z(n72) );
  EOP U135 ( .A(\CARRYB[6][38] ), .B(n72), .Z(\SUMB[7][38] ) );
  ND2 U136 ( .A(\CARRYB[6][38] ), .B(\SUMB[6][39] ), .Z(n73) );
  ND2 U137 ( .A(\CARRYB[6][38] ), .B(n1288), .Z(n74) );
  ND2 U138 ( .A(\SUMB[6][39] ), .B(n1288), .Z(n75) );
  ND3 U139 ( .A(n73), .B(n74), .C(n75), .Z(\CARRYB[7][38] ) );
  EO U140 ( .A(\CARRYB[43][22] ), .B(\ab[44][22] ), .Z(n76) );
  EO U141 ( .A(\SUMB[43][23] ), .B(n76), .Z(\SUMB[44][22] ) );
  ND2P U142 ( .A(\SUMB[43][23] ), .B(\CARRYB[43][22] ), .Z(n77) );
  ND2P U143 ( .A(\SUMB[43][23] ), .B(\ab[44][22] ), .Z(n78) );
  ND2 U144 ( .A(\CARRYB[43][22] ), .B(\ab[44][22] ), .Z(n79) );
  ND3P U145 ( .A(n77), .B(n78), .C(n79), .Z(\CARRYB[44][22] ) );
  EOP U146 ( .A(\CARRYB[2][40] ), .B(n288), .Z(n80) );
  EOP U147 ( .A(\SUMB[2][41] ), .B(n80), .Z(\SUMB[3][40] ) );
  ND2 U148 ( .A(\SUMB[2][41] ), .B(\CARRYB[2][40] ), .Z(n81) );
  ND2 U149 ( .A(\SUMB[2][41] ), .B(n288), .Z(n82) );
  ND2 U150 ( .A(\CARRYB[2][40] ), .B(n288), .Z(n83) );
  ND3 U151 ( .A(n81), .B(n82), .C(n83), .Z(\CARRYB[3][40] ) );
  B4IP U152 ( .A(\ab[19][19] ), .Z(n1471) );
  AN2P U153 ( .A(n1345), .B(n1374), .Z(\CARRYB[1][37] ) );
  ND3P U154 ( .A(n657), .B(n658), .C(n659), .Z(\CARRYB[30][30] ) );
  AN2 U155 ( .A(n268), .B(n310), .Z(\CARRYB[1][21] ) );
  ND2P U156 ( .A(n395), .B(\SUMB[5][33] ), .Z(n866) );
  EO U157 ( .A(\CARRYB[42][20] ), .B(n179), .Z(\SUMB[43][20] ) );
  AN2 U158 ( .A(n1332), .B(n1327), .Z(\CARRYB[1][46] ) );
  EO3P U159 ( .A(\CARRYB[10][16] ), .B(n589), .C(\SUMB[10][17] ), .Z(
        \SUMB[11][16] ) );
  EOP U160 ( .A(\CARRYB[47][9] ), .B(\SUMB[47][10] ), .Z(\A1[55] ) );
  EO3P U161 ( .A(\CARRYB[28][9] ), .B(n509), .C(\SUMB[28][10] ), .Z(
        \SUMB[29][9] ) );
  AN2P U162 ( .A(\CARRYB[47][33] ), .B(\SUMB[47][34] ), .Z(\A2[80] ) );
  ND3 U163 ( .A(n1125), .B(n1126), .C(n1127), .Z(\CARRYB[27][4] ) );
  ND3P U164 ( .A(n214), .B(n215), .C(n216), .Z(\CARRYB[6][41] ) );
  ND2P U165 ( .A(\CARRYB[20][7] ), .B(\SUMB[20][8] ), .Z(n98) );
  ND2P U166 ( .A(\CARRYB[20][7] ), .B(n469), .Z(n99) );
  EOP U167 ( .A(\CARRYB[13][16] ), .B(n638), .Z(n670) );
  EOP U168 ( .A(\CARRYB[3][20] ), .B(n349), .Z(n674) );
  EOP U169 ( .A(n1398), .B(n1414), .Z(\SUMB[1][20] ) );
  ND2P U170 ( .A(n186), .B(n979), .Z(n189) );
  IV U171 ( .A(\SUMB[19][36] ), .Z(n186) );
  EO3 U172 ( .A(\CARRYB[16][34] ), .B(\ab[34][17] ), .C(\SUMB[16][35] ), .Z(
        \SUMB[17][34] ) );
  ND3P U173 ( .A(n252), .B(n253), .C(n254), .Z(\CARRYB[21][44] ) );
  ND2 U174 ( .A(\SUMB[40][3] ), .B(\CARRYB[40][2] ), .Z(n1227) );
  EOP U175 ( .A(\CARRYB[36][2] ), .B(n1121), .Z(\SUMB[37][2] ) );
  ND2P U176 ( .A(\CARRYB[37][3] ), .B(n343), .Z(n1204) );
  ND2P U177 ( .A(\CARRYB[37][3] ), .B(\SUMB[37][4] ), .Z(n1203) );
  EO U178 ( .A(n653), .B(\SUMB[29][31] ), .Z(\SUMB[30][30] ) );
  EOP U179 ( .A(\CARRYB[37][3] ), .B(n1202), .Z(\SUMB[38][3] ) );
  ND2P U180 ( .A(\CARRYB[35][0] ), .B(\SUMB[35][1] ), .Z(n1212) );
  EOP U181 ( .A(n1350), .B(n1143), .Z(\SUMB[1][41] ) );
  EOP U182 ( .A(\CARRYB[47][20] ), .B(\SUMB[47][21] ), .Z(\A1[66] ) );
  ND2P U183 ( .A(n287), .B(\CARRYB[2][23] ), .Z(n1067) );
  ND2P U184 ( .A(n1360), .B(n1399), .Z(n718) );
  EOP U185 ( .A(\SUMB[45][31] ), .B(n914), .Z(\SUMB[46][30] ) );
  EOP U186 ( .A(\CARRYB[45][30] ), .B(\ab[46][30] ), .Z(n914) );
  EO U187 ( .A(n151), .B(\CARRYB[45][1] ), .Z(\SUMB[46][1] ) );
  ND3P U188 ( .A(n1255), .B(n1256), .C(n1257), .Z(\CARRYB[39][1] ) );
  EO3P U189 ( .A(\CARRYB[14][15] ), .B(n1461), .C(\SUMB[14][16] ), .Z(
        \SUMB[15][15] ) );
  EOP U190 ( .A(\CARRYB[32][29] ), .B(\ab[33][29] ), .Z(n711) );
  EOP U191 ( .A(\SUMB[35][29] ), .B(n1092), .Z(\SUMB[36][28] ) );
  EOP U192 ( .A(\CARRYB[35][28] ), .B(\ab[36][28] ), .Z(n1092) );
  EOP U193 ( .A(A[30]), .B(\CARRYB[29][30] ), .Z(n653) );
  EOP U194 ( .A(\SUMB[13][20] ), .B(n636), .Z(n1020) );
  EO3P U195 ( .A(\CARRYB[22][16] ), .B(\ab[23][16] ), .C(\SUMB[22][17] ), .Z(
        \SUMB[23][16] ) );
  EOP U196 ( .A(\CARRYB[44][3] ), .B(n1242), .Z(\SUMB[45][3] ) );
  AN2 U197 ( .A(n267), .B(n1395), .Z(\CARRYB[1][15] ) );
  ND3P U198 ( .A(n865), .B(n866), .C(n867), .Z(\CARRYB[6][32] ) );
  ND3P U199 ( .A(n739), .B(n740), .C(n741), .Z(\CARRYB[5][38] ) );
  ND2P U200 ( .A(\CARRYB[39][2] ), .B(\SUMB[39][3] ), .Z(n1223) );
  ND2P U201 ( .A(n1319), .B(\CARRYB[39][2] ), .Z(n1221) );
  ND2P U202 ( .A(\CARRYB[27][3] ), .B(\SUMB[27][4] ), .Z(n1083) );
  ND2P U203 ( .A(n286), .B(\CARRYB[27][3] ), .Z(n1081) );
  EOP U204 ( .A(\CARRYB[47][41] ), .B(\SUMB[47][42] ), .Z(\A1[87] ) );
  ND3P U205 ( .A(n117), .B(n118), .C(n119), .Z(\CARRYB[46][29] ) );
  ND3P U206 ( .A(n853), .B(n854), .C(n855), .Z(\CARRYB[25][34] ) );
  EOP U207 ( .A(\CARRYB[47][42] ), .B(\SUMB[47][43] ), .Z(\A1[88] ) );
  EOP U208 ( .A(n1311), .B(\SUMB[40][3] ), .Z(n1224) );
  ND2 U209 ( .A(n286), .B(\SUMB[27][4] ), .Z(n1082) );
  ND3P U210 ( .A(n1034), .B(n1035), .C(n1036), .Z(\CARRYB[29][9] ) );
  EOP U211 ( .A(n1351), .B(n1370), .Z(\SUMB[1][13] ) );
  AN2 U212 ( .A(n1376), .B(n1431), .Z(\CARRYB[1][14] ) );
  EOP U213 ( .A(\CARRYB[10][34] ), .B(n583), .Z(n1009) );
  B4IP U214 ( .A(n1506), .Z(n1505) );
  B4IP U215 ( .A(\ab[37][37] ), .Z(n1506) );
  ND3P U216 ( .A(n968), .B(n969), .C(n970), .Z(\CARRYB[23][15] ) );
  ND3P U217 ( .A(n1188), .B(n1189), .C(n1190), .Z(\CARRYB[11][2] ) );
  AN2P U218 ( .A(\CARRYB[47][1] ), .B(\SUMB[47][2] ), .Z(\A2[48] ) );
  B4IP U219 ( .A(n1434), .Z(n1433) );
  B4IP U220 ( .A(\ab[2][2] ), .Z(n1434) );
  ND3P U221 ( .A(n1225), .B(n1226), .C(n1227), .Z(\CARRYB[41][2] ) );
  ND3 U222 ( .A(n1118), .B(n1119), .C(n1120), .Z(\CARRYB[37][36] ) );
  EOP U223 ( .A(\CARRYB[47][34] ), .B(\SUMB[47][35] ), .Z(\A1[80] ) );
  EOP U224 ( .A(\CARRYB[47][18] ), .B(\SUMB[47][19] ), .Z(\A1[64] ) );
  EO U225 ( .A(\SUMB[25][10] ), .B(n168), .Z(\SUMB[26][9] ) );
  B4IP U226 ( .A(\ab[36][36] ), .Z(n1504) );
  ND2P U227 ( .A(\CARRYB[36][2] ), .B(n309), .Z(n1123) );
  ND2P U228 ( .A(\CARRYB[36][2] ), .B(\SUMB[36][3] ), .Z(n1122) );
  ND2P U229 ( .A(\CARRYB[13][2] ), .B(n342), .Z(n1197) );
  EOP U230 ( .A(n1390), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  ND3P U231 ( .A(n1031), .B(n1032), .C(n1033), .Z(\CARRYB[38][0] ) );
  EO3P U232 ( .A(\CARRYB[14][6] ), .B(n442), .C(\SUMB[14][7] ), .Z(
        \SUMB[15][6] ) );
  ND2 U233 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(n84) );
  ND2 U234 ( .A(\CARRYB[14][6] ), .B(n442), .Z(n85) );
  ND2 U235 ( .A(\SUMB[14][7] ), .B(n442), .Z(n86) );
  ND3P U236 ( .A(n84), .B(n85), .C(n86), .Z(\CARRYB[15][6] ) );
  EOP U237 ( .A(\CARRYB[13][7] ), .B(n1160), .Z(\SUMB[14][7] ) );
  EO3P U238 ( .A(n1144), .B(\CARRYB[40][1] ), .C(\SUMB[40][2] ), .Z(
        \SUMB[41][1] ) );
  ND2 U239 ( .A(n1144), .B(\CARRYB[40][1] ), .Z(n87) );
  ND2 U240 ( .A(n1144), .B(\SUMB[40][2] ), .Z(n88) );
  ND2 U241 ( .A(\CARRYB[40][1] ), .B(\SUMB[40][2] ), .Z(n89) );
  ND3P U242 ( .A(n87), .B(n88), .C(n89), .Z(\CARRYB[41][1] ) );
  EOP U243 ( .A(n1333), .B(\SUMB[41][2] ), .Z(n90) );
  EOP U244 ( .A(n90), .B(\CARRYB[41][1] ), .Z(\SUMB[42][1] ) );
  ND2 U245 ( .A(n1333), .B(\SUMB[41][2] ), .Z(n91) );
  ND2P U246 ( .A(n1333), .B(\CARRYB[41][1] ), .Z(n92) );
  ND2P U247 ( .A(\SUMB[41][2] ), .B(\CARRYB[41][1] ), .Z(n93) );
  ND3P U248 ( .A(n91), .B(n92), .C(n93), .Z(\CARRYB[42][1] ) );
  EO3 U249 ( .A(\CARRYB[17][44] ), .B(\ab[44][18] ), .C(\SUMB[17][45] ), .Z(
        \SUMB[18][44] ) );
  ND2 U250 ( .A(\CARRYB[17][44] ), .B(\SUMB[17][45] ), .Z(n94) );
  ND2 U251 ( .A(\CARRYB[17][44] ), .B(\ab[44][18] ), .Z(n95) );
  ND2 U252 ( .A(\SUMB[17][45] ), .B(\ab[44][18] ), .Z(n96) );
  ND3P U253 ( .A(n94), .B(n95), .C(n96), .Z(\CARRYB[18][44] ) );
  EOP U254 ( .A(\SUMB[20][8] ), .B(n469), .Z(n97) );
  EOP U255 ( .A(\CARRYB[20][7] ), .B(n97), .Z(\SUMB[21][7] ) );
  ND2P U256 ( .A(\SUMB[20][8] ), .B(n469), .Z(n100) );
  ND3P U257 ( .A(n98), .B(n99), .C(n100), .Z(\CARRYB[21][7] ) );
  EOP U258 ( .A(\CARRYB[21][7] ), .B(n1156), .Z(\SUMB[22][7] ) );
  ND2 U259 ( .A(\CARRYB[10][16] ), .B(\SUMB[10][17] ), .Z(n101) );
  ND2 U260 ( .A(\CARRYB[10][16] ), .B(n589), .Z(n102) );
  ND2 U261 ( .A(\SUMB[10][17] ), .B(n589), .Z(n103) );
  ND3P U262 ( .A(n101), .B(n102), .C(n103), .Z(\CARRYB[11][16] ) );
  EO3P U263 ( .A(\CARRYB[10][17] ), .B(n581), .C(\SUMB[10][18] ), .Z(
        \SUMB[11][17] ) );
  ND2 U264 ( .A(\CARRYB[10][17] ), .B(\SUMB[10][18] ), .Z(n104) );
  ND2 U265 ( .A(\CARRYB[10][17] ), .B(n581), .Z(n105) );
  ND2 U266 ( .A(\SUMB[10][18] ), .B(n581), .Z(n106) );
  ND3 U267 ( .A(n104), .B(n105), .C(n106), .Z(\CARRYB[11][17] ) );
  EO3 U268 ( .A(\CARRYB[25][18] ), .B(\ab[26][18] ), .C(\SUMB[25][19] ), .Z(
        \SUMB[26][18] ) );
  ND2 U269 ( .A(\CARRYB[25][18] ), .B(\SUMB[25][19] ), .Z(n107) );
  ND2 U270 ( .A(\CARRYB[25][18] ), .B(\ab[26][18] ), .Z(n108) );
  ND2 U271 ( .A(\SUMB[25][19] ), .B(\ab[26][18] ), .Z(n109) );
  ND3P U272 ( .A(n107), .B(n108), .C(n109), .Z(\CARRYB[26][18] ) );
  EO3P U273 ( .A(\ab[37][31] ), .B(\CARRYB[30][37] ), .C(\SUMB[30][38] ), .Z(
        \SUMB[31][37] ) );
  EOP U274 ( .A(\ab[36][32] ), .B(\CARRYB[31][36] ), .Z(n110) );
  EOP U275 ( .A(n110), .B(\SUMB[31][37] ), .Z(\SUMB[32][36] ) );
  ND2 U276 ( .A(\ab[37][31] ), .B(\CARRYB[30][37] ), .Z(n111) );
  ND2 U277 ( .A(\ab[37][31] ), .B(\SUMB[30][38] ), .Z(n112) );
  ND2 U278 ( .A(\CARRYB[30][37] ), .B(\SUMB[30][38] ), .Z(n113) );
  ND3 U279 ( .A(n111), .B(n112), .C(n113), .Z(\CARRYB[31][37] ) );
  ND2P U280 ( .A(\ab[36][32] ), .B(\CARRYB[31][36] ), .Z(n114) );
  ND2P U281 ( .A(\ab[36][32] ), .B(\SUMB[31][37] ), .Z(n115) );
  ND2P U282 ( .A(\CARRYB[31][36] ), .B(\SUMB[31][37] ), .Z(n116) );
  ND3P U283 ( .A(n114), .B(n115), .C(n116), .Z(\CARRYB[32][36] ) );
  EO3 U284 ( .A(\CARRYB[45][29] ), .B(\ab[46][29] ), .C(\SUMB[45][30] ), .Z(
        \SUMB[46][29] ) );
  ND2 U285 ( .A(\CARRYB[45][29] ), .B(\SUMB[45][30] ), .Z(n117) );
  ND2 U286 ( .A(\CARRYB[45][29] ), .B(\ab[46][29] ), .Z(n118) );
  ND2 U287 ( .A(\SUMB[45][30] ), .B(\ab[46][29] ), .Z(n119) );
  EO3 U288 ( .A(\CARRYB[27][35] ), .B(\ab[35][28] ), .C(\SUMB[27][36] ), .Z(
        \SUMB[28][35] ) );
  ND2 U289 ( .A(\CARRYB[27][35] ), .B(\SUMB[27][36] ), .Z(n120) );
  ND2 U290 ( .A(\CARRYB[27][35] ), .B(\ab[35][28] ), .Z(n121) );
  ND2 U291 ( .A(\SUMB[27][36] ), .B(\ab[35][28] ), .Z(n122) );
  ND3P U292 ( .A(n120), .B(n121), .C(n122), .Z(\CARRYB[28][35] ) );
  EOP U293 ( .A(\SUMB[17][36] ), .B(\ab[35][18] ), .Z(n123) );
  EOP U294 ( .A(\CARRYB[17][35] ), .B(n123), .Z(\SUMB[18][35] ) );
  ND2 U295 ( .A(\CARRYB[17][35] ), .B(\SUMB[17][36] ), .Z(n124) );
  ND2 U296 ( .A(\CARRYB[17][35] ), .B(\ab[35][18] ), .Z(n125) );
  ND2 U297 ( .A(\SUMB[17][36] ), .B(\ab[35][18] ), .Z(n126) );
  ND3P U298 ( .A(n124), .B(n125), .C(n126), .Z(\CARRYB[18][35] ) );
  EO3 U299 ( .A(\CARRYB[2][11] ), .B(n331), .C(\SUMB[2][12] ), .Z(
        \SUMB[3][11] ) );
  ND2 U300 ( .A(\CARRYB[2][11] ), .B(\SUMB[2][12] ), .Z(n127) );
  ND2 U301 ( .A(\CARRYB[2][11] ), .B(n331), .Z(n128) );
  ND2 U302 ( .A(\SUMB[2][12] ), .B(n331), .Z(n129) );
  ND3P U303 ( .A(n127), .B(n128), .C(n129), .Z(\CARRYB[3][11] ) );
  EO3 U304 ( .A(\CARRYB[19][34] ), .B(\ab[34][20] ), .C(\SUMB[19][35] ), .Z(
        \SUMB[20][34] ) );
  ND2 U305 ( .A(\CARRYB[19][34] ), .B(\SUMB[19][35] ), .Z(n130) );
  ND2 U306 ( .A(\CARRYB[19][34] ), .B(\ab[34][20] ), .Z(n131) );
  ND2 U307 ( .A(\SUMB[19][35] ), .B(\ab[34][20] ), .Z(n132) );
  ND3P U308 ( .A(n130), .B(n131), .C(n132), .Z(\CARRYB[20][34] ) );
  EO3P U309 ( .A(\CARRYB[7][11] ), .B(n533), .C(\SUMB[7][12] ), .Z(
        \SUMB[8][11] ) );
  ND2 U310 ( .A(\CARRYB[7][11] ), .B(\SUMB[7][12] ), .Z(n133) );
  ND2 U311 ( .A(\CARRYB[7][11] ), .B(n533), .Z(n134) );
  ND2 U312 ( .A(\SUMB[7][12] ), .B(n533), .Z(n135) );
  ND3 U313 ( .A(n133), .B(n134), .C(n135), .Z(\CARRYB[8][11] ) );
  EO3 U314 ( .A(\CARRYB[15][31] ), .B(\ab[31][16] ), .C(\SUMB[15][32] ), .Z(
        \SUMB[16][31] ) );
  ND2 U315 ( .A(\CARRYB[15][31] ), .B(\SUMB[15][32] ), .Z(n136) );
  ND2 U316 ( .A(\CARRYB[15][31] ), .B(\ab[31][16] ), .Z(n137) );
  ND2 U317 ( .A(\SUMB[15][32] ), .B(\ab[31][16] ), .Z(n138) );
  ND3P U318 ( .A(n136), .B(n137), .C(n138), .Z(\CARRYB[16][31] ) );
  EO3 U319 ( .A(\CARRYB[30][4] ), .B(n365), .C(\SUMB[30][5] ), .Z(
        \SUMB[31][4] ) );
  ND2 U320 ( .A(\CARRYB[30][4] ), .B(\SUMB[30][5] ), .Z(n139) );
  ND2 U321 ( .A(\CARRYB[30][4] ), .B(n365), .Z(n140) );
  ND2 U322 ( .A(\SUMB[30][5] ), .B(n365), .Z(n141) );
  ND3P U323 ( .A(n139), .B(n140), .C(n141), .Z(\CARRYB[31][4] ) );
  EO3P U324 ( .A(\CARRYB[16][14] ), .B(n643), .C(\SUMB[16][15] ), .Z(
        \SUMB[17][14] ) );
  ND2P U325 ( .A(\CARRYB[16][14] ), .B(\SUMB[16][15] ), .Z(n142) );
  ND2P U326 ( .A(\CARRYB[16][14] ), .B(n643), .Z(n143) );
  ND2 U327 ( .A(\SUMB[16][15] ), .B(n643), .Z(n144) );
  ND3P U328 ( .A(n142), .B(n143), .C(n144), .Z(\CARRYB[17][14] ) );
  EO3 U329 ( .A(\CARRYB[5][33] ), .B(n434), .C(\SUMB[5][34] ), .Z(
        \SUMB[6][33] ) );
  ND2 U330 ( .A(\CARRYB[5][33] ), .B(\SUMB[5][34] ), .Z(n145) );
  ND2 U331 ( .A(\CARRYB[5][33] ), .B(n434), .Z(n146) );
  ND2 U332 ( .A(\SUMB[5][34] ), .B(n434), .Z(n147) );
  ND3P U333 ( .A(n145), .B(n146), .C(n147), .Z(\CARRYB[6][33] ) );
  ND2P U334 ( .A(\CARRYB[6][33] ), .B(n445), .Z(n264) );
  EO3P U335 ( .A(n304), .B(\CARRYB[44][1] ), .C(\SUMB[44][2] ), .Z(
        \SUMB[45][1] ) );
  ND2 U336 ( .A(n304), .B(\CARRYB[44][1] ), .Z(n148) );
  ND2 U337 ( .A(n304), .B(\SUMB[44][2] ), .Z(n149) );
  ND2 U338 ( .A(\CARRYB[44][1] ), .B(\SUMB[44][2] ), .Z(n150) );
  ND3P U339 ( .A(n148), .B(n149), .C(n150), .Z(\CARRYB[45][1] ) );
  EOP U340 ( .A(n1332), .B(\SUMB[45][2] ), .Z(n151) );
  ND2 U341 ( .A(n1332), .B(\SUMB[45][2] ), .Z(n152) );
  ND2 U342 ( .A(n1332), .B(\CARRYB[45][1] ), .Z(n153) );
  ND2 U343 ( .A(\SUMB[45][2] ), .B(\CARRYB[45][1] ), .Z(n154) );
  ND3P U344 ( .A(n152), .B(n153), .C(n154), .Z(\CARRYB[46][1] ) );
  EOP U345 ( .A(\SUMB[24][7] ), .B(n405), .Z(n155) );
  EOP U346 ( .A(\CARRYB[24][6] ), .B(n155), .Z(\SUMB[25][6] ) );
  ND2P U347 ( .A(\CARRYB[24][6] ), .B(\SUMB[24][7] ), .Z(n156) );
  ND2P U348 ( .A(\CARRYB[24][6] ), .B(n405), .Z(n157) );
  ND2 U349 ( .A(\SUMB[24][7] ), .B(n405), .Z(n158) );
  ND3P U350 ( .A(n156), .B(n157), .C(n158), .Z(\CARRYB[25][6] ) );
  EO U351 ( .A(\CARRYB[29][6] ), .B(n373), .Z(n159) );
  EO U352 ( .A(\SUMB[29][7] ), .B(n159), .Z(\SUMB[30][6] ) );
  EO3 U353 ( .A(\CARRYB[3][43] ), .B(n337), .C(\SUMB[3][44] ), .Z(
        \SUMB[4][43] ) );
  ND2 U354 ( .A(\CARRYB[3][43] ), .B(\SUMB[3][44] ), .Z(n160) );
  ND2 U355 ( .A(\CARRYB[3][43] ), .B(n337), .Z(n161) );
  ND2 U356 ( .A(\SUMB[3][44] ), .B(n337), .Z(n162) );
  ND3P U357 ( .A(n160), .B(n161), .C(n162), .Z(\CARRYB[4][43] ) );
  EOP U358 ( .A(\SUMB[7][41] ), .B(n454), .Z(n163) );
  EOP U359 ( .A(\CARRYB[7][40] ), .B(n163), .Z(\SUMB[8][40] ) );
  ND2 U360 ( .A(n529), .B(\SUMB[8][40] ), .Z(n208) );
  ND2 U361 ( .A(\CARRYB[8][39] ), .B(\SUMB[8][40] ), .Z(n209) );
  EO U362 ( .A(\SUMB[12][12] ), .B(n587), .Z(n164) );
  EO U363 ( .A(\CARRYB[12][11] ), .B(n164), .Z(\SUMB[13][11] ) );
  ND2 U364 ( .A(\CARRYB[12][11] ), .B(\SUMB[12][12] ), .Z(n165) );
  ND2 U365 ( .A(\CARRYB[12][11] ), .B(n587), .Z(n166) );
  ND2 U366 ( .A(\SUMB[12][12] ), .B(n587), .Z(n167) );
  ND3 U367 ( .A(n165), .B(n166), .C(n167), .Z(\CARRYB[13][11] ) );
  EOP U368 ( .A(\CARRYB[25][9] ), .B(n523), .Z(n168) );
  ND2P U369 ( .A(\SUMB[25][10] ), .B(\CARRYB[25][9] ), .Z(n169) );
  ND2P U370 ( .A(\SUMB[25][10] ), .B(n523), .Z(n170) );
  ND2 U371 ( .A(\CARRYB[25][9] ), .B(n523), .Z(n171) );
  ND3P U372 ( .A(n169), .B(n170), .C(n171), .Z(\CARRYB[26][9] ) );
  EO3 U373 ( .A(\ab[43][22] ), .B(\CARRYB[21][43] ), .C(\SUMB[21][44] ), .Z(
        \SUMB[22][43] ) );
  ND2P U374 ( .A(\ab[43][22] ), .B(\CARRYB[21][43] ), .Z(n172) );
  ND2 U375 ( .A(\ab[43][22] ), .B(\SUMB[21][44] ), .Z(n173) );
  ND2P U376 ( .A(\CARRYB[21][43] ), .B(\SUMB[21][44] ), .Z(n174) );
  ND3P U377 ( .A(n172), .B(n173), .C(n174), .Z(\CARRYB[22][43] ) );
  EO U378 ( .A(\ab[43][23] ), .B(\SUMB[22][44] ), .Z(n175) );
  EOP U379 ( .A(n175), .B(\CARRYB[22][43] ), .Z(\SUMB[23][43] ) );
  ND2 U380 ( .A(\ab[43][23] ), .B(\SUMB[22][44] ), .Z(n176) );
  ND2P U381 ( .A(\ab[43][23] ), .B(\CARRYB[22][43] ), .Z(n177) );
  ND2P U382 ( .A(\SUMB[22][44] ), .B(\CARRYB[22][43] ), .Z(n178) );
  ND3P U383 ( .A(n176), .B(n177), .C(n178), .Z(\CARRYB[23][43] ) );
  EOP U384 ( .A(\SUMB[42][21] ), .B(\ab[43][20] ), .Z(n179) );
  ND2P U385 ( .A(\CARRYB[42][20] ), .B(\SUMB[42][21] ), .Z(n180) );
  ND2P U386 ( .A(\CARRYB[42][20] ), .B(\ab[43][20] ), .Z(n181) );
  ND2 U387 ( .A(\SUMB[42][21] ), .B(\ab[43][20] ), .Z(n182) );
  ND3P U388 ( .A(n180), .B(n181), .C(n182), .Z(\CARRYB[43][20] ) );
  EO3P U389 ( .A(\CARRYB[4][21] ), .B(n400), .C(\SUMB[4][22] ), .Z(
        \SUMB[5][21] ) );
  ND2P U390 ( .A(\CARRYB[4][21] ), .B(\SUMB[4][22] ), .Z(n183) );
  ND2P U391 ( .A(\CARRYB[4][21] ), .B(n400), .Z(n184) );
  ND2 U392 ( .A(\SUMB[4][22] ), .B(n400), .Z(n185) );
  ND3P U393 ( .A(n183), .B(n184), .C(n185), .Z(\CARRYB[5][21] ) );
  ND2P U394 ( .A(\SUMB[19][36] ), .B(n187), .Z(n188) );
  ND2P U395 ( .A(n188), .B(n189), .Z(\SUMB[20][35] ) );
  IVAP U396 ( .A(n979), .Z(n187) );
  EOP U397 ( .A(\CARRYB[19][35] ), .B(\ab[35][20] ), .Z(n979) );
  EO3 U398 ( .A(\CARRYB[20][34] ), .B(\ab[34][21] ), .C(\SUMB[20][35] ), .Z(
        \SUMB[21][34] ) );
  EO U399 ( .A(\ab[46][17] ), .B(\ab[47][16] ), .Z(n190) );
  EOP U400 ( .A(\CARRYB[16][46] ), .B(n190), .Z(\SUMB[17][46] ) );
  ND2P U401 ( .A(\CARRYB[16][46] ), .B(\ab[46][17] ), .Z(n191) );
  ND2P U402 ( .A(\CARRYB[16][46] ), .B(\ab[47][16] ), .Z(n192) );
  ND2 U403 ( .A(\ab[46][17] ), .B(\ab[47][16] ), .Z(n193) );
  ND3P U404 ( .A(n191), .B(n192), .C(n193), .Z(\CARRYB[17][46] ) );
  EO3P U405 ( .A(\CARRYB[43][1] ), .B(n1357), .C(\SUMB[43][2] ), .Z(
        \SUMB[44][1] ) );
  ND2 U406 ( .A(\CARRYB[43][1] ), .B(\SUMB[43][2] ), .Z(n194) );
  ND2 U407 ( .A(\CARRYB[43][1] ), .B(n1357), .Z(n195) );
  ND2 U408 ( .A(\SUMB[43][2] ), .B(n1357), .Z(n196) );
  ND3 U409 ( .A(n194), .B(n195), .C(n196), .Z(\CARRYB[44][1] ) );
  ND3P U410 ( .A(n1267), .B(n1268), .C(n1269), .Z(\CARRYB[43][1] ) );
  EO3P U411 ( .A(\CARRYB[24][10] ), .B(n540), .C(\SUMB[24][11] ), .Z(
        \SUMB[25][10] ) );
  ND2 U412 ( .A(\CARRYB[24][10] ), .B(\SUMB[24][11] ), .Z(n197) );
  ND2 U413 ( .A(\CARRYB[24][10] ), .B(n540), .Z(n198) );
  ND2 U414 ( .A(\SUMB[24][11] ), .B(n540), .Z(n199) );
  ND3P U415 ( .A(n197), .B(n198), .C(n199), .Z(\CARRYB[25][10] ) );
  ND2 U416 ( .A(\CARRYB[14][15] ), .B(\SUMB[14][16] ), .Z(n200) );
  ND2 U417 ( .A(\CARRYB[14][15] ), .B(n1461), .Z(n201) );
  ND2 U418 ( .A(\SUMB[14][16] ), .B(n1461), .Z(n202) );
  ND3P U419 ( .A(n200), .B(n201), .C(n202), .Z(\CARRYB[15][15] ) );
  IVA U420 ( .A(n1463), .Z(n1461) );
  EOP U421 ( .A(\SUMB[13][17] ), .B(n670), .Z(\SUMB[14][16] ) );
  EOP U422 ( .A(n529), .B(\CARRYB[8][39] ), .Z(n203) );
  EOP U423 ( .A(n203), .B(\SUMB[8][40] ), .Z(\SUMB[9][39] ) );
  ND2 U424 ( .A(n454), .B(\CARRYB[7][40] ), .Z(n204) );
  ND2 U425 ( .A(n454), .B(n45), .Z(n205) );
  ND2 U426 ( .A(\CARRYB[7][40] ), .B(n45), .Z(n206) );
  ND3P U427 ( .A(n204), .B(n205), .C(n206), .Z(\CARRYB[8][40] ) );
  ND2 U428 ( .A(n529), .B(\CARRYB[8][39] ), .Z(n207) );
  ND3 U429 ( .A(n207), .B(n208), .C(n209), .Z(\CARRYB[9][39] ) );
  EOP U430 ( .A(\SUMB[15][23] ), .B(\ab[22][16] ), .Z(n210) );
  EOP U431 ( .A(\CARRYB[15][22] ), .B(n210), .Z(\SUMB[16][22] ) );
  ND2P U432 ( .A(\CARRYB[15][22] ), .B(\SUMB[15][23] ), .Z(n211) );
  ND2P U433 ( .A(\CARRYB[15][22] ), .B(\ab[22][16] ), .Z(n212) );
  ND2 U434 ( .A(\SUMB[15][23] ), .B(\ab[22][16] ), .Z(n213) );
  ND3P U435 ( .A(n211), .B(n212), .C(n213), .Z(\CARRYB[16][22] ) );
  EO3P U436 ( .A(\CARRYB[5][41] ), .B(n443), .C(\SUMB[5][42] ), .Z(
        \SUMB[6][41] ) );
  ND2 U437 ( .A(\CARRYB[5][41] ), .B(\SUMB[5][42] ), .Z(n214) );
  ND2 U438 ( .A(\CARRYB[5][41] ), .B(n443), .Z(n215) );
  ND2 U439 ( .A(\SUMB[5][42] ), .B(n443), .Z(n216) );
  EO3 U440 ( .A(\CARRYB[38][21] ), .B(\ab[39][21] ), .C(\SUMB[38][22] ), .Z(
        \SUMB[39][21] ) );
  ND2 U441 ( .A(\CARRYB[38][21] ), .B(\SUMB[38][22] ), .Z(n217) );
  ND2 U442 ( .A(\CARRYB[38][21] ), .B(\ab[39][21] ), .Z(n218) );
  ND2 U443 ( .A(\SUMB[38][22] ), .B(\ab[39][21] ), .Z(n219) );
  ND3P U444 ( .A(n217), .B(n218), .C(n219), .Z(\CARRYB[39][21] ) );
  EOP U445 ( .A(\SUMB[19][42] ), .B(\ab[41][20] ), .Z(n220) );
  EOP U446 ( .A(\CARRYB[19][41] ), .B(n220), .Z(\SUMB[20][41] ) );
  ND2P U447 ( .A(\CARRYB[19][41] ), .B(\SUMB[19][42] ), .Z(n221) );
  ND2P U448 ( .A(\CARRYB[19][41] ), .B(\ab[41][20] ), .Z(n222) );
  ND2 U449 ( .A(\SUMB[19][42] ), .B(\ab[41][20] ), .Z(n223) );
  ND3P U450 ( .A(n221), .B(n222), .C(n223), .Z(\CARRYB[20][41] ) );
  EO3 U451 ( .A(\CARRYB[7][9] ), .B(n526), .C(\SUMB[7][10] ), .Z(\SUMB[8][9] )
         );
  ND2 U452 ( .A(\CARRYB[7][9] ), .B(\SUMB[7][10] ), .Z(n224) );
  ND2 U453 ( .A(\CARRYB[7][9] ), .B(n526), .Z(n225) );
  ND2 U454 ( .A(\SUMB[7][10] ), .B(n526), .Z(n226) );
  ND3P U455 ( .A(n224), .B(n225), .C(n226), .Z(\CARRYB[8][9] ) );
  EOP U456 ( .A(\SUMB[6][22] ), .B(n469), .Z(n227) );
  EOP U457 ( .A(\CARRYB[6][21] ), .B(n227), .Z(\SUMB[7][21] ) );
  ND2P U458 ( .A(\CARRYB[6][21] ), .B(\SUMB[6][22] ), .Z(n228) );
  ND2P U459 ( .A(\CARRYB[6][21] ), .B(n469), .Z(n229) );
  ND2 U460 ( .A(\SUMB[6][22] ), .B(n469), .Z(n230) );
  ND3P U461 ( .A(n228), .B(n229), .C(n230), .Z(\CARRYB[7][21] ) );
  EO3 U462 ( .A(\CARRYB[18][45] ), .B(\ab[45][19] ), .C(\SUMB[18][46] ), .Z(
        \SUMB[19][45] ) );
  ND2 U463 ( .A(\CARRYB[18][45] ), .B(\SUMB[18][46] ), .Z(n231) );
  ND2 U464 ( .A(\CARRYB[18][45] ), .B(\ab[45][19] ), .Z(n232) );
  ND2 U465 ( .A(\SUMB[18][46] ), .B(\ab[45][19] ), .Z(n233) );
  ND3 U466 ( .A(n231), .B(n232), .C(n233), .Z(\CARRYB[19][45] ) );
  EO U467 ( .A(\SUMB[29][43] ), .B(\ab[42][30] ), .Z(n234) );
  EO U468 ( .A(\CARRYB[29][42] ), .B(n234), .Z(\SUMB[30][42] ) );
  ND2P U469 ( .A(\CARRYB[29][42] ), .B(\SUMB[29][43] ), .Z(n235) );
  ND2P U470 ( .A(\CARRYB[29][42] ), .B(\ab[42][30] ), .Z(n236) );
  ND2 U471 ( .A(\SUMB[29][43] ), .B(\ab[42][30] ), .Z(n237) );
  ND3P U472 ( .A(n235), .B(n236), .C(n237), .Z(\CARRYB[30][42] ) );
  EO3 U473 ( .A(\CARRYB[6][42] ), .B(n498), .C(\SUMB[6][43] ), .Z(
        \SUMB[7][42] ) );
  ND2 U474 ( .A(\CARRYB[6][42] ), .B(\SUMB[6][43] ), .Z(n238) );
  ND2 U475 ( .A(\CARRYB[6][42] ), .B(n498), .Z(n239) );
  ND2 U476 ( .A(\SUMB[6][43] ), .B(n498), .Z(n240) );
  ND3P U477 ( .A(n238), .B(n239), .C(n240), .Z(\CARRYB[7][42] ) );
  ND2 U478 ( .A(\CARRYB[12][40] ), .B(n242), .Z(n243) );
  ND2 U479 ( .A(n241), .B(n1037), .Z(n244) );
  ND2 U480 ( .A(n243), .B(n244), .Z(\SUMB[13][40] ) );
  IVDA U481 ( .A(\CARRYB[12][40] ), .Y(n241) );
  IV U482 ( .A(n1037), .Z(n242) );
  EOP U483 ( .A(\SUMB[12][41] ), .B(\ab[40][13] ), .Z(n1037) );
  EO3P U484 ( .A(\CARRYB[9][8] ), .B(n508), .C(\SUMB[9][9] ), .Z(\SUMB[10][8] ) );
  ND2 U485 ( .A(\CARRYB[9][8] ), .B(\SUMB[9][9] ), .Z(n245) );
  ND2 U486 ( .A(\CARRYB[9][8] ), .B(n508), .Z(n246) );
  ND2 U487 ( .A(\SUMB[9][9] ), .B(n508), .Z(n247) );
  ND3P U488 ( .A(n245), .B(n246), .C(n247), .Z(\CARRYB[10][8] ) );
  ND2P U489 ( .A(\CARRYB[29][32] ), .B(n249), .Z(n250) );
  ND2 U490 ( .A(n248), .B(n694), .Z(n251) );
  ND2P U491 ( .A(n250), .B(n251), .Z(\SUMB[30][32] ) );
  IVDA U492 ( .A(\CARRYB[29][32] ), .Y(n248) );
  EOP U493 ( .A(\SUMB[29][33] ), .B(\ab[32][30] ), .Z(n694) );
  EO3P U494 ( .A(\CARRYB[20][44] ), .B(\ab[44][21] ), .C(\SUMB[20][45] ), .Z(
        \SUMB[21][44] ) );
  ND2 U495 ( .A(\CARRYB[20][44] ), .B(\SUMB[20][45] ), .Z(n252) );
  ND2 U496 ( .A(\CARRYB[20][44] ), .B(\ab[44][21] ), .Z(n253) );
  ND2 U497 ( .A(\SUMB[20][45] ), .B(\ab[44][21] ), .Z(n254) );
  ND2P U498 ( .A(\CARRYB[47][7] ), .B(n256), .Z(n257) );
  ND2 U499 ( .A(n255), .B(\SUMB[47][8] ), .Z(n258) );
  ND2P U500 ( .A(n257), .B(n258), .Z(\A1[53] ) );
  IVDA U501 ( .A(\CARRYB[47][7] ), .Y(n255) );
  IVP U502 ( .A(\SUMB[47][8] ), .Z(n256) );
  EOP U503 ( .A(\SUMB[39][43] ), .B(\ab[42][40] ), .Z(n259) );
  EOP U504 ( .A(\CARRYB[39][42] ), .B(n259), .Z(\SUMB[40][42] ) );
  ND2 U505 ( .A(\CARRYB[39][42] ), .B(\SUMB[39][43] ), .Z(n260) );
  ND2 U506 ( .A(\CARRYB[39][42] ), .B(\ab[42][40] ), .Z(n261) );
  ND2 U507 ( .A(\SUMB[39][43] ), .B(\ab[42][40] ), .Z(n262) );
  ND3 U508 ( .A(n260), .B(n261), .C(n262), .Z(\CARRYB[40][42] ) );
  EO3P U509 ( .A(\CARRYB[6][33] ), .B(n445), .C(\SUMB[6][34] ), .Z(
        \SUMB[7][33] ) );
  ND2 U510 ( .A(\CARRYB[6][33] ), .B(\SUMB[6][34] ), .Z(n263) );
  ND2 U511 ( .A(\SUMB[6][34] ), .B(n445), .Z(n265) );
  ND3P U512 ( .A(n263), .B(n264), .C(n265), .Z(\CARRYB[7][33] ) );
  ND3P U513 ( .A(n1053), .B(n1054), .C(n1055), .Z(\CARRYB[31][1] ) );
  ND3P U514 ( .A(n956), .B(n957), .C(n958), .Z(\CARRYB[37][21] ) );
  EOP U515 ( .A(n1224), .B(\CARRYB[40][2] ), .Z(\SUMB[41][2] ) );
  EOP U516 ( .A(\SUMB[30][13] ), .B(n873), .Z(\SUMB[31][12] ) );
  EOP U517 ( .A(n1349), .B(n1372), .Z(\SUMB[1][33] ) );
  ND2P U518 ( .A(\ab[1][1] ), .B(n1349), .Z(n725) );
  AN2P U519 ( .A(\ab[34][34] ), .B(\B[0] ), .Z(n1349) );
  ND2P U520 ( .A(n716), .B(\CARRYB[35][0] ), .Z(n1210) );
  AN2 U521 ( .A(n1357), .B(n1415), .Z(\CARRYB[1][44] ) );
  EOP U522 ( .A(n1415), .B(n1357), .Z(\SUMB[1][44] ) );
  EOP U523 ( .A(\CARRYB[47][28] ), .B(\SUMB[47][29] ), .Z(\A1[74] ) );
  EOP U524 ( .A(\SUMB[42][2] ), .B(n1422), .Z(n1266) );
  ND3P U525 ( .A(n996), .B(n997), .C(n998), .Z(\CARRYB[35][8] ) );
  ND3P U526 ( .A(n925), .B(n926), .C(n927), .Z(\CARRYB[33][10] ) );
  B4IP U527 ( .A(\ab[3][3] ), .Z(n1439) );
  ND2P U528 ( .A(\CARRYB[17][6] ), .B(n428), .Z(n1141) );
  NR2P U529 ( .A(n1457), .B(n872), .Z(n1386) );
  B4I U530 ( .A(\ab[8][8] ), .Z(n1457) );
  ND3P U531 ( .A(n922), .B(n923), .C(n924), .Z(\CARRYB[30][6] ) );
  ND3P U532 ( .A(n985), .B(n986), .C(n987), .Z(\CARRYB[29][7] ) );
  ND3P U533 ( .A(n1136), .B(n1137), .C(n1138), .Z(\CARRYB[35][4] ) );
  EOP U534 ( .A(n1327), .B(n1332), .Z(\SUMB[1][46] ) );
  ND2 U535 ( .A(n1364), .B(\SUMB[36][1] ), .Z(n1214) );
  ND2 U536 ( .A(n1364), .B(\CARRYB[36][0] ), .Z(n1215) );
  ND2 U537 ( .A(\SUMB[1][41] ), .B(\CARRYB[1][40] ), .Z(n780) );
  ND2 U538 ( .A(\CARRYB[14][30] ), .B(\ab[30][15] ), .Z(n901) );
  ND2 U539 ( .A(\CARRYB[14][30] ), .B(\SUMB[14][31] ), .Z(n900) );
  ND2 U540 ( .A(\CARRYB[14][36] ), .B(\ab[36][15] ), .Z(n828) );
  ND2 U541 ( .A(\CARRYB[17][38] ), .B(\ab[38][18] ), .Z(n789) );
  ND3 U542 ( .A(n1165), .B(n1166), .C(n1167), .Z(\CARRYB[15][34] ) );
  ND3 U543 ( .A(n931), .B(n932), .C(n933), .Z(\CARRYB[21][34] ) );
  ND3 U544 ( .A(n731), .B(n732), .C(n733), .Z(\CARRYB[21][14] ) );
  ND2 U545 ( .A(\SUMB[30][13] ), .B(\CARRYB[30][12] ), .Z(n874) );
  ND2 U546 ( .A(\CARRYB[36][36] ), .B(\SUMB[36][37] ), .Z(n1118) );
  ND2 U547 ( .A(\CARRYB[35][7] ), .B(\SUMB[35][8] ), .Z(n1001) );
  ND3 U548 ( .A(n1239), .B(n1240), .C(n1241), .Z(\CARRYB[4][4] ) );
  ND2 U549 ( .A(n1440), .B(\SUMB[3][5] ), .Z(n1239) );
  ND3 U550 ( .A(n1228), .B(n1229), .C(n1230), .Z(\CARRYB[34][3] ) );
  ND3 U551 ( .A(n1263), .B(n1264), .C(n1265), .Z(\CARRYB[35][1] ) );
  ND3 U552 ( .A(n796), .B(n797), .C(n798), .Z(\CARRYB[3][45] ) );
  ND2 U553 ( .A(\SUMB[2][42] ), .B(n282), .Z(n778) );
  ND3 U554 ( .A(n1006), .B(n1007), .C(n1008), .Z(\CARRYB[2][42] ) );
  EO U555 ( .A(\CARRYB[2][45] ), .B(n795), .Z(\SUMB[3][45] ) );
  EO U556 ( .A(\SUMB[2][46] ), .B(n285), .Z(n795) );
  ND2 U557 ( .A(\CARRYB[2][41] ), .B(n282), .Z(n779) );
  ND2 U558 ( .A(\SUMB[2][42] ), .B(\CARRYB[2][41] ), .Z(n777) );
  ND3 U559 ( .A(n1114), .B(n1115), .C(n1116), .Z(\CARRYB[5][39] ) );
  EO U560 ( .A(n1362), .B(n1359), .Z(\SUMB[1][34] ) );
  EO U561 ( .A(\SUMB[8][39] ), .B(n522), .Z(n1171) );
  ND2 U562 ( .A(\CARRYB[6][31] ), .B(\SUMB[6][32] ), .Z(n870) );
  EO U563 ( .A(n715), .B(n1361), .Z(\SUMB[1][31] ) );
  ND3 U564 ( .A(n886), .B(n887), .C(n888), .Z(\CARRYB[11][30] ) );
  ND3 U565 ( .A(n804), .B(n805), .C(n806), .Z(\CARRYB[8][30] ) );
  ND2 U566 ( .A(\SUMB[7][31] ), .B(n275), .Z(n806) );
  ND2 U567 ( .A(\CARRYB[7][30] ), .B(\SUMB[7][31] ), .Z(n804) );
  ND3 U568 ( .A(n816), .B(n817), .C(n818), .Z(\CARRYB[2][28] ) );
  ND3 U569 ( .A(n827), .B(n828), .C(n829), .Z(\CARRYB[15][36] ) );
  ND2 U570 ( .A(\CARRYB[14][36] ), .B(\SUMB[14][37] ), .Z(n827) );
  ND2 U571 ( .A(n770), .B(n771), .Z(\SUMB[2][28] ) );
  ND2 U572 ( .A(\CARRYB[1][28] ), .B(n769), .Z(n770) );
  ND3 U573 ( .A(n788), .B(n789), .C(n790), .Z(\CARRYB[18][38] ) );
  ND2 U574 ( .A(\CARRYB[17][38] ), .B(\SUMB[17][39] ), .Z(n788) );
  EO U575 ( .A(n1367), .B(n1408), .Z(\SUMB[1][26] ) );
  EO U576 ( .A(\CARRYB[17][38] ), .B(n787), .Z(\SUMB[18][38] ) );
  EO U577 ( .A(\SUMB[14][27] ), .B(n903), .Z(\SUMB[15][26] ) );
  ND3 U578 ( .A(n893), .B(n894), .C(n895), .Z(\CARRYB[4][23] ) );
  EO U579 ( .A(\SUMB[23][28] ), .B(n721), .Z(\SUMB[24][27] ) );
  EO U580 ( .A(\CARRYB[23][27] ), .B(\ab[27][24] ), .Z(n721) );
  ND3 U581 ( .A(n722), .B(n723), .C(n724), .Z(\CARRYB[24][27] ) );
  ND3 U582 ( .A(n799), .B(n800), .C(n801), .Z(\CARRYB[10][23] ) );
  EO U583 ( .A(\SUMB[9][24] ), .B(n758), .Z(\SUMB[10][23] ) );
  EO U584 ( .A(\CARRYB[9][23] ), .B(n561), .Z(n758) );
  EO U585 ( .A(\CARRYB[22][33] ), .B(n753), .Z(\SUMB[23][33] ) );
  EO U586 ( .A(\SUMB[22][34] ), .B(\ab[33][23] ), .Z(n753) );
  ND3 U587 ( .A(n754), .B(n755), .C(n756), .Z(\CARRYB[23][33] ) );
  EO U588 ( .A(\SUMB[18][25] ), .B(n877), .Z(\SUMB[19][24] ) );
  EO U589 ( .A(\SUMB[9][23] ), .B(n841), .Z(\SUMB[10][22] ) );
  EO U590 ( .A(\CARRYB[26][43] ), .B(n934), .Z(\SUMB[27][43] ) );
  EO U591 ( .A(\SUMB[26][44] ), .B(\ab[43][27] ), .Z(n934) );
  ND3 U592 ( .A(n935), .B(n936), .C(n937), .Z(\CARRYB[27][43] ) );
  ND2 U593 ( .A(\CARRYB[26][43] ), .B(\SUMB[26][44] ), .Z(n935) );
  EO U594 ( .A(n1338), .B(n1393), .Z(\SUMB[1][22] ) );
  ND2 U595 ( .A(\CARRYB[27][31] ), .B(\ab[31][28] ), .Z(n835) );
  ND2 U596 ( .A(\CARRYB[27][31] ), .B(\SUMB[27][32] ), .Z(n834) );
  EO U597 ( .A(\CARRYB[13][19] ), .B(n1020), .Z(\SUMB[14][19] ) );
  ND3 U598 ( .A(n1021), .B(n1022), .C(n1023), .Z(\CARRYB[14][19] ) );
  ND2 U599 ( .A(\CARRYB[13][19] ), .B(\SUMB[13][20] ), .Z(n1021) );
  ND3 U600 ( .A(n695), .B(n696), .C(n697), .Z(\CARRYB[30][32] ) );
  EO U601 ( .A(\CARRYB[22][18] ), .B(\ab[23][18] ), .Z(n860) );
  ND3 U602 ( .A(n773), .B(n774), .C(n775), .Z(\CARRYB[30][15] ) );
  ND2 U603 ( .A(\SUMB[29][16] ), .B(\CARRYB[29][15] ), .Z(n773) );
  ND3 U604 ( .A(n671), .B(n672), .C(n673), .Z(\CARRYB[14][16] ) );
  ND3 U605 ( .A(n992), .B(n993), .C(n994), .Z(\CARRYB[34][20] ) );
  EO U606 ( .A(\SUMB[29][16] ), .B(n772), .Z(\SUMB[30][15] ) );
  EO U607 ( .A(\CARRYB[29][15] ), .B(\ab[30][15] ), .Z(n772) );
  EO U608 ( .A(\SUMB[18][19] ), .B(n988), .Z(\SUMB[19][18] ) );
  EO U609 ( .A(\CARRYB[20][14] ), .B(n639), .Z(n717) );
  ND2 U610 ( .A(\CARRYB[35][28] ), .B(\ab[36][28] ), .Z(n1095) );
  ND2 U611 ( .A(\SUMB[35][29] ), .B(\CARRYB[35][28] ), .Z(n1093) );
  EO U612 ( .A(\CARRYB[26][13] ), .B(n918), .Z(\SUMB[27][13] ) );
  EO U613 ( .A(\SUMB[26][14] ), .B(n613), .Z(n918) );
  ND2 U614 ( .A(\CARRYB[22][13] ), .B(n619), .Z(n813) );
  ND3 U615 ( .A(n1050), .B(n1051), .C(n1052), .Z(\CARRYB[15][11] ) );
  ND2 U616 ( .A(\CARRYB[36][36] ), .B(\ab[37][36] ), .Z(n1119) );
  EO U617 ( .A(\CARRYB[36][36] ), .B(n1117), .Z(\SUMB[37][36] ) );
  EO U618 ( .A(\SUMB[36][37] ), .B(\ab[37][36] ), .Z(n1117) );
  ND3 U619 ( .A(n747), .B(n748), .C(n749), .Z(\CARRYB[34][11] ) );
  EO U620 ( .A(n1358), .B(n1354), .Z(\SUMB[1][12] ) );
  ND3 U621 ( .A(n809), .B(n810), .C(n811), .Z(\CARRYB[27][11] ) );
  ND2 U622 ( .A(\SUMB[26][12] ), .B(n543), .Z(n810) );
  EO U623 ( .A(\SUMB[25][13] ), .B(n830), .Z(\SUMB[26][12] ) );
  EO U624 ( .A(\CARRYB[25][12] ), .B(n595), .Z(n830) );
  EO U625 ( .A(\SUMB[14][12] ), .B(n585), .Z(n1049) );
  EO U626 ( .A(n1371), .B(n1346), .Z(\SUMB[1][10] ) );
  ND3 U627 ( .A(n1056), .B(n1057), .C(n1058), .Z(\CARRYB[40][38] ) );
  ND2 U628 ( .A(\SUMB[40][39] ), .B(\CARRYB[40][38] ), .Z(n1062) );
  EO U629 ( .A(n1059), .B(\CARRYB[40][38] ), .Z(\SUMB[41][38] ) );
  EO U630 ( .A(\ab[41][38] ), .B(\SUMB[40][39] ), .Z(n1059) );
  ND3 U631 ( .A(n1060), .B(n1061), .C(n1062), .Z(\CARRYB[41][38] ) );
  ND2 U632 ( .A(\ab[41][38] ), .B(\SUMB[40][39] ), .Z(n1060) );
  ND2 U633 ( .A(\ab[41][38] ), .B(\CARRYB[40][38] ), .Z(n1061) );
  EO U634 ( .A(\CARRYB[40][13] ), .B(n1045), .Z(\SUMB[41][13] ) );
  EO U635 ( .A(\SUMB[40][14] ), .B(\ab[41][13] ), .Z(n1045) );
  ND3 U636 ( .A(n999), .B(n1000), .C(n1001), .Z(\CARRYB[36][7] ) );
  ND2 U637 ( .A(n470), .B(\SUMB[35][8] ), .Z(n1000) );
  ND3 U638 ( .A(n1157), .B(n1158), .C(n1159), .Z(\CARRYB[22][7] ) );
  ND2 U639 ( .A(\CARRYB[21][7] ), .B(\SUMB[21][8] ), .Z(n1157) );
  ND2 U640 ( .A(\CARRYB[21][7] ), .B(n416), .Z(n1158) );
  EO U641 ( .A(n1385), .B(n1378), .Z(\SUMB[1][9] ) );
  ND3 U642 ( .A(n1089), .B(n1090), .C(n1091), .Z(\CARRYB[43][18] ) );
  ND3 U643 ( .A(n1078), .B(n1079), .C(n1080), .Z(\CARRYB[43][16] ) );
  ND3 U644 ( .A(n1295), .B(n1296), .C(n1297), .Z(\CARRYB[29][5] ) );
  IVP U645 ( .A(\ab[27][27] ), .Z(n1486) );
  EO U646 ( .A(\SUMB[13][8] ), .B(n459), .Z(n1160) );
  ND3 U647 ( .A(n1161), .B(n1162), .C(n1163), .Z(\CARRYB[14][7] ) );
  ND3 U648 ( .A(n1180), .B(n1181), .C(n1182), .Z(\CARRYB[5][5] ) );
  ND3 U649 ( .A(n1176), .B(n1177), .C(n1178), .Z(\CARRYB[45][4] ) );
  EO U650 ( .A(\CARRYB[28][5] ), .B(n1294), .Z(\SUMB[29][5] ) );
  EO U651 ( .A(\SUMB[28][6] ), .B(n1276), .Z(n1294) );
  ND3 U652 ( .A(n1017), .B(n1018), .C(n1019), .Z(\CARRYB[20][5] ) );
  IVP U653 ( .A(\ab[22][22] ), .Z(n1477) );
  IVP U654 ( .A(n1448), .Z(n1445) );
  ND3 U655 ( .A(n1132), .B(n1133), .C(n1134), .Z(\CARRYB[45][26] ) );
  ND3 U656 ( .A(n953), .B(n954), .C(n955), .Z(\CARRYB[46][31] ) );
  ND2 U657 ( .A(\CARRYB[45][31] ), .B(\SUMB[45][32] ), .Z(n953) );
  ND3 U658 ( .A(n1085), .B(n1086), .C(n1087), .Z(\CARRYB[29][3] ) );
  ND3 U659 ( .A(n1104), .B(n1105), .C(n1106), .Z(\CARRYB[7][3] ) );
  IVP U660 ( .A(\ab[4][4] ), .Z(n1444) );
  ND3 U661 ( .A(n915), .B(n916), .C(n917), .Z(\CARRYB[46][30] ) );
  EO U662 ( .A(\CARRYB[47][6] ), .B(\SUMB[47][7] ), .Z(\A1[52] ) );
  EO U663 ( .A(\CARRYB[47][2] ), .B(\SUMB[47][3] ), .Z(\A1[48] ) );
  EO U664 ( .A(\CARRYB[19][4] ), .B(n1231), .Z(\SUMB[20][4] ) );
  EO U665 ( .A(\SUMB[19][5] ), .B(n349), .Z(n1231) );
  ND2 U666 ( .A(\CARRYB[17][1] ), .B(n1329), .Z(n1150) );
  ND3 U667 ( .A(n1100), .B(n1101), .C(n1102), .Z(\CARRYB[12][3] ) );
  EO U668 ( .A(\CARRYB[11][3] ), .B(n1099), .Z(\SUMB[12][3] ) );
  EO U669 ( .A(\SUMB[11][4] ), .B(n346), .Z(n1099) );
  EO U670 ( .A(\CARRYB[6][3] ), .B(n1103), .Z(\SUMB[7][3] ) );
  EO U671 ( .A(\SUMB[6][4] ), .B(n345), .Z(n1103) );
  ND2 U672 ( .A(n1311), .B(\CARRYB[40][2] ), .Z(n1226) );
  ND2 U673 ( .A(n1311), .B(\SUMB[40][3] ), .Z(n1225) );
  EO U674 ( .A(\CARRYB[34][1] ), .B(n1262), .Z(\SUMB[35][1] ) );
  EO U675 ( .A(n1084), .B(\CARRYB[28][3] ), .Z(\SUMB[29][3] ) );
  EO U676 ( .A(n297), .B(\SUMB[28][4] ), .Z(n1084) );
  ND3 U677 ( .A(n1153), .B(n1154), .C(n1155), .Z(\CARRYB[23][1] ) );
  ND2 U678 ( .A(\CARRYB[22][1] ), .B(\SUMB[22][2] ), .Z(n1153) );
  ND2 U679 ( .A(\CARRYB[22][1] ), .B(n1420), .Z(n1154) );
  EO U680 ( .A(\CARRYB[10][2] ), .B(n1187), .Z(\SUMB[11][2] ) );
  EO U681 ( .A(\SUMB[10][3] ), .B(n312), .Z(n1187) );
  NR2 U682 ( .A(n1434), .B(n1249), .Z(\CARRYB[1][1] ) );
  ND3 U683 ( .A(n1218), .B(n1219), .C(n1220), .Z(\CARRYB[28][0] ) );
  EO U684 ( .A(\CARRYB[24][1] ), .B(n1258), .Z(\SUMB[25][1] ) );
  EO U685 ( .A(\CARRYB[22][1] ), .B(n1152), .Z(\SUMB[23][1] ) );
  EO U686 ( .A(\CARRYB[17][1] ), .B(n1148), .Z(\SUMB[18][1] ) );
  IVP U687 ( .A(\ab[33][33] ), .Z(n1499) );
  IVP U688 ( .A(\ab[29][29] ), .Z(n1492) );
  IVP U689 ( .A(\ab[11][11] ), .Z(n1458) );
  AN2P U690 ( .A(\ab[15][15] ), .B(\ab[1][1] ), .Z(n267) );
  IVP U691 ( .A(\ab[23][23] ), .Z(n1478) );
  IVP U692 ( .A(\ab[21][21] ), .Z(n1473) );
  IVP U693 ( .A(\ab[20][20] ), .Z(n1472) );
  IVP U694 ( .A(\ab[43][43] ), .Z(n1522) );
  IVP U695 ( .A(\ab[46][46] ), .Z(n1527) );
  IVP U696 ( .A(\ab[45][45] ), .Z(n1524) );
  AN2P U697 ( .A(A[21]), .B(\ab[1][1] ), .Z(n268) );
  AN2P U698 ( .A(n1507), .B(A[3]), .Z(n269) );
  AN2P U699 ( .A(n1435), .B(A[47]), .Z(n270) );
  AN2P U700 ( .A(A[2]), .B(A[47]), .Z(n271) );
  AN2P U701 ( .A(n1440), .B(A[47]), .Z(n272) );
  AN2P U702 ( .A(A[44]), .B(A[6]), .Z(n273) );
  AN2P U703 ( .A(n1445), .B(A[47]), .Z(n274) );
  AN2P U704 ( .A(A[30]), .B(A[8]), .Z(n275) );
  AN2P U705 ( .A(n1500), .B(A[8]), .Z(n276) );
  AN2P U706 ( .A(n1487), .B(A[8]), .Z(n277) );
  AN2P U707 ( .A(A[32]), .B(A[8]), .Z(n278) );
  AN2P U708 ( .A(n1521), .B(A[7]), .Z(n279) );
  AN2P U709 ( .A(n1475), .B(A[9]), .Z(n280) );
  AN2P U710 ( .A(n1475), .B(A[10]), .Z(n281) );
  IVP U711 ( .A(\ab[14][14] ), .Z(n1460) );
  AN2P U712 ( .A(A[41]), .B(A[3]), .Z(n282) );
  AN2P U713 ( .A(n1505), .B(A[3]), .Z(n283) );
  AN2P U714 ( .A(A[25]), .B(n1437), .Z(n284) );
  AN2P U715 ( .A(A[45]), .B(A[3]), .Z(n285) );
  AN2P U716 ( .A(A[28]), .B(n1437), .Z(n286) );
  AN2P U717 ( .A(A[23]), .B(n1436), .Z(n287) );
  AN2P U718 ( .A(n1512), .B(A[3]), .Z(n288) );
  AN2P U719 ( .A(\ab[36][36] ), .B(A[3]), .Z(n289) );
  AN2P U720 ( .A(A[30]), .B(n1433), .Z(n290) );
  AN2P U721 ( .A(n1469), .B(A[2]), .Z(n291) );
  AN2P U722 ( .A(n1485), .B(n1437), .Z(n292) );
  AN2P U723 ( .A(\ab[36][36] ), .B(A[2]), .Z(n293) );
  AN2P U724 ( .A(n1466), .B(A[2]), .Z(n294) );
  AN2P U725 ( .A(A[46]), .B(A[3]), .Z(n295) );
  AN2P U726 ( .A(\ab[31][31] ), .B(n1437), .Z(n296) );
  AN2P U727 ( .A(n1491), .B(n1437), .Z(n297) );
  AN2P U728 ( .A(n1502), .B(n1437), .Z(n298) );
  AN2P U729 ( .A(\ab[26][26] ), .B(A[2]), .Z(n299) );
  AN2P U730 ( .A(A[30]), .B(n1437), .Z(n300) );
  AN2P U731 ( .A(A[3]), .B(A[2]), .Z(n301) );
  AN2P U732 ( .A(A[23]), .B(A[2]), .Z(n302) );
  AN2P U733 ( .A(A[10]), .B(A[2]), .Z(n303) );
  AN2P U734 ( .A(A[45]), .B(\ab[1][1] ), .Z(n304) );
  AN2P U735 ( .A(\ab[34][34] ), .B(n1437), .Z(n305) );
  AN2P U736 ( .A(A[44]), .B(\B[0] ), .Z(n306) );
  AN2P U737 ( .A(n1480), .B(n1437), .Z(n307) );
  IVP U738 ( .A(\ab[24][24] ), .Z(n1481) );
  AN2P U739 ( .A(\ab[44][44] ), .B(A[2]), .Z(n308) );
  AN2P U740 ( .A(A[37]), .B(A[2]), .Z(n309) );
  AN2P U741 ( .A(A[22]), .B(\B[0] ), .Z(n310) );
  AN2P U742 ( .A(A[23]), .B(n1441), .Z(n311) );
  AN2P U743 ( .A(A[11]), .B(A[2]), .Z(n312) );
  AN2P U744 ( .A(n1474), .B(n1441), .Z(n313) );
  AN2P U745 ( .A(\ab[6][6] ), .B(n1435), .Z(n314) );
  AN2P U746 ( .A(\ab[6][6] ), .B(n1440), .Z(n315) );
  AN2P U747 ( .A(A[9]), .B(A[2]), .Z(n316) );
  AN2P U748 ( .A(A[13]), .B(A[2]), .Z(n317) );
  AN2P U749 ( .A(A[33]), .B(n1437), .Z(n318) );
  AN2P U750 ( .A(A[30]), .B(n1447), .Z(n319) );
  AN2P U751 ( .A(A[41]), .B(n1441), .Z(n320) );
  AN2P U752 ( .A(A[32]), .B(n1437), .Z(n321) );
  AN2P U753 ( .A(\ab[42][42] ), .B(n1441), .Z(n322) );
  AN2P U754 ( .A(n1511), .B(n1441), .Z(n323) );
  AN2P U755 ( .A(n1446), .B(n1435), .Z(n324) );
  AN2P U756 ( .A(\ab[6][6] ), .B(A[2]), .Z(n325) );
  AN2P U757 ( .A(A[8]), .B(n1435), .Z(n326) );
  AN2P U758 ( .A(A[25]), .B(A[2]), .Z(n327) );
  AN2P U759 ( .A(A[10]), .B(n1435), .Z(n328) );
  AN2P U760 ( .A(n1468), .B(n1436), .Z(n329) );
  AN2P U761 ( .A(A[21]), .B(n1436), .Z(n330) );
  AN2P U762 ( .A(A[11]), .B(n1435), .Z(n331) );
  AN2P U763 ( .A(A[12]), .B(A[2]), .Z(n332) );
  AN2P U764 ( .A(n1464), .B(n1436), .Z(n333) );
  AN2P U765 ( .A(n1525), .B(n1441), .Z(n334) );
  AN2P U766 ( .A(A[38]), .B(n1440), .Z(n335) );
  AN2P U767 ( .A(\ab[26][26] ), .B(n1437), .Z(n336) );
  AN2P U768 ( .A(n1520), .B(n1440), .Z(n337) );
  AN2P U769 ( .A(n1459), .B(n1436), .Z(n338) );
  AN2P U770 ( .A(A[30]), .B(n1442), .Z(n339) );
  AN2P U771 ( .A(A[8]), .B(A[2]), .Z(n340) );
  AN2P U772 ( .A(A[44]), .B(A[3]), .Z(n341) );
  AN2P U773 ( .A(A[14]), .B(A[2]), .Z(n342) );
  AN2P U774 ( .A(A[38]), .B(A[3]), .Z(n343) );
  AN2P U775 ( .A(n1523), .B(n1440), .Z(n344) );
  AN2P U776 ( .A(\ab[7][7] ), .B(n1435), .Z(n345) );
  AN2P U777 ( .A(A[12]), .B(n1436), .Z(n346) );
  AN2P U778 ( .A(A[9]), .B(n1435), .Z(n347) );
  AN2P U779 ( .A(\ab[7][7] ), .B(A[2]), .Z(n348) );
  IVP U780 ( .A(\ab[39][39] ), .Z(n1509) );
  IVP U781 ( .A(n1509), .Z(n1507) );
  IVP U782 ( .A(n1509), .Z(n1508) );
  AN2P U783 ( .A(\ab[20][20] ), .B(n1441), .Z(n349) );
  AN2P U784 ( .A(\ab[18][18] ), .B(n1441), .Z(n350) );
  AN2P U785 ( .A(n1489), .B(n1442), .Z(n351) );
  AN2P U786 ( .A(\ab[34][34] ), .B(n1442), .Z(n352) );
  AN2P U787 ( .A(A[33]), .B(n1442), .Z(n353) );
  AN2P U788 ( .A(A[44]), .B(n1441), .Z(n354) );
  AN2P U789 ( .A(n1508), .B(n1440), .Z(n355) );
  AN2P U790 ( .A(n1484), .B(n1442), .Z(n356) );
  AN2P U791 ( .A(A[25]), .B(n1441), .Z(n357) );
  AN2P U792 ( .A(n1442), .B(n1435), .Z(n358) );
  AN2P U793 ( .A(A[5]), .B(A[2]), .Z(n359) );
  AN2P U794 ( .A(A[13]), .B(n1436), .Z(n360) );
  AN2P U795 ( .A(\ab[16][16] ), .B(n1441), .Z(n361) );
  AN2P U796 ( .A(n1462), .B(n1441), .Z(n362) );
  AN2P U797 ( .A(A[21]), .B(n1441), .Z(n363) );
  AN2P U798 ( .A(\ab[26][26] ), .B(n1442), .Z(n364) );
  AN2P U799 ( .A(\ab[31][31] ), .B(n1442), .Z(n365) );
  AN2P U800 ( .A(A[14]), .B(n1441), .Z(n366) );
  AN2P U801 ( .A(\ab[36][36] ), .B(n1442), .Z(n367) );
  AN2P U802 ( .A(n1501), .B(n1442), .Z(n368) );
  AN2P U803 ( .A(\ab[7][7] ), .B(n1440), .Z(n369) );
  AN2P U804 ( .A(A[4]), .B(A[2]), .Z(n370) );
  AN2P U805 ( .A(n1475), .B(n1446), .Z(n371) );
  AN2P U806 ( .A(A[8]), .B(n1440), .Z(n372) );
  AN2P U807 ( .A(A[30]), .B(n1451), .Z(n373) );
  AN2P U808 ( .A(n1483), .B(n1446), .Z(n374) );
  AN2P U809 ( .A(A[9]), .B(n1440), .Z(n375) );
  AN2P U810 ( .A(A[32]), .B(n1442), .Z(n376) );
  AN2P U811 ( .A(n1510), .B(n1445), .Z(n377) );
  AN2P U812 ( .A(A[10]), .B(n1440), .Z(n378) );
  AN2P U813 ( .A(n1447), .B(n1440), .Z(n379) );
  AN2P U814 ( .A(A[12]), .B(n1440), .Z(n380) );
  AN2P U815 ( .A(A[11]), .B(n1440), .Z(n381) );
  AN2P U816 ( .A(n1500), .B(n1447), .Z(n382) );
  AN2P U817 ( .A(\ab[20][20] ), .B(n1446), .Z(n383) );
  AN2P U818 ( .A(n1507), .B(n1447), .Z(n384) );
  AN2P U819 ( .A(A[41]), .B(n1445), .Z(n385) );
  AN2P U820 ( .A(A[33]), .B(n1447), .Z(n386) );
  AN2P U821 ( .A(n1510), .B(n1451), .Z(n387) );
  AN2P U822 ( .A(n1526), .B(n1445), .Z(n388) );
  AN2P U823 ( .A(\ab[26][26] ), .B(n1446), .Z(n389) );
  AN2P U824 ( .A(A[32]), .B(n1447), .Z(n390) );
  AN2P U825 ( .A(A[13]), .B(n1440), .Z(n391) );
  AN2P U826 ( .A(\ab[34][34] ), .B(n1447), .Z(n392) );
  AN2P U827 ( .A(n1488), .B(n1447), .Z(n393) );
  AN2P U828 ( .A(A[23]), .B(n1446), .Z(n394) );
  AN2P U829 ( .A(A[32]), .B(n1451), .Z(n395) );
  AN2P U830 ( .A(n1487), .B(n1450), .Z(n396) );
  AN2P U831 ( .A(n1483), .B(n1450), .Z(n397) );
  AN2P U832 ( .A(\ab[18][18] ), .B(n1446), .Z(n398) );
  AN2P U833 ( .A(n1521), .B(n1445), .Z(n399) );
  AN2P U834 ( .A(A[21]), .B(n1446), .Z(n400) );
  AN2P U835 ( .A(n1523), .B(n1445), .Z(n401) );
  AN2P U836 ( .A(\ab[42][42] ), .B(n1445), .Z(n402) );
  AN2P U837 ( .A(\ab[31][31] ), .B(n1447), .Z(n403) );
  AN2P U838 ( .A(\ab[16][16] ), .B(n1446), .Z(n404) );
  AN2P U839 ( .A(A[25]), .B(n1450), .Z(n405) );
  AN2P U840 ( .A(A[25]), .B(n1446), .Z(n406) );
  AN2P U841 ( .A(\ab[36][36] ), .B(n1447), .Z(n407) );
  AN2P U842 ( .A(n1475), .B(n1450), .Z(n408) );
  AN2P U843 ( .A(n1500), .B(n1451), .Z(n409) );
  AN2P U844 ( .A(\ab[6][6] ), .B(n1445), .Z(n410) );
  AN2P U845 ( .A(A[30]), .B(n1455), .Z(n411) );
  AN2P U846 ( .A(A[11]), .B(n1445), .Z(n412) );
  AN2P U847 ( .A(n1461), .B(n1445), .Z(n413) );
  AN2P U848 ( .A(A[14]), .B(n1445), .Z(n414) );
  AN2P U849 ( .A(A[44]), .B(n1445), .Z(n415) );
  AN2P U850 ( .A(n1475), .B(n1454), .Z(n416) );
  AN2P U851 ( .A(n1500), .B(n1455), .Z(n417) );
  AN2P U852 ( .A(n1510), .B(n1455), .Z(n418) );
  AN2P U853 ( .A(A[25]), .B(n1454), .Z(n419) );
  AN2P U854 ( .A(\ab[6][6] ), .B(n1526), .Z(n420) );
  AN2P U855 ( .A(A[13]), .B(n1445), .Z(n421) );
  AN2P U856 ( .A(A[23]), .B(n1450), .Z(n422) );
  AN2P U857 ( .A(n1483), .B(n1454), .Z(n423) );
  AN2P U858 ( .A(n1487), .B(n1454), .Z(n424) );
  AN2P U859 ( .A(A[8]), .B(n1445), .Z(n425) );
  AN2P U860 ( .A(\ab[7][7] ), .B(n1445), .Z(n426) );
  AN2P U861 ( .A(A[9]), .B(n1445), .Z(n427) );
  AN2P U862 ( .A(\ab[18][18] ), .B(n1450), .Z(n428) );
  AN2P U863 ( .A(\ab[20][20] ), .B(n1450), .Z(n429) );
  AN2P U864 ( .A(\ab[34][34] ), .B(n1451), .Z(n430) );
  AN2P U865 ( .A(\ab[16][16] ), .B(n1449), .Z(n431) );
  AN2P U866 ( .A(n1507), .B(n1451), .Z(n432) );
  AN2P U867 ( .A(\ab[26][26] ), .B(n1450), .Z(n433) );
  AN2P U868 ( .A(A[33]), .B(n1451), .Z(n434) );
  AN2P U869 ( .A(n1523), .B(\ab[6][6] ), .Z(n435) );
  AN2P U870 ( .A(\ab[36][36] ), .B(n1451), .Z(n436) );
  AN2P U871 ( .A(A[10]), .B(n1445), .Z(n437) );
  AN2P U872 ( .A(A[14]), .B(n1449), .Z(n438) );
  AN2P U873 ( .A(A[21]), .B(n1450), .Z(n439) );
  AN2P U874 ( .A(A[32]), .B(n1455), .Z(n440) );
  AN2P U875 ( .A(A[12]), .B(n1445), .Z(n441) );
  AN2P U876 ( .A(n1461), .B(n1449), .Z(n442) );
  AN2P U877 ( .A(A[41]), .B(\ab[6][6] ), .Z(n443) );
  IVP U878 ( .A(\ab[6][6] ), .Z(n1452) );
  AN2P U879 ( .A(A[33]), .B(n1455), .Z(n445) );
  AN2P U880 ( .A(n1483), .B(A[8]), .Z(n446) );
  AN2P U881 ( .A(n1521), .B(\ab[6][6] ), .Z(n447) );
  AN2P U882 ( .A(n1465), .B(n1454), .Z(n448) );
  AN2P U883 ( .A(A[9]), .B(n1449), .Z(n449) );
  AN2P U884 ( .A(A[13]), .B(n1449), .Z(n450) );
  AN2P U885 ( .A(n1470), .B(n1454), .Z(n451) );
  AN2P U886 ( .A(n1475), .B(A[8]), .Z(n452) );
  AN2P U887 ( .A(\ab[31][31] ), .B(n1451), .Z(n453) );
  AN2P U888 ( .A(n1510), .B(A[8]), .Z(n454) );
  AN2P U889 ( .A(\ab[42][42] ), .B(\ab[6][6] ), .Z(n455) );
  AN2P U890 ( .A(A[8]), .B(n1449), .Z(n456) );
  AN2P U891 ( .A(A[11]), .B(n1449), .Z(n457) );
  AN2P U892 ( .A(\ab[20][20] ), .B(n1454), .Z(n458) );
  AN2P U893 ( .A(A[14]), .B(n1453), .Z(n459) );
  AN2P U894 ( .A(\ab[31][31] ), .B(n1455), .Z(n460) );
  AN2P U895 ( .A(A[37]), .B(n1455), .Z(n461) );
  AN2P U896 ( .A(A[30]), .B(A[9]), .Z(n462) );
  AN2P U897 ( .A(A[41]), .B(\ab[7][7] ), .Z(n463) );
  AN2P U898 ( .A(A[10]), .B(n1449), .Z(n464) );
  AN2P U899 ( .A(A[13]), .B(n1453), .Z(n465) );
  AN2P U900 ( .A(A[23]), .B(n1454), .Z(n466) );
  AN2P U901 ( .A(A[44]), .B(\ab[7][7] ), .Z(n467) );
  AN2P U902 ( .A(A[25]), .B(A[8]), .Z(n468) );
  AN2P U903 ( .A(A[21]), .B(n1454), .Z(n469) );
  AN2P U904 ( .A(\ab[36][36] ), .B(n1455), .Z(n470) );
  AN2P U905 ( .A(n1461), .B(n1453), .Z(n471) );
  AN2P U906 ( .A(\ab[26][26] ), .B(n1454), .Z(n472) );
  AN2P U907 ( .A(\ab[7][7] ), .B(n1523), .Z(n473) );
  AN2P U908 ( .A(\ab[18][18] ), .B(n1454), .Z(n474) );
  AN2P U909 ( .A(n1507), .B(n1455), .Z(n475) );
  AN2P U910 ( .A(A[12]), .B(n1449), .Z(n476) );
  AN2P U911 ( .A(\ab[34][34] ), .B(n1455), .Z(n477) );
  AN2P U912 ( .A(\ab[20][20] ), .B(A[8]), .Z(n478) );
  AN2P U913 ( .A(\ab[16][16] ), .B(n1453), .Z(n479) );
  AN2P U914 ( .A(\ab[7][7] ), .B(n1449), .Z(n480) );
  AN2P U915 ( .A(n1507), .B(A[8]), .Z(n482) );
  AN2P U916 ( .A(A[25]), .B(A[9]), .Z(n483) );
  AN2P U917 ( .A(n1470), .B(A[8]), .Z(n484) );
  AN2P U918 ( .A(\ab[31][31] ), .B(A[8]), .Z(n485) );
  AN2P U919 ( .A(A[37]), .B(A[8]), .Z(n486) );
  AN2P U920 ( .A(A[13]), .B(A[8]), .Z(n487) );
  AN2P U921 ( .A(\ab[34][34] ), .B(A[8]), .Z(n488) );
  AN2P U922 ( .A(A[33]), .B(A[8]), .Z(n489) );
  AN2P U923 ( .A(A[21]), .B(A[8]), .Z(n490) );
  AN2P U924 ( .A(n1483), .B(A[9]), .Z(n491) );
  AN2P U925 ( .A(n1461), .B(A[8]), .Z(n492) );
  AN2P U926 ( .A(A[8]), .B(n1453), .Z(n493) );
  AN2P U927 ( .A(A[11]), .B(n1453), .Z(n494) );
  AN2P U928 ( .A(A[14]), .B(A[8]), .Z(n495) );
  AN2P U929 ( .A(n1500), .B(A[9]), .Z(n496) );
  AN2P U930 ( .A(\ab[26][26] ), .B(A[8]), .Z(n497) );
  AN2P U931 ( .A(\ab[42][42] ), .B(\ab[7][7] ), .Z(n498) );
  AN2P U932 ( .A(A[23]), .B(A[8]), .Z(n499) );
  AN2P U933 ( .A(n1465), .B(A[8]), .Z(n500) );
  AN2P U934 ( .A(A[32]), .B(A[9]), .Z(n501) );
  AN2P U935 ( .A(n1487), .B(A[9]), .Z(n502) );
  AN2P U936 ( .A(A[10]), .B(n1453), .Z(n503) );
  IVP U937 ( .A(\ab[7][7] ), .Z(n1456) );
  AN2P U938 ( .A(\ab[18][18] ), .B(A[8]), .Z(n506) );
  AN2P U939 ( .A(A[30]), .B(A[10]), .Z(n507) );
  AN2P U940 ( .A(A[10]), .B(A[8]), .Z(n508) );
  AN2P U941 ( .A(A[29]), .B(A[9]), .Z(n509) );
  AN2P U942 ( .A(A[12]), .B(n1453), .Z(n510) );
  AN2P U943 ( .A(A[8]), .B(n1521), .Z(n511) );
  AN2P U944 ( .A(A[21]), .B(A[9]), .Z(n512) );
  AN2P U945 ( .A(n1479), .B(A[9]), .Z(n513) );
  AN2P U946 ( .A(A[9]), .B(n1453), .Z(n514) );
  AN2P U947 ( .A(n1465), .B(A[9]), .Z(n515) );
  AN2P U948 ( .A(A[33]), .B(A[9]), .Z(n516) );
  AN2P U949 ( .A(\ab[36][36] ), .B(A[8]), .Z(n517) );
  AN2P U950 ( .A(\ab[16][16] ), .B(A[8]), .Z(n518) );
  AN2P U951 ( .A(A[41]), .B(A[8]), .Z(n519) );
  AN2P U952 ( .A(n1483), .B(A[10]), .Z(n520) );
  AN2P U953 ( .A(A[23]), .B(A[9]), .Z(n521) );
  AN2P U954 ( .A(A[38]), .B(A[9]), .Z(n522) );
  AN2P U955 ( .A(\ab[26][26] ), .B(A[9]), .Z(n523) );
  AN2P U956 ( .A(\ab[31][31] ), .B(A[9]), .Z(n524) );
  AN2P U957 ( .A(\ab[20][20] ), .B(A[9]), .Z(n525) );
  AN2P U958 ( .A(A[9]), .B(A[8]), .Z(n526) );
  AN2P U959 ( .A(n1461), .B(A[9]), .Z(n527) );
  AN2P U960 ( .A(\ab[18][18] ), .B(A[9]), .Z(n528) );
  AN2P U961 ( .A(A[9]), .B(n1507), .Z(n529) );
  AN2P U962 ( .A(A[13]), .B(A[9]), .Z(n530) );
  AN2P U963 ( .A(n1468), .B(A[9]), .Z(n531) );
  AN2P U964 ( .A(n1500), .B(A[10]), .Z(n532) );
  AN2P U965 ( .A(A[11]), .B(A[8]), .Z(n533) );
  AN2P U966 ( .A(\ab[42][42] ), .B(A[8]), .Z(n534) );
  AN2P U967 ( .A(\ab[16][16] ), .B(A[9]), .Z(n535) );
  AN2P U968 ( .A(A[14]), .B(A[9]), .Z(n536) );
  AN2P U969 ( .A(\ab[36][36] ), .B(A[9]), .Z(n537) );
  AN2P U970 ( .A(A[12]), .B(A[8]), .Z(n538) );
  AN2P U971 ( .A(\ab[34][34] ), .B(A[9]), .Z(n539) );
  AN2P U972 ( .A(A[25]), .B(A[10]), .Z(n540) );
  AN2P U973 ( .A(A[33]), .B(A[10]), .Z(n542) );
  AN2P U974 ( .A(n1483), .B(A[11]), .Z(n543) );
  AN2P U975 ( .A(\ab[26][26] ), .B(A[10]), .Z(n544) );
  AN2P U976 ( .A(\ab[31][31] ), .B(A[10]), .Z(n545) );
  AN2P U977 ( .A(A[37]), .B(A[9]), .Z(n546) );
  AN2P U978 ( .A(A[21]), .B(A[10]), .Z(n547) );
  AN2P U979 ( .A(n1487), .B(A[10]), .Z(n548) );
  AN2P U980 ( .A(\ab[20][20] ), .B(A[10]), .Z(n549) );
  AN2P U981 ( .A(A[30]), .B(A[11]), .Z(n550) );
  AN2P U982 ( .A(A[32]), .B(A[10]), .Z(n551) );
  AN2P U983 ( .A(A[10]), .B(A[9]), .Z(n552) );
  AN2P U984 ( .A(A[12]), .B(A[9]), .Z(n553) );
  AN2P U985 ( .A(n1479), .B(A[10]), .Z(n554) );
  AN2P U986 ( .A(A[29]), .B(A[10]), .Z(n555) );
  AN2P U987 ( .A(n1465), .B(A[10]), .Z(n556) );
  AN2P U988 ( .A(\ab[18][18] ), .B(A[10]), .Z(n557) );
  AN2P U989 ( .A(n1461), .B(A[10]), .Z(n558) );
  AN2P U990 ( .A(\ab[16][16] ), .B(A[10]), .Z(n559) );
  AN2P U991 ( .A(n1470), .B(A[10]), .Z(n560) );
  AN2P U992 ( .A(A[23]), .B(A[10]), .Z(n561) );
  AN2P U993 ( .A(n1487), .B(A[11]), .Z(n562) );
  AN2P U994 ( .A(A[25]), .B(A[11]), .Z(n563) );
  AN2P U995 ( .A(\ab[34][34] ), .B(A[10]), .Z(n564) );
  AN2P U996 ( .A(n1475), .B(A[11]), .Z(n565) );
  AN2P U997 ( .A(A[13]), .B(A[10]), .Z(n566) );
  AN2P U998 ( .A(A[10]), .B(n1505), .Z(n567) );
  AN2P U999 ( .A(A[11]), .B(A[9]), .Z(n568) );
  AN2P U1000 ( .A(A[14]), .B(A[10]), .Z(n569) );
  AN2P U1001 ( .A(A[29]), .B(A[11]), .Z(n571) );
  AN2P U1002 ( .A(n1468), .B(A[11]), .Z(n572) );
  AN2P U1003 ( .A(A[33]), .B(A[11]), .Z(n573) );
  AN2P U1004 ( .A(\ab[36][36] ), .B(A[10]), .Z(n574) );
  AN2P U1005 ( .A(A[11]), .B(A[10]), .Z(n575) );
  AN2P U1006 ( .A(A[12]), .B(A[10]), .Z(n576) );
  AN2P U1007 ( .A(A[32]), .B(A[11]), .Z(n577) );
  AN2P U1008 ( .A(\ab[26][26] ), .B(A[11]), .Z(n578) );
  AN2P U1009 ( .A(n1496), .B(A[11]), .Z(n579) );
  AN2P U1010 ( .A(A[21]), .B(A[11]), .Z(n580) );
  AN2P U1011 ( .A(n1465), .B(A[11]), .Z(n581) );
  AN2P U1012 ( .A(A[23]), .B(A[11]), .Z(n582) );
  AN2P U1013 ( .A(A[11]), .B(\ab[34][34] ), .Z(n583) );
  AN2P U1014 ( .A(\ab[18][18] ), .B(A[11]), .Z(n584) );
  AN2P U1015 ( .A(n1461), .B(A[11]), .Z(n585) );
  AN2P U1016 ( .A(A[14]), .B(A[11]), .Z(n586) );
  AN2P U1017 ( .A(A[13]), .B(A[11]), .Z(n587) );
  AN2P U1018 ( .A(n1479), .B(A[11]), .Z(n588) );
  AN2P U1019 ( .A(\ab[16][16] ), .B(A[11]), .Z(n589) );
  AN2P U1020 ( .A(n1495), .B(A[12]), .Z(n591) );
  AN2P U1021 ( .A(n1489), .B(A[12]), .Z(n592) );
  AN2P U1022 ( .A(n1479), .B(A[12]), .Z(n593) );
  AN2P U1023 ( .A(n1476), .B(A[12]), .Z(n594) );
  AN2P U1024 ( .A(\ab[26][26] ), .B(A[12]), .Z(n595) );
  AN2P U1025 ( .A(A[21]), .B(A[12]), .Z(n596) );
  AN2P U1026 ( .A(A[20]), .B(A[12]), .Z(n597) );
  AN2P U1027 ( .A(A[30]), .B(A[12]), .Z(n598) );
  AN2P U1028 ( .A(\ab[18][18] ), .B(A[12]), .Z(n599) );
  AN2P U1029 ( .A(A[23]), .B(A[12]), .Z(n600) );
  AN2P U1030 ( .A(A[12]), .B(A[32]), .Z(n601) );
  AN2P U1031 ( .A(A[12]), .B(A[11]), .Z(n602) );
  AN2P U1032 ( .A(n1485), .B(A[12]), .Z(n603) );
  AN2P U1033 ( .A(A[13]), .B(A[12]), .Z(n604) );
  AN2P U1034 ( .A(n1470), .B(A[12]), .Z(n605) );
  AN2P U1035 ( .A(n1466), .B(A[12]), .Z(n608) );
  AN2P U1036 ( .A(A[29]), .B(A[12]), .Z(n609) );
  AN2P U1037 ( .A(A[25]), .B(A[12]), .Z(n610) );
  AN2P U1038 ( .A(A[14]), .B(A[12]), .Z(n611) );
  AN2P U1039 ( .A(A[16]), .B(A[12]), .Z(n612) );
  AN2P U1040 ( .A(n1485), .B(A[13]), .Z(n613) );
  AN2P U1041 ( .A(A[13]), .B(A[30]), .Z(n614) );
  AN2P U1042 ( .A(A[20]), .B(A[13]), .Z(n615) );
  AN2P U1043 ( .A(\ab[26][26] ), .B(A[13]), .Z(n616) );
  AN2P U1044 ( .A(n1462), .B(A[12]), .Z(n617) );
  AN2P U1045 ( .A(A[23]), .B(A[13]), .Z(n619) );
  AN2P U1046 ( .A(n1476), .B(A[13]), .Z(n620) );
  AN2P U1047 ( .A(A[29]), .B(A[13]), .Z(n621) );
  AN2P U1048 ( .A(A[14]), .B(A[13]), .Z(n622) );
  AN2P U1049 ( .A(\ab[18][18] ), .B(A[13]), .Z(n623) );
  AN2P U1050 ( .A(A[16]), .B(A[13]), .Z(n624) );
  AN2P U1051 ( .A(A[25]), .B(A[13]), .Z(n625) );
  AN2P U1052 ( .A(A[21]), .B(A[13]), .Z(n626) );
  AN2P U1053 ( .A(n1489), .B(A[13]), .Z(n627) );
  AN2P U1054 ( .A(n1462), .B(A[13]), .Z(n628) );
  AN2P U1055 ( .A(n1466), .B(A[13]), .Z(n629) );
  AN2P U1056 ( .A(n1470), .B(A[13]), .Z(n630) );
  AN2P U1057 ( .A(n1479), .B(A[13]), .Z(n631) );
  AN2P U1058 ( .A(A[25]), .B(A[14]), .Z(n635) );
  AN2P U1059 ( .A(n1470), .B(A[14]), .Z(n636) );
  AN2P U1060 ( .A(A[20]), .B(A[14]), .Z(n637) );
  AN2P U1061 ( .A(A[16]), .B(A[14]), .Z(n638) );
  AN2P U1062 ( .A(A[21]), .B(A[14]), .Z(n639) );
  AN2P U1063 ( .A(n1479), .B(A[14]), .Z(n640) );
  AN2P U1064 ( .A(n1462), .B(A[14]), .Z(n641) );
  AN2P U1065 ( .A(A[23]), .B(A[14]), .Z(n642) );
  AN2P U1066 ( .A(n1466), .B(A[14]), .Z(n643) );
  AN2P U1067 ( .A(\ab[18][18] ), .B(A[14]), .Z(n644) );
  AN2P U1068 ( .A(A[14]), .B(\ab[26][26] ), .Z(n645) );
  AN2P U1069 ( .A(n1476), .B(A[14]), .Z(n646) );
  IVP U1070 ( .A(\ab[15][15] ), .Z(n1463) );
  AN2P U1071 ( .A(A[21]), .B(\B[0] ), .Z(n651) );
  AN2P U1072 ( .A(\ab[31][31] ), .B(\B[0] ), .Z(n1342) );
  AN2 U1073 ( .A(\CARRYB[47][0] ), .B(\SUMB[47][1] ), .Z(\A2[47] ) );
  AN2 U1074 ( .A(n1534), .B(n1530), .Z(\CARRYB[1][2] ) );
  EO3P U1075 ( .A(\ab[31][29] ), .B(\CARRYB[28][31] ), .C(\SUMB[28][32] ), .Z(
        \SUMB[29][31] ) );
  ND2 U1076 ( .A(\ab[31][29] ), .B(\CARRYB[28][31] ), .Z(n654) );
  ND2 U1077 ( .A(\ab[31][29] ), .B(\SUMB[28][32] ), .Z(n655) );
  ND2 U1078 ( .A(\CARRYB[28][31] ), .B(\SUMB[28][32] ), .Z(n656) );
  ND3 U1079 ( .A(n654), .B(n655), .C(n656), .Z(\CARRYB[29][31] ) );
  ND2 U1080 ( .A(A[30]), .B(\CARRYB[29][30] ), .Z(n657) );
  ND2 U1081 ( .A(A[30]), .B(\SUMB[29][31] ), .Z(n658) );
  ND2 U1082 ( .A(\CARRYB[29][30] ), .B(\SUMB[29][31] ), .Z(n659) );
  EO3P U1083 ( .A(\CARRYB[19][36] ), .B(\ab[36][20] ), .C(\SUMB[19][37] ), .Z(
        \SUMB[20][36] ) );
  ND2 U1084 ( .A(\CARRYB[19][36] ), .B(\SUMB[19][37] ), .Z(n660) );
  ND2 U1085 ( .A(\CARRYB[19][36] ), .B(\ab[36][20] ), .Z(n661) );
  ND2 U1086 ( .A(\SUMB[19][37] ), .B(\ab[36][20] ), .Z(n662) );
  ND3 U1087 ( .A(n660), .B(n661), .C(n662), .Z(\CARRYB[20][36] ) );
  EOP U1088 ( .A(\CARRYB[7][39] ), .B(n482), .Z(n663) );
  EOP U1089 ( .A(\SUMB[7][40] ), .B(n663), .Z(\SUMB[8][39] ) );
  ND2 U1090 ( .A(\SUMB[7][40] ), .B(\CARRYB[7][39] ), .Z(n664) );
  ND2 U1091 ( .A(\SUMB[7][40] ), .B(n482), .Z(n665) );
  ND2 U1092 ( .A(\CARRYB[7][39] ), .B(n482), .Z(n666) );
  ND3P U1093 ( .A(n664), .B(n665), .C(n666), .Z(\CARRYB[8][39] ) );
  EO3P U1094 ( .A(\CARRYB[23][12] ), .B(n593), .C(\SUMB[23][13] ), .Z(
        \SUMB[24][12] ) );
  ND2 U1095 ( .A(\CARRYB[23][12] ), .B(\SUMB[23][13] ), .Z(n667) );
  ND2 U1096 ( .A(\CARRYB[23][12] ), .B(n593), .Z(n668) );
  ND2 U1097 ( .A(\SUMB[23][13] ), .B(n593), .Z(n669) );
  ND3 U1098 ( .A(n667), .B(n668), .C(n669), .Z(\CARRYB[24][12] ) );
  ND2 U1099 ( .A(\SUMB[13][17] ), .B(\CARRYB[13][16] ), .Z(n671) );
  ND2 U1100 ( .A(\SUMB[13][17] ), .B(n638), .Z(n672) );
  ND2 U1101 ( .A(\CARRYB[13][16] ), .B(n638), .Z(n673) );
  EO U1102 ( .A(\SUMB[3][21] ), .B(n674), .Z(\SUMB[4][20] ) );
  ND2 U1103 ( .A(\SUMB[3][21] ), .B(\CARRYB[3][20] ), .Z(n675) );
  ND2 U1104 ( .A(\SUMB[3][21] ), .B(n349), .Z(n676) );
  ND2 U1105 ( .A(\CARRYB[3][20] ), .B(n349), .Z(n677) );
  ND3 U1106 ( .A(n675), .B(n676), .C(n677), .Z(\CARRYB[4][20] ) );
  EO U1107 ( .A(\CARRYB[22][31] ), .B(\ab[31][23] ), .Z(n678) );
  EO U1108 ( .A(\SUMB[22][32] ), .B(n678), .Z(\SUMB[23][31] ) );
  ND2 U1109 ( .A(\SUMB[22][32] ), .B(\CARRYB[22][31] ), .Z(n679) );
  ND2 U1110 ( .A(\SUMB[22][32] ), .B(\ab[31][23] ), .Z(n680) );
  ND2 U1111 ( .A(\CARRYB[22][31] ), .B(\ab[31][23] ), .Z(n681) );
  ND3P U1112 ( .A(n679), .B(n680), .C(n681), .Z(\CARRYB[23][31] ) );
  EOP U1113 ( .A(\CARRYB[23][31] ), .B(\ab[31][24] ), .Z(n682) );
  EOP U1114 ( .A(\SUMB[23][32] ), .B(n682), .Z(\SUMB[24][31] ) );
  ND2 U1115 ( .A(\SUMB[23][32] ), .B(\CARRYB[23][31] ), .Z(n683) );
  ND2 U1116 ( .A(\SUMB[23][32] ), .B(\ab[31][24] ), .Z(n684) );
  ND2 U1117 ( .A(\CARRYB[23][31] ), .B(\ab[31][24] ), .Z(n685) );
  ND3 U1118 ( .A(n683), .B(n684), .C(n685), .Z(\CARRYB[24][31] ) );
  ND3P U1119 ( .A(n792), .B(n793), .C(n794), .Z(\CARRYB[2][46] ) );
  EOP U1120 ( .A(\CARRYB[23][16] ), .B(\ab[24][16] ), .Z(n686) );
  EOP U1121 ( .A(\SUMB[23][17] ), .B(n686), .Z(\SUMB[24][16] ) );
  ND2 U1122 ( .A(\SUMB[23][17] ), .B(\CARRYB[23][16] ), .Z(n687) );
  ND2 U1123 ( .A(\SUMB[23][17] ), .B(\ab[24][16] ), .Z(n688) );
  ND2 U1124 ( .A(\CARRYB[23][16] ), .B(\ab[24][16] ), .Z(n689) );
  ND3P U1125 ( .A(n687), .B(n688), .C(n689), .Z(\CARRYB[24][16] ) );
  ND2 U1126 ( .A(n1063), .B(n691), .Z(n692) );
  ND2 U1127 ( .A(n690), .B(\SUMB[2][24] ), .Z(n693) );
  IV U1128 ( .A(n1063), .Z(n690) );
  IVDA U1129 ( .A(\SUMB[2][24] ), .Y(n691) );
  NR2P U1130 ( .A(n1473), .B(n872), .Z(n1398) );
  ND2 U1131 ( .A(\CARRYB[29][13] ), .B(n614), .Z(n892) );
  ND2 U1132 ( .A(\CARRYB[29][32] ), .B(\SUMB[29][33] ), .Z(n695) );
  ND2 U1133 ( .A(\CARRYB[29][32] ), .B(\ab[32][30] ), .Z(n696) );
  ND2 U1134 ( .A(\SUMB[29][33] ), .B(\ab[32][30] ), .Z(n697) );
  ND2 U1135 ( .A(\SUMB[29][14] ), .B(n614), .Z(n891) );
  ND2 U1136 ( .A(\SUMB[29][14] ), .B(\CARRYB[29][13] ), .Z(n890) );
  ND2 U1137 ( .A(\SUMB[1][25] ), .B(n963), .Z(n964) );
  EOP U1138 ( .A(\CARRYB[23][21] ), .B(\ab[24][21] ), .Z(n698) );
  EOP U1139 ( .A(\SUMB[23][22] ), .B(n698), .Z(\SUMB[24][21] ) );
  ND2 U1140 ( .A(\SUMB[23][22] ), .B(\CARRYB[23][21] ), .Z(n699) );
  ND2 U1141 ( .A(\SUMB[23][22] ), .B(\ab[24][21] ), .Z(n700) );
  ND2 U1142 ( .A(\CARRYB[23][21] ), .B(\ab[24][21] ), .Z(n701) );
  ND3P U1143 ( .A(n699), .B(n700), .C(n701), .Z(\CARRYB[24][21] ) );
  EO3P U1144 ( .A(\CARRYB[6][20] ), .B(n458), .C(\SUMB[6][21] ), .Z(
        \SUMB[7][20] ) );
  ND2 U1145 ( .A(\CARRYB[6][20] ), .B(\SUMB[6][21] ), .Z(n702) );
  ND2 U1146 ( .A(\CARRYB[6][20] ), .B(n458), .Z(n703) );
  ND2 U1147 ( .A(\SUMB[6][21] ), .B(n458), .Z(n704) );
  ND3 U1148 ( .A(n702), .B(n703), .C(n704), .Z(\CARRYB[7][20] ) );
  ND2 U1149 ( .A(\CARRYB[22][16] ), .B(\SUMB[22][17] ), .Z(n705) );
  ND2 U1150 ( .A(\CARRYB[22][16] ), .B(\ab[23][16] ), .Z(n706) );
  ND2 U1151 ( .A(\SUMB[22][17] ), .B(\ab[23][16] ), .Z(n707) );
  ND3P U1152 ( .A(n705), .B(n706), .C(n707), .Z(\CARRYB[23][16] ) );
  EO3 U1153 ( .A(\SUMB[33][29] ), .B(\ab[34][28] ), .C(\CARRYB[33][28] ), .Z(
        \SUMB[34][28] ) );
  ND2P U1154 ( .A(\SUMB[33][29] ), .B(\CARRYB[33][28] ), .Z(n708) );
  ND2P U1155 ( .A(\SUMB[33][29] ), .B(\ab[34][28] ), .Z(n709) );
  ND2 U1156 ( .A(\CARRYB[33][28] ), .B(\ab[34][28] ), .Z(n710) );
  ND3P U1157 ( .A(n708), .B(n709), .C(n710), .Z(\CARRYB[34][28] ) );
  EOP U1158 ( .A(\SUMB[32][30] ), .B(n711), .Z(\SUMB[33][29] ) );
  ND2 U1159 ( .A(\SUMB[32][30] ), .B(\CARRYB[32][29] ), .Z(n712) );
  ND2 U1160 ( .A(\SUMB[32][30] ), .B(\ab[33][29] ), .Z(n713) );
  ND2 U1161 ( .A(\CARRYB[32][29] ), .B(\ab[33][29] ), .Z(n714) );
  ND3P U1162 ( .A(n712), .B(n713), .C(n714), .Z(\CARRYB[33][29] ) );
  EO U1163 ( .A(\CARRYB[14][11] ), .B(n1049), .Z(\SUMB[15][11] ) );
  AN2 U1164 ( .A(n1356), .B(n1350), .Z(\CARRYB[1][41] ) );
  AN2P U1165 ( .A(\ab[42][42] ), .B(\B[0] ), .Z(n1350) );
  ND3 U1166 ( .A(n949), .B(n950), .C(n951), .Z(\CARRYB[35][18] ) );
  NR2P U1167 ( .A(n1498), .B(n872), .Z(n715) );
  IVDA U1168 ( .A(n1363), .Z(n716) );
  ENP U1169 ( .A(n718), .B(n1300), .Z(n1016) );
  EO U1170 ( .A(n1366), .B(n1331), .Z(\SUMB[1][28] ) );
  B4IP U1171 ( .A(\ab[30][30] ), .Z(n719) );
  B4IP U1172 ( .A(\ab[30][30] ), .Z(n720) );
  AN2 U1173 ( .A(n1324), .B(n1396), .Z(\CARRYB[1][29] ) );
  EO3P U1174 ( .A(\CARRYB[2][25] ), .B(n284), .C(\SUMB[2][26] ), .Z(
        \SUMB[3][25] ) );
  ND2 U1175 ( .A(\SUMB[23][28] ), .B(\CARRYB[23][27] ), .Z(n722) );
  ND2 U1176 ( .A(\SUMB[23][28] ), .B(\ab[27][24] ), .Z(n723) );
  ND2 U1177 ( .A(\CARRYB[23][27] ), .B(\ab[27][24] ), .Z(n724) );
  NR2P U1178 ( .A(n1499), .B(n872), .Z(n1326) );
  NR2P U1179 ( .A(n1499), .B(n725), .Z(\CARRYB[1][33] ) );
  AN2P U1180 ( .A(\ab[31][31] ), .B(\ab[1][1] ), .Z(n726) );
  EOP U1181 ( .A(\CARRYB[21][13] ), .B(n620), .Z(n727) );
  EOP U1182 ( .A(\SUMB[21][14] ), .B(n727), .Z(\SUMB[22][13] ) );
  ND2 U1183 ( .A(\CARRYB[21][13] ), .B(n620), .Z(n730) );
  ND3P U1184 ( .A(n728), .B(n729), .C(n730), .Z(\CARRYB[22][13] ) );
  ND2 U1185 ( .A(\CARRYB[20][14] ), .B(\SUMB[20][15] ), .Z(n731) );
  ND2 U1186 ( .A(\CARRYB[20][14] ), .B(n639), .Z(n732) );
  ND2 U1187 ( .A(\SUMB[20][15] ), .B(n639), .Z(n733) );
  IVP U1188 ( .A(\ab[28][28] ), .Z(n1490) );
  B4IP U1189 ( .A(\ab[25][25] ), .Z(n736) );
  EO U1190 ( .A(\CARRYB[4][38] ), .B(n1273), .Z(n738) );
  EO U1191 ( .A(\SUMB[4][39] ), .B(n738), .Z(\SUMB[5][38] ) );
  ND2 U1192 ( .A(\SUMB[4][39] ), .B(\CARRYB[4][38] ), .Z(n739) );
  ND2 U1193 ( .A(\SUMB[4][39] ), .B(n1273), .Z(n740) );
  ND2 U1194 ( .A(\CARRYB[4][38] ), .B(n1273), .Z(n741) );
  IVP U1195 ( .A(\ab[40][40] ), .Z(n1513) );
  IVDA U1196 ( .A(n1355), .Z(n743) );
  EO3 U1197 ( .A(\CARRYB[24][32] ), .B(\ab[32][25] ), .C(\SUMB[24][33] ), .Z(
        \SUMB[25][32] ) );
  ND2 U1198 ( .A(\CARRYB[24][32] ), .B(\SUMB[24][33] ), .Z(n744) );
  ND2 U1199 ( .A(\CARRYB[24][32] ), .B(\ab[32][25] ), .Z(n745) );
  ND2 U1200 ( .A(\SUMB[24][33] ), .B(\ab[32][25] ), .Z(n746) );
  ND3 U1201 ( .A(n744), .B(n745), .C(n746), .Z(\CARRYB[25][32] ) );
  EO3P U1202 ( .A(\CARRYB[33][11] ), .B(n583), .C(\SUMB[33][12] ), .Z(
        \SUMB[34][11] ) );
  ND2 U1203 ( .A(\CARRYB[33][11] ), .B(\SUMB[33][12] ), .Z(n747) );
  ND2 U1204 ( .A(\CARRYB[33][11] ), .B(n583), .Z(n748) );
  ND2 U1205 ( .A(\SUMB[33][12] ), .B(n583), .Z(n749) );
  EO3 U1206 ( .A(\CARRYB[27][17] ), .B(\ab[28][17] ), .C(\SUMB[27][18] ), .Z(
        \SUMB[28][17] ) );
  ND2 U1207 ( .A(\CARRYB[27][17] ), .B(\SUMB[27][18] ), .Z(n750) );
  ND2 U1208 ( .A(\CARRYB[27][17] ), .B(\ab[28][17] ), .Z(n751) );
  ND2 U1209 ( .A(\SUMB[27][18] ), .B(\ab[28][17] ), .Z(n752) );
  ND3P U1210 ( .A(n750), .B(n751), .C(n752), .Z(\CARRYB[28][17] ) );
  ND2 U1211 ( .A(\CARRYB[22][33] ), .B(\SUMB[22][34] ), .Z(n754) );
  ND2 U1212 ( .A(\CARRYB[22][33] ), .B(\ab[33][23] ), .Z(n755) );
  ND2 U1213 ( .A(\SUMB[22][34] ), .B(\ab[33][23] ), .Z(n756) );
  IVDA U1214 ( .A(n1361), .Z(n757) );
  EO U1215 ( .A(\CARRYB[34][4] ), .B(n1135), .Z(\SUMB[35][4] ) );
  EO U1216 ( .A(\SUMB[34][5] ), .B(n368), .Z(n1135) );
  ND3 U1217 ( .A(n1140), .B(n1141), .C(n1142), .Z(\CARRYB[18][6] ) );
  AN2 U1218 ( .A(n1360), .B(n1399), .Z(n759) );
  EO U1219 ( .A(\CARRYB[12][31] ), .B(\ab[31][13] ), .Z(n760) );
  EO U1220 ( .A(\SUMB[12][32] ), .B(n760), .Z(\SUMB[13][31] ) );
  ND2 U1221 ( .A(\SUMB[12][32] ), .B(\CARRYB[12][31] ), .Z(n761) );
  ND2 U1222 ( .A(\SUMB[12][32] ), .B(\ab[31][13] ), .Z(n762) );
  ND2 U1223 ( .A(\CARRYB[12][31] ), .B(\ab[31][13] ), .Z(n763) );
  ND3P U1224 ( .A(n761), .B(n762), .C(n763), .Z(\CARRYB[13][31] ) );
  EOP U1225 ( .A(\CARRYB[11][28] ), .B(n592), .Z(n764) );
  ND2 U1226 ( .A(\SUMB[11][29] ), .B(\CARRYB[11][28] ), .Z(n765) );
  ND2 U1227 ( .A(\SUMB[11][29] ), .B(n592), .Z(n766) );
  ND2 U1228 ( .A(\CARRYB[11][28] ), .B(n592), .Z(n767) );
  ND3 U1229 ( .A(n765), .B(n766), .C(n767), .Z(\CARRYB[12][28] ) );
  AN2P U1230 ( .A(n1347), .B(n1352), .Z(\CARRYB[1][39] ) );
  ND2 U1231 ( .A(n768), .B(n815), .Z(n771) );
  IVDA U1232 ( .A(\CARRYB[1][28] ), .Y(n768) );
  IVP U1233 ( .A(n815), .Z(n769) );
  ND2P U1234 ( .A(\SUMB[29][16] ), .B(\ab[30][15] ), .Z(n774) );
  ND2 U1235 ( .A(\CARRYB[29][15] ), .B(\ab[30][15] ), .Z(n775) );
  AN2P U1236 ( .A(A[43]), .B(A[2]), .Z(n1302) );
  EO3 U1237 ( .A(\SUMB[2][42] ), .B(n282), .C(\CARRYB[2][41] ), .Z(
        \SUMB[3][41] ) );
  ND2 U1238 ( .A(\SUMB[18][25] ), .B(\ab[24][19] ), .Z(n879) );
  ND2 U1239 ( .A(\SUMB[18][25] ), .B(\CARRYB[18][24] ), .Z(n878) );
  EO3P U1240 ( .A(\SUMB[1][41] ), .B(n1319), .C(\CARRYB[1][40] ), .Z(
        \SUMB[2][40] ) );
  ND2P U1241 ( .A(\SUMB[1][41] ), .B(n1319), .Z(n781) );
  ND2P U1242 ( .A(\CARRYB[1][40] ), .B(n1319), .Z(n782) );
  ND3P U1243 ( .A(n780), .B(n781), .C(n782), .Z(\CARRYB[2][40] ) );
  EOP U1244 ( .A(\CARRYB[10][41] ), .B(\ab[41][11] ), .Z(n783) );
  EOP U1245 ( .A(\SUMB[10][42] ), .B(n783), .Z(\SUMB[11][41] ) );
  ND2 U1246 ( .A(\SUMB[10][42] ), .B(\CARRYB[10][41] ), .Z(n784) );
  ND2 U1247 ( .A(\SUMB[10][42] ), .B(\ab[41][11] ), .Z(n785) );
  ND2 U1248 ( .A(\CARRYB[10][41] ), .B(\ab[41][11] ), .Z(n786) );
  ND3P U1249 ( .A(n784), .B(n785), .C(n786), .Z(\CARRYB[11][41] ) );
  EOP U1250 ( .A(\SUMB[17][39] ), .B(\ab[38][18] ), .Z(n787) );
  ND2 U1251 ( .A(\SUMB[17][39] ), .B(\ab[38][18] ), .Z(n790) );
  EO U1252 ( .A(n1308), .B(n1343), .Z(n791) );
  EOP U1253 ( .A(\CARRYB[1][46] ), .B(n791), .Z(\SUMB[2][46] ) );
  ND2 U1254 ( .A(\CARRYB[1][46] ), .B(n1308), .Z(n792) );
  ND2 U1255 ( .A(\CARRYB[1][46] ), .B(n1343), .Z(n793) );
  ND2 U1256 ( .A(n1308), .B(n1343), .Z(n794) );
  ND2 U1257 ( .A(\CARRYB[2][45] ), .B(\SUMB[2][46] ), .Z(n796) );
  ND2 U1258 ( .A(\CARRYB[2][45] ), .B(n285), .Z(n797) );
  ND2 U1259 ( .A(\SUMB[2][46] ), .B(n285), .Z(n798) );
  ND2 U1260 ( .A(\SUMB[9][24] ), .B(\CARRYB[9][23] ), .Z(n799) );
  ND2 U1261 ( .A(\SUMB[9][24] ), .B(n561), .Z(n800) );
  ND2 U1262 ( .A(\CARRYB[9][23] ), .B(n561), .Z(n801) );
  AN2P U1263 ( .A(A[36]), .B(A[0]), .Z(n1363) );
  AN2 U1264 ( .A(n1393), .B(n1338), .Z(\CARRYB[1][22] ) );
  ND2 U1265 ( .A(\SUMB[26][12] ), .B(\CARRYB[26][11] ), .Z(n809) );
  EO3 U1266 ( .A(\CARRYB[7][30] ), .B(n275), .C(\SUMB[7][31] ), .Z(
        \SUMB[8][30] ) );
  ND2P U1267 ( .A(\CARRYB[7][30] ), .B(n275), .Z(n805) );
  NR2 U1268 ( .A(n1514), .B(n1400), .Z(n1356) );
  B4IP U1269 ( .A(\ab[1][1] ), .Z(n807) );
  EOP U1270 ( .A(\CARRYB[26][11] ), .B(n543), .Z(n808) );
  EOP U1271 ( .A(n808), .B(\SUMB[26][12] ), .Z(\SUMB[27][11] ) );
  ND2 U1272 ( .A(\CARRYB[26][11] ), .B(n543), .Z(n811) );
  EO3P U1273 ( .A(\CARRYB[22][13] ), .B(n619), .C(\SUMB[22][14] ), .Z(
        \SUMB[23][13] ) );
  ND2 U1274 ( .A(\CARRYB[22][13] ), .B(\SUMB[22][14] ), .Z(n812) );
  ND2 U1275 ( .A(\SUMB[22][14] ), .B(n619), .Z(n814) );
  ND3 U1276 ( .A(n812), .B(n813), .C(n814), .Z(\CARRYB[23][13] ) );
  EOP U1277 ( .A(\SUMB[1][29] ), .B(n1309), .Z(n815) );
  ND2 U1278 ( .A(\CARRYB[1][28] ), .B(\SUMB[1][29] ), .Z(n816) );
  ND2 U1279 ( .A(\CARRYB[1][28] ), .B(n1309), .Z(n817) );
  ND2 U1280 ( .A(\SUMB[1][29] ), .B(n1309), .Z(n818) );
  EO3 U1281 ( .A(\CARRYB[18][25] ), .B(\ab[25][19] ), .C(\SUMB[18][26] ), .Z(
        \SUMB[19][25] ) );
  ND2 U1282 ( .A(\CARRYB[18][25] ), .B(\SUMB[18][26] ), .Z(n819) );
  ND2 U1283 ( .A(\CARRYB[18][25] ), .B(\ab[25][19] ), .Z(n820) );
  ND2 U1284 ( .A(\SUMB[18][26] ), .B(\ab[25][19] ), .Z(n821) );
  ND3 U1285 ( .A(n819), .B(n820), .C(n821), .Z(\CARRYB[19][25] ) );
  EOP U1286 ( .A(n1396), .B(n1324), .Z(\SUMB[1][29] ) );
  NR2P U1287 ( .A(n1504), .B(n1411), .Z(n1403) );
  EOP U1288 ( .A(\CARRYB[33][24] ), .B(\ab[34][24] ), .Z(n822) );
  EOP U1289 ( .A(\SUMB[33][25] ), .B(n822), .Z(\SUMB[34][24] ) );
  ND2 U1290 ( .A(\SUMB[33][25] ), .B(\CARRYB[33][24] ), .Z(n823) );
  ND2 U1291 ( .A(\SUMB[33][25] ), .B(\ab[34][24] ), .Z(n824) );
  ND2 U1292 ( .A(\CARRYB[33][24] ), .B(\ab[34][24] ), .Z(n825) );
  ND3P U1293 ( .A(n823), .B(n824), .C(n825), .Z(\CARRYB[34][24] ) );
  EOP U1294 ( .A(\SUMB[14][37] ), .B(\ab[36][15] ), .Z(n826) );
  EOP U1295 ( .A(\CARRYB[14][36] ), .B(n826), .Z(\SUMB[15][36] ) );
  ND2 U1296 ( .A(\SUMB[14][37] ), .B(\ab[36][15] ), .Z(n829) );
  EO3P U1297 ( .A(\CARRYB[12][35] ), .B(\ab[35][13] ), .C(\SUMB[12][36] ), .Z(
        \SUMB[13][35] ) );
  ND2 U1298 ( .A(\SUMB[25][13] ), .B(\CARRYB[25][12] ), .Z(n831) );
  ND2 U1299 ( .A(\SUMB[25][13] ), .B(n595), .Z(n832) );
  ND2 U1300 ( .A(\CARRYB[25][12] ), .B(n595), .Z(n833) );
  ND3 U1301 ( .A(n831), .B(n832), .C(n833), .Z(\CARRYB[26][12] ) );
  ND3P U1302 ( .A(n939), .B(n940), .C(n941), .Z(\CARRYB[13][35] ) );
  EO3 U1303 ( .A(\CARRYB[27][31] ), .B(\ab[31][28] ), .C(\SUMB[27][32] ), .Z(
        \SUMB[28][31] ) );
  ND2 U1304 ( .A(\SUMB[27][32] ), .B(\ab[31][28] ), .Z(n836) );
  ND3P U1305 ( .A(n834), .B(n835), .C(n836), .Z(\CARRYB[28][31] ) );
  EO3P U1306 ( .A(\CARRYB[18][33] ), .B(\ab[33][19] ), .C(\SUMB[18][34] ), .Z(
        \SUMB[19][33] ) );
  ND2P U1307 ( .A(\CARRYB[18][33] ), .B(\SUMB[18][34] ), .Z(n837) );
  ND2P U1308 ( .A(\CARRYB[18][33] ), .B(\ab[33][19] ), .Z(n838) );
  ND2 U1309 ( .A(\SUMB[18][34] ), .B(\ab[33][19] ), .Z(n839) );
  ND3P U1310 ( .A(n837), .B(n838), .C(n839), .Z(\CARRYB[19][33] ) );
  ND3 U1311 ( .A(n981), .B(n982), .C(n983), .Z(\CARRYB[20][33] ) );
  EO3 U1312 ( .A(\SUMB[24][35] ), .B(\ab[34][25] ), .C(\CARRYB[24][34] ), .Z(
        \SUMB[25][34] ) );
  EOP U1313 ( .A(\CARRYB[9][22] ), .B(n281), .Z(n841) );
  ND2 U1314 ( .A(\SUMB[9][23] ), .B(\CARRYB[9][22] ), .Z(n842) );
  ND2 U1315 ( .A(\SUMB[9][23] ), .B(n281), .Z(n843) );
  ND2 U1316 ( .A(\CARRYB[9][22] ), .B(n281), .Z(n844) );
  ND3 U1317 ( .A(n842), .B(n843), .C(n844), .Z(\CARRYB[10][22] ) );
  EOP U1318 ( .A(\CARRYB[15][20] ), .B(\ab[20][16] ), .Z(n845) );
  EOP U1319 ( .A(\SUMB[15][21] ), .B(n845), .Z(\SUMB[16][20] ) );
  ND2 U1320 ( .A(\SUMB[15][21] ), .B(\CARRYB[15][20] ), .Z(n846) );
  ND2 U1321 ( .A(\SUMB[15][21] ), .B(\ab[20][16] ), .Z(n847) );
  ND2 U1322 ( .A(\CARRYB[15][20] ), .B(\ab[20][16] ), .Z(n848) );
  ND3P U1323 ( .A(n846), .B(n847), .C(n848), .Z(\CARRYB[16][20] ) );
  ND3P U1324 ( .A(n1122), .B(n1123), .C(n1124), .Z(\CARRYB[37][2] ) );
  EOP U1325 ( .A(\CARRYB[26][33] ), .B(\ab[33][27] ), .Z(n849) );
  EOP U1326 ( .A(\SUMB[26][34] ), .B(n849), .Z(\SUMB[27][33] ) );
  ND2 U1327 ( .A(\SUMB[26][34] ), .B(\CARRYB[26][33] ), .Z(n850) );
  ND2 U1328 ( .A(\SUMB[26][34] ), .B(\ab[33][27] ), .Z(n851) );
  ND2 U1329 ( .A(\CARRYB[26][33] ), .B(\ab[33][27] ), .Z(n852) );
  ND3P U1330 ( .A(n850), .B(n851), .C(n852), .Z(\CARRYB[27][33] ) );
  ND2 U1331 ( .A(\SUMB[24][35] ), .B(\CARRYB[24][34] ), .Z(n853) );
  ND2 U1332 ( .A(\CARRYB[24][34] ), .B(\ab[34][25] ), .Z(n855) );
  EO3 U1333 ( .A(\CARRYB[20][30] ), .B(\ab[30][21] ), .C(\SUMB[20][31] ), .Z(
        \SUMB[21][30] ) );
  EOP U1334 ( .A(\SUMB[32][17] ), .B(\ab[33][16] ), .Z(n856) );
  EOP U1335 ( .A(\CARRYB[32][16] ), .B(n856), .Z(\SUMB[33][16] ) );
  ND2 U1336 ( .A(\CARRYB[32][16] ), .B(\SUMB[32][17] ), .Z(n857) );
  ND2 U1337 ( .A(\CARRYB[32][16] ), .B(\ab[33][16] ), .Z(n858) );
  ND2 U1338 ( .A(\SUMB[32][17] ), .B(\ab[33][16] ), .Z(n859) );
  ND3 U1339 ( .A(n857), .B(n858), .C(n859), .Z(\CARRYB[33][16] ) );
  ND2 U1340 ( .A(\SUMB[22][19] ), .B(\CARRYB[22][18] ), .Z(n861) );
  ND2 U1341 ( .A(\SUMB[22][19] ), .B(\ab[23][18] ), .Z(n862) );
  ND2 U1342 ( .A(\CARRYB[22][18] ), .B(\ab[23][18] ), .Z(n863) );
  ND3 U1343 ( .A(n861), .B(n862), .C(n863), .Z(\CARRYB[23][18] ) );
  EO3P U1344 ( .A(\CARRYB[5][32] ), .B(n395), .C(\SUMB[5][33] ), .Z(
        \SUMB[6][32] ) );
  EOP U1345 ( .A(n460), .B(\CARRYB[6][31] ), .Z(n864) );
  EOP U1346 ( .A(n864), .B(\SUMB[6][32] ), .Z(\SUMB[7][31] ) );
  ND2 U1347 ( .A(n395), .B(\CARRYB[5][32] ), .Z(n865) );
  ND2 U1348 ( .A(n460), .B(\CARRYB[6][31] ), .Z(n868) );
  ND2P U1349 ( .A(n460), .B(\SUMB[6][32] ), .Z(n869) );
  ND3P U1350 ( .A(n868), .B(n869), .C(n870), .Z(\CARRYB[7][31] ) );
  NR2P U1351 ( .A(n1498), .B(n872), .Z(n871) );
  B4IP U1352 ( .A(\B[0] ), .Z(n872) );
  EOP U1353 ( .A(\CARRYB[30][12] ), .B(n591), .Z(n873) );
  ND2P U1354 ( .A(\SUMB[30][13] ), .B(n591), .Z(n875) );
  ND2 U1355 ( .A(\CARRYB[30][12] ), .B(n591), .Z(n876) );
  ND3P U1356 ( .A(n874), .B(n875), .C(n876), .Z(\CARRYB[31][12] ) );
  EOP U1357 ( .A(\CARRYB[18][24] ), .B(\ab[24][19] ), .Z(n877) );
  ND2 U1358 ( .A(\CARRYB[18][24] ), .B(\ab[24][19] ), .Z(n880) );
  EOP U1359 ( .A(n1342), .B(n1405), .Z(\SUMB[1][30] ) );
  EOP U1360 ( .A(\CARRYB[37][14] ), .B(\ab[38][14] ), .Z(n881) );
  EOP U1361 ( .A(\SUMB[37][15] ), .B(n881), .Z(\SUMB[38][14] ) );
  ND2 U1362 ( .A(\SUMB[37][15] ), .B(\CARRYB[37][14] ), .Z(n882) );
  ND2 U1363 ( .A(\SUMB[37][15] ), .B(\ab[38][14] ), .Z(n883) );
  ND2 U1364 ( .A(\CARRYB[37][14] ), .B(\ab[38][14] ), .Z(n884) );
  ND3P U1365 ( .A(n882), .B(n883), .C(n884), .Z(\CARRYB[38][14] ) );
  EOP U1366 ( .A(\CARRYB[10][30] ), .B(n550), .Z(n885) );
  EOP U1367 ( .A(\SUMB[10][31] ), .B(n885), .Z(\SUMB[11][30] ) );
  ND2 U1368 ( .A(\SUMB[10][31] ), .B(\CARRYB[10][30] ), .Z(n886) );
  ND2 U1369 ( .A(\SUMB[10][31] ), .B(n550), .Z(n887) );
  ND2 U1370 ( .A(\CARRYB[10][30] ), .B(n550), .Z(n888) );
  EO U1371 ( .A(\SUMB[9][39] ), .B(n910), .Z(\SUMB[10][38] ) );
  EOP U1372 ( .A(\CARRYB[29][13] ), .B(n614), .Z(n889) );
  EOP U1373 ( .A(\SUMB[29][14] ), .B(n889), .Z(\SUMB[30][13] ) );
  ND3P U1374 ( .A(n890), .B(n891), .C(n892), .Z(\CARRYB[30][13] ) );
  EO3P U1375 ( .A(\SUMB[3][24] ), .B(n311), .C(\CARRYB[3][23] ), .Z(
        \SUMB[4][23] ) );
  ND2 U1376 ( .A(\SUMB[3][24] ), .B(\CARRYB[3][23] ), .Z(n893) );
  ND2 U1377 ( .A(\SUMB[3][24] ), .B(n311), .Z(n894) );
  ND2 U1378 ( .A(\CARRYB[3][23] ), .B(n311), .Z(n895) );
  AN2 U1379 ( .A(n1408), .B(n1367), .Z(\CARRYB[1][26] ) );
  EO3P U1380 ( .A(\SUMB[26][22] ), .B(\ab[27][21] ), .C(\CARRYB[26][21] ), .Z(
        \SUMB[27][21] ) );
  ND2 U1381 ( .A(\SUMB[26][22] ), .B(\CARRYB[26][21] ), .Z(n896) );
  ND2 U1382 ( .A(\SUMB[26][22] ), .B(\ab[27][21] ), .Z(n897) );
  ND2 U1383 ( .A(\CARRYB[26][21] ), .B(\ab[27][21] ), .Z(n898) );
  ND3 U1384 ( .A(n896), .B(n897), .C(n898), .Z(\CARRYB[27][21] ) );
  EO3 U1385 ( .A(\CARRYB[14][30] ), .B(\ab[30][15] ), .C(\SUMB[14][31] ), .Z(
        \SUMB[15][30] ) );
  ND2 U1386 ( .A(\SUMB[14][31] ), .B(\ab[30][15] ), .Z(n902) );
  ND3P U1387 ( .A(n900), .B(n901), .C(n902), .Z(\CARRYB[15][30] ) );
  IVP U1388 ( .A(\ab[35][35] ), .Z(n1503) );
  IVP U1389 ( .A(n1503), .Z(n1502) );
  ND2 U1390 ( .A(\CARRYB[20][34] ), .B(\SUMB[20][35] ), .Z(n931) );
  EOP U1391 ( .A(\CARRYB[14][26] ), .B(\ab[26][15] ), .Z(n903) );
  ND2 U1392 ( .A(\SUMB[14][27] ), .B(\CARRYB[14][26] ), .Z(n904) );
  ND2 U1393 ( .A(\SUMB[14][27] ), .B(\ab[26][15] ), .Z(n905) );
  ND2 U1394 ( .A(\CARRYB[14][26] ), .B(\ab[26][15] ), .Z(n906) );
  ND3P U1395 ( .A(n904), .B(n905), .C(n906), .Z(\CARRYB[15][26] ) );
  AN2P U1396 ( .A(\ab[16][16] ), .B(\B[0] ), .Z(n1395) );
  EO3 U1397 ( .A(\CARRYB[31][24] ), .B(\ab[32][24] ), .C(\SUMB[31][25] ), .Z(
        \SUMB[32][24] ) );
  ND2 U1398 ( .A(\CARRYB[31][24] ), .B(\SUMB[31][25] ), .Z(n907) );
  ND2 U1399 ( .A(\CARRYB[31][24] ), .B(\ab[32][24] ), .Z(n908) );
  ND2 U1400 ( .A(\SUMB[31][25] ), .B(\ab[32][24] ), .Z(n909) );
  ND3P U1401 ( .A(n907), .B(n908), .C(n909), .Z(\CARRYB[32][24] ) );
  ND3P U1402 ( .A(n989), .B(n990), .C(n991), .Z(\CARRYB[19][18] ) );
  AN2P U1403 ( .A(\ab[27][27] ), .B(\B[0] ), .Z(n1367) );
  IV U1404 ( .A(\SUMB[1][25] ), .Z(n962) );
  AN2 U1405 ( .A(n1412), .B(n1337), .Z(\CARRYB[1][25] ) );
  EO U1406 ( .A(\CARRYB[8][38] ), .B(n1171), .Z(\SUMB[9][38] ) );
  EO U1407 ( .A(\CARRYB[37][39] ), .B(n975), .Z(\SUMB[38][39] ) );
  EOP U1408 ( .A(\CARRYB[9][38] ), .B(\ab[38][10] ), .Z(n910) );
  ND2 U1409 ( .A(\SUMB[9][39] ), .B(\CARRYB[9][38] ), .Z(n911) );
  ND2 U1410 ( .A(\SUMB[9][39] ), .B(\ab[38][10] ), .Z(n912) );
  ND2 U1411 ( .A(\CARRYB[9][38] ), .B(\ab[38][10] ), .Z(n913) );
  ND2 U1412 ( .A(\SUMB[45][31] ), .B(\CARRYB[45][30] ), .Z(n915) );
  ND2 U1413 ( .A(\SUMB[45][31] ), .B(\ab[46][30] ), .Z(n916) );
  ND2 U1414 ( .A(\CARRYB[45][30] ), .B(\ab[46][30] ), .Z(n917) );
  ND2 U1415 ( .A(\CARRYB[26][13] ), .B(\SUMB[26][14] ), .Z(n919) );
  ND2 U1416 ( .A(\CARRYB[26][13] ), .B(n613), .Z(n920) );
  ND2 U1417 ( .A(\SUMB[26][14] ), .B(n613), .Z(n921) );
  ND2 U1418 ( .A(\CARRYB[29][6] ), .B(\SUMB[29][7] ), .Z(n922) );
  ND2 U1419 ( .A(\CARRYB[29][6] ), .B(n373), .Z(n923) );
  ND2 U1420 ( .A(\SUMB[29][7] ), .B(n373), .Z(n924) );
  EO3 U1421 ( .A(\CARRYB[32][10] ), .B(n542), .C(\SUMB[32][11] ), .Z(
        \SUMB[33][10] ) );
  ND2 U1422 ( .A(\CARRYB[32][10] ), .B(\SUMB[32][11] ), .Z(n925) );
  ND2 U1423 ( .A(\CARRYB[32][10] ), .B(n542), .Z(n926) );
  ND2 U1424 ( .A(\SUMB[32][11] ), .B(n542), .Z(n927) );
  EO3 U1425 ( .A(\SUMB[17][38] ), .B(\ab[37][18] ), .C(\CARRYB[17][37] ), .Z(
        \SUMB[18][37] ) );
  ND2 U1426 ( .A(\CARRYB[17][37] ), .B(\SUMB[17][38] ), .Z(n928) );
  ND2 U1427 ( .A(\CARRYB[17][37] ), .B(\ab[37][18] ), .Z(n929) );
  ND2 U1428 ( .A(\SUMB[17][38] ), .B(\ab[37][18] ), .Z(n930) );
  ND3 U1429 ( .A(n928), .B(n929), .C(n930), .Z(\CARRYB[18][37] ) );
  ND2P U1430 ( .A(\CARRYB[20][34] ), .B(\ab[34][21] ), .Z(n932) );
  ND2 U1431 ( .A(\SUMB[20][35] ), .B(\ab[34][21] ), .Z(n933) );
  ND2P U1432 ( .A(\CARRYB[26][43] ), .B(\ab[43][27] ), .Z(n936) );
  ND2 U1433 ( .A(\SUMB[26][44] ), .B(\ab[43][27] ), .Z(n937) );
  EO U1434 ( .A(\CARRYB[34][18] ), .B(\ab[35][18] ), .Z(n938) );
  EO U1435 ( .A(\SUMB[34][19] ), .B(n938), .Z(\SUMB[35][18] ) );
  ND2 U1436 ( .A(\CARRYB[12][35] ), .B(\SUMB[12][36] ), .Z(n939) );
  ND2 U1437 ( .A(\CARRYB[12][35] ), .B(\ab[35][13] ), .Z(n940) );
  ND2 U1438 ( .A(\SUMB[12][36] ), .B(\ab[35][13] ), .Z(n941) );
  EO3 U1439 ( .A(\CARRYB[34][22] ), .B(\ab[35][22] ), .C(\SUMB[34][23] ), .Z(
        \SUMB[35][22] ) );
  ND2 U1440 ( .A(\CARRYB[34][22] ), .B(\SUMB[34][23] ), .Z(n942) );
  ND2 U1441 ( .A(\CARRYB[34][22] ), .B(\ab[35][22] ), .Z(n943) );
  ND2 U1442 ( .A(\SUMB[34][23] ), .B(\ab[35][22] ), .Z(n944) );
  ND3P U1443 ( .A(n942), .B(n943), .C(n944), .Z(\CARRYB[35][22] ) );
  EOP U1444 ( .A(\SUMB[24][15] ), .B(n635), .Z(n945) );
  EOP U1445 ( .A(\CARRYB[24][14] ), .B(n945), .Z(\SUMB[25][14] ) );
  ND2 U1446 ( .A(\CARRYB[24][14] ), .B(\SUMB[24][15] ), .Z(n946) );
  ND2 U1447 ( .A(\CARRYB[24][14] ), .B(n635), .Z(n947) );
  ND2 U1448 ( .A(\SUMB[24][15] ), .B(n635), .Z(n948) );
  ND3 U1449 ( .A(n946), .B(n947), .C(n948), .Z(\CARRYB[25][14] ) );
  ND2 U1450 ( .A(\CARRYB[34][18] ), .B(\SUMB[34][19] ), .Z(n949) );
  ND2 U1451 ( .A(\CARRYB[34][18] ), .B(\ab[35][18] ), .Z(n950) );
  ND2 U1452 ( .A(\SUMB[34][19] ), .B(\ab[35][18] ), .Z(n951) );
  EOP U1453 ( .A(\SUMB[45][32] ), .B(\ab[46][31] ), .Z(n952) );
  EOP U1454 ( .A(\CARRYB[45][31] ), .B(n952), .Z(\SUMB[46][31] ) );
  ND2P U1455 ( .A(\CARRYB[45][31] ), .B(\ab[46][31] ), .Z(n954) );
  ND2 U1456 ( .A(\SUMB[45][32] ), .B(\ab[46][31] ), .Z(n955) );
  EO3 U1457 ( .A(\CARRYB[36][21] ), .B(\ab[37][21] ), .C(\SUMB[36][22] ), .Z(
        \SUMB[37][21] ) );
  ND2 U1458 ( .A(\CARRYB[36][21] ), .B(\SUMB[36][22] ), .Z(n956) );
  ND2 U1459 ( .A(\CARRYB[36][21] ), .B(\ab[37][21] ), .Z(n957) );
  ND2 U1460 ( .A(\SUMB[36][22] ), .B(\ab[37][21] ), .Z(n958) );
  ND2 U1461 ( .A(\CARRYB[20][30] ), .B(\SUMB[20][31] ), .Z(n959) );
  ND2 U1462 ( .A(\CARRYB[20][30] ), .B(\ab[30][21] ), .Z(n960) );
  ND2 U1463 ( .A(\SUMB[20][31] ), .B(\ab[30][21] ), .Z(n961) );
  ND3P U1464 ( .A(n959), .B(n960), .C(n961), .Z(\CARRYB[21][30] ) );
  ND2 U1465 ( .A(n962), .B(n1016), .Z(n965) );
  ND2P U1466 ( .A(n964), .B(n965), .Z(\SUMB[2][24] ) );
  IVP U1467 ( .A(n1016), .Z(n963) );
  EOP U1468 ( .A(\CARRYB[15][13] ), .B(n624), .Z(n966) );
  EOP U1469 ( .A(\SUMB[15][14] ), .B(n966), .Z(\SUMB[16][13] ) );
  ND2P U1470 ( .A(n608), .B(\SUMB[16][13] ), .Z(n1075) );
  ND2P U1471 ( .A(\CARRYB[16][12] ), .B(\SUMB[16][13] ), .Z(n1076) );
  EOP U1472 ( .A(\CARRYB[22][15] ), .B(n967), .Z(\SUMB[23][15] ) );
  ND2 U1473 ( .A(\CARRYB[22][15] ), .B(\SUMB[22][16] ), .Z(n968) );
  ND2 U1474 ( .A(\CARRYB[22][15] ), .B(\ab[23][15] ), .Z(n969) );
  ND2 U1475 ( .A(\SUMB[22][16] ), .B(\ab[23][15] ), .Z(n970) );
  EOP U1476 ( .A(\SUMB[20][17] ), .B(\ab[21][16] ), .Z(n971) );
  EOP U1477 ( .A(\CARRYB[20][16] ), .B(n971), .Z(\SUMB[21][16] ) );
  ND2 U1478 ( .A(\CARRYB[20][16] ), .B(\SUMB[20][17] ), .Z(n972) );
  ND2 U1479 ( .A(\CARRYB[20][16] ), .B(\ab[21][16] ), .Z(n973) );
  ND2 U1480 ( .A(\SUMB[20][17] ), .B(\ab[21][16] ), .Z(n974) );
  ND3 U1481 ( .A(n972), .B(n973), .C(n974), .Z(\CARRYB[21][16] ) );
  ND2 U1482 ( .A(\CARRYB[37][39] ), .B(\SUMB[37][40] ), .Z(n976) );
  ND2 U1483 ( .A(\CARRYB[37][39] ), .B(\ab[39][38] ), .Z(n977) );
  ND2 U1484 ( .A(\SUMB[37][40] ), .B(\ab[39][38] ), .Z(n978) );
  ND3P U1485 ( .A(n976), .B(n977), .C(n978), .Z(\CARRYB[38][39] ) );
  EOP U1486 ( .A(\CARRYB[19][33] ), .B(\ab[33][20] ), .Z(n980) );
  EOP U1487 ( .A(\SUMB[19][34] ), .B(n980), .Z(\SUMB[20][33] ) );
  ND2 U1488 ( .A(\SUMB[19][34] ), .B(\CARRYB[19][33] ), .Z(n981) );
  ND2 U1489 ( .A(\SUMB[19][34] ), .B(\ab[33][20] ), .Z(n982) );
  ND2 U1490 ( .A(\CARRYB[19][33] ), .B(\ab[33][20] ), .Z(n983) );
  EOP U1491 ( .A(\SUMB[28][8] ), .B(n1287), .Z(n984) );
  EOP U1492 ( .A(\CARRYB[28][7] ), .B(n984), .Z(\SUMB[29][7] ) );
  ND2 U1493 ( .A(\CARRYB[28][7] ), .B(\SUMB[28][8] ), .Z(n985) );
  ND2 U1494 ( .A(\CARRYB[28][7] ), .B(n1287), .Z(n986) );
  ND2 U1495 ( .A(\SUMB[28][8] ), .B(n1287), .Z(n987) );
  EOP U1496 ( .A(\CARRYB[18][18] ), .B(\ab[19][18] ), .Z(n988) );
  ND2 U1497 ( .A(\SUMB[18][19] ), .B(\CARRYB[18][18] ), .Z(n989) );
  ND2 U1498 ( .A(\SUMB[18][19] ), .B(\ab[19][18] ), .Z(n990) );
  ND2 U1499 ( .A(\CARRYB[18][18] ), .B(\ab[19][18] ), .Z(n991) );
  EO3 U1500 ( .A(\CARRYB[33][20] ), .B(\ab[34][20] ), .C(\SUMB[33][21] ), .Z(
        \SUMB[34][20] ) );
  ND2 U1501 ( .A(\CARRYB[33][20] ), .B(\SUMB[33][21] ), .Z(n992) );
  ND2 U1502 ( .A(\CARRYB[33][20] ), .B(\ab[34][20] ), .Z(n993) );
  ND2 U1503 ( .A(\SUMB[33][21] ), .B(\ab[34][20] ), .Z(n994) );
  EO3P U1504 ( .A(n276), .B(\CARRYB[34][8] ), .C(\SUMB[34][9] ), .Z(
        \SUMB[35][8] ) );
  EOP U1505 ( .A(n470), .B(\CARRYB[35][7] ), .Z(n995) );
  EOP U1506 ( .A(n995), .B(\SUMB[35][8] ), .Z(\SUMB[36][7] ) );
  ND2 U1507 ( .A(n276), .B(\CARRYB[34][8] ), .Z(n996) );
  ND2 U1508 ( .A(n276), .B(\SUMB[34][9] ), .Z(n997) );
  ND2 U1509 ( .A(\CARRYB[34][8] ), .B(\SUMB[34][9] ), .Z(n998) );
  ND2 U1510 ( .A(n470), .B(\CARRYB[35][7] ), .Z(n999) );
  ND2 U1511 ( .A(n1325), .B(n1003), .Z(n1004) );
  ND2 U1512 ( .A(n1002), .B(n1419), .Z(n1005) );
  ND2 U1513 ( .A(n1004), .B(n1005), .Z(\SUMB[1][23] ) );
  IV U1514 ( .A(n1419), .Z(n1003) );
  AN2P U1515 ( .A(\ab[24][24] ), .B(\B[0] ), .Z(n1325) );
  NR2P U1516 ( .A(n1478), .B(n1400), .Z(n1419) );
  EO3P U1517 ( .A(\SUMB[1][43] ), .B(n1328), .C(\CARRYB[1][42] ), .Z(
        \SUMB[2][42] ) );
  ND2 U1518 ( .A(\CARRYB[1][42] ), .B(\SUMB[1][43] ), .Z(n1006) );
  ND2 U1519 ( .A(\CARRYB[1][42] ), .B(n1328), .Z(n1007) );
  ND2 U1520 ( .A(\SUMB[1][43] ), .B(n1328), .Z(n1008) );
  EOP U1521 ( .A(n306), .B(n1422), .Z(\SUMB[1][43] ) );
  EOP U1522 ( .A(\SUMB[10][35] ), .B(n1009), .Z(\SUMB[11][34] ) );
  ND2P U1523 ( .A(\SUMB[10][35] ), .B(\CARRYB[10][34] ), .Z(n1010) );
  ND2P U1524 ( .A(\SUMB[10][35] ), .B(n583), .Z(n1011) );
  ND2 U1525 ( .A(\CARRYB[10][34] ), .B(n583), .Z(n1012) );
  ND3P U1526 ( .A(n1010), .B(n1011), .C(n1012), .Z(\CARRYB[11][34] ) );
  EO3 U1527 ( .A(\CARRYB[2][37] ), .B(n283), .C(\SUMB[2][38] ), .Z(
        \SUMB[3][37] ) );
  ND2P U1528 ( .A(\CARRYB[2][37] ), .B(\SUMB[2][38] ), .Z(n1013) );
  ND2P U1529 ( .A(\CARRYB[2][37] ), .B(n283), .Z(n1014) );
  ND3P U1530 ( .A(n1013), .B(n1014), .C(n1015), .Z(\CARRYB[3][37] ) );
  EO3 U1531 ( .A(\CARRYB[19][5] ), .B(n383), .C(\SUMB[19][6] ), .Z(
        \SUMB[20][5] ) );
  ND2 U1532 ( .A(\CARRYB[19][5] ), .B(\SUMB[19][6] ), .Z(n1017) );
  ND2 U1533 ( .A(\CARRYB[19][5] ), .B(n383), .Z(n1018) );
  ND2 U1534 ( .A(\SUMB[19][6] ), .B(n383), .Z(n1019) );
  ND2P U1535 ( .A(\CARRYB[13][19] ), .B(n636), .Z(n1022) );
  ND2 U1536 ( .A(\SUMB[13][20] ), .B(n636), .Z(n1023) );
  ND2 U1537 ( .A(\CARRYB[19][35] ), .B(\SUMB[19][36] ), .Z(n1024) );
  ND2 U1538 ( .A(\CARRYB[19][35] ), .B(\ab[35][20] ), .Z(n1025) );
  ND2 U1539 ( .A(\SUMB[19][36] ), .B(\ab[35][20] ), .Z(n1026) );
  ND3 U1540 ( .A(n1024), .B(n1025), .C(n1026), .Z(\CARRYB[20][35] ) );
  ND2 U1541 ( .A(\CARRYB[2][25] ), .B(\SUMB[2][26] ), .Z(n1027) );
  ND2 U1542 ( .A(\CARRYB[2][25] ), .B(n284), .Z(n1028) );
  ND2 U1543 ( .A(\SUMB[2][26] ), .B(n284), .Z(n1029) );
  ND3 U1544 ( .A(n1027), .B(n1028), .C(n1029), .Z(\CARRYB[3][25] ) );
  EO U1545 ( .A(\SUMB[37][1] ), .B(n1374), .Z(n1030) );
  EO U1546 ( .A(\CARRYB[37][0] ), .B(n1030), .Z(\A1[36] ) );
  ND2 U1547 ( .A(\CARRYB[37][0] ), .B(\SUMB[37][1] ), .Z(n1031) );
  ND2 U1548 ( .A(\CARRYB[37][0] ), .B(n1374), .Z(n1032) );
  ND2 U1549 ( .A(\SUMB[37][1] ), .B(n1374), .Z(n1033) );
  AN2P U1550 ( .A(\ab[38][38] ), .B(\B[0] ), .Z(n1374) );
  ND2 U1551 ( .A(\CARRYB[28][9] ), .B(\SUMB[28][10] ), .Z(n1034) );
  ND2 U1552 ( .A(\CARRYB[28][9] ), .B(n509), .Z(n1035) );
  ND2 U1553 ( .A(\SUMB[28][10] ), .B(n509), .Z(n1036) );
  ND2 U1554 ( .A(\CARRYB[12][40] ), .B(\SUMB[12][41] ), .Z(n1038) );
  ND2 U1555 ( .A(\CARRYB[12][40] ), .B(\ab[40][13] ), .Z(n1039) );
  ND2 U1556 ( .A(\SUMB[12][41] ), .B(\ab[40][13] ), .Z(n1040) );
  ND3P U1557 ( .A(n1038), .B(n1039), .C(n1040), .Z(\CARRYB[13][40] ) );
  EOP U1558 ( .A(\CARRYB[17][11] ), .B(n584), .Z(n1041) );
  EOP U1559 ( .A(\SUMB[17][12] ), .B(n1041), .Z(\SUMB[18][11] ) );
  ND2P U1560 ( .A(\SUMB[17][12] ), .B(\CARRYB[17][11] ), .Z(n1042) );
  ND2P U1561 ( .A(\SUMB[17][12] ), .B(n584), .Z(n1043) );
  ND2 U1562 ( .A(\CARRYB[17][11] ), .B(n584), .Z(n1044) );
  ND3P U1563 ( .A(n1042), .B(n1043), .C(n1044), .Z(\CARRYB[18][11] ) );
  ND2 U1564 ( .A(\CARRYB[40][13] ), .B(\SUMB[40][14] ), .Z(n1046) );
  ND2 U1565 ( .A(\CARRYB[40][13] ), .B(\ab[41][13] ), .Z(n1047) );
  ND2 U1566 ( .A(\SUMB[40][14] ), .B(\ab[41][13] ), .Z(n1048) );
  ND3 U1567 ( .A(n1046), .B(n1047), .C(n1048), .Z(\CARRYB[41][13] ) );
  ND2 U1568 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(n1050) );
  ND2 U1569 ( .A(\CARRYB[14][11] ), .B(n585), .Z(n1051) );
  ND2 U1570 ( .A(\SUMB[14][12] ), .B(n585), .Z(n1052) );
  EO3 U1571 ( .A(\CARRYB[30][1] ), .B(n757), .C(\SUMB[30][2] ), .Z(
        \SUMB[31][1] ) );
  ND2 U1572 ( .A(\CARRYB[30][1] ), .B(\SUMB[30][2] ), .Z(n1053) );
  ND2 U1573 ( .A(\CARRYB[30][1] ), .B(n757), .Z(n1054) );
  ND2 U1574 ( .A(\SUMB[30][2] ), .B(n726), .Z(n1055) );
  ND2 U1575 ( .A(\ab[40][38] ), .B(\CARRYB[39][38] ), .Z(n1056) );
  ND2 U1576 ( .A(\ab[40][38] ), .B(\SUMB[39][39] ), .Z(n1057) );
  ND2 U1577 ( .A(\CARRYB[39][38] ), .B(\SUMB[39][39] ), .Z(n1058) );
  EOP U1578 ( .A(n287), .B(\CARRYB[2][23] ), .Z(n1063) );
  ND2 U1579 ( .A(n1300), .B(n759), .Z(n1064) );
  ND2 U1580 ( .A(n1300), .B(\SUMB[1][25] ), .Z(n1065) );
  ND2 U1581 ( .A(n759), .B(\SUMB[1][25] ), .Z(n1066) );
  ND3 U1582 ( .A(n1064), .B(n1065), .C(n1066), .Z(\CARRYB[2][24] ) );
  ND2P U1583 ( .A(n287), .B(\SUMB[2][24] ), .Z(n1068) );
  ND2P U1584 ( .A(\CARRYB[2][23] ), .B(\SUMB[2][24] ), .Z(n1069) );
  ND3P U1585 ( .A(n1067), .B(n1068), .C(n1069), .Z(\CARRYB[3][23] ) );
  EOP U1586 ( .A(n1070), .B(\SUMB[16][13] ), .Z(\SUMB[17][12] ) );
  ND2 U1587 ( .A(n624), .B(\CARRYB[15][13] ), .Z(n1071) );
  ND2 U1588 ( .A(n624), .B(\SUMB[15][14] ), .Z(n1072) );
  ND2 U1589 ( .A(\CARRYB[15][13] ), .B(\SUMB[15][14] ), .Z(n1073) );
  ND3 U1590 ( .A(n1071), .B(n1072), .C(n1073), .Z(\CARRYB[16][13] ) );
  ND2 U1591 ( .A(n608), .B(\CARRYB[16][12] ), .Z(n1074) );
  ND3P U1592 ( .A(n1074), .B(n1075), .C(n1076), .Z(\CARRYB[17][12] ) );
  EOP U1593 ( .A(\CARRYB[42][16] ), .B(\ab[43][16] ), .Z(n1077) );
  ND2 U1594 ( .A(\SUMB[42][17] ), .B(\CARRYB[42][16] ), .Z(n1078) );
  ND2 U1595 ( .A(\SUMB[42][17] ), .B(\ab[43][16] ), .Z(n1079) );
  ND2 U1596 ( .A(\CARRYB[42][16] ), .B(\ab[43][16] ), .Z(n1080) );
  EO3P U1597 ( .A(n286), .B(\CARRYB[27][3] ), .C(\SUMB[27][4] ), .Z(
        \SUMB[28][3] ) );
  ND3P U1598 ( .A(n1081), .B(n1082), .C(n1083), .Z(\CARRYB[28][3] ) );
  ND2 U1599 ( .A(n297), .B(\SUMB[28][4] ), .Z(n1085) );
  ND2 U1600 ( .A(n297), .B(\CARRYB[28][3] ), .Z(n1086) );
  ND2 U1601 ( .A(\SUMB[28][4] ), .B(\CARRYB[28][3] ), .Z(n1087) );
  ND2 U1602 ( .A(\CARRYB[42][18] ), .B(\SUMB[42][19] ), .Z(n1089) );
  ND2 U1603 ( .A(\CARRYB[42][18] ), .B(\ab[43][18] ), .Z(n1090) );
  ND2 U1604 ( .A(\SUMB[42][19] ), .B(\ab[43][18] ), .Z(n1091) );
  ND2P U1605 ( .A(\SUMB[35][29] ), .B(\ab[36][28] ), .Z(n1094) );
  AN2P U1606 ( .A(n304), .B(n1336), .Z(\CARRYB[1][45] ) );
  B4IP U1607 ( .A(\ab[1][1] ), .Z(n1411) );
  AN2P U1608 ( .A(A[26]), .B(\B[0] ), .Z(n1337) );
  EOP U1609 ( .A(n1363), .B(n1355), .Z(\SUMB[1][35] ) );
  EOP U1610 ( .A(\CARRYB[47][29] ), .B(\SUMB[47][30] ), .Z(\A1[75] ) );
  EOP U1611 ( .A(n1386), .B(n1381), .Z(\SUMB[1][7] ) );
  EOP U1612 ( .A(n1374), .B(n1345), .Z(\SUMB[1][37] ) );
  EOP U1613 ( .A(\CARRYB[3][35] ), .B(n1098), .Z(\SUMB[4][35] ) );
  EOP U1614 ( .A(\SUMB[3][36] ), .B(n368), .Z(n1098) );
  ND2 U1615 ( .A(\CARRYB[11][3] ), .B(\SUMB[11][4] ), .Z(n1100) );
  ND2 U1616 ( .A(\CARRYB[11][3] ), .B(n346), .Z(n1101) );
  ND2 U1617 ( .A(\SUMB[11][4] ), .B(n346), .Z(n1102) );
  ND2 U1618 ( .A(\CARRYB[6][3] ), .B(\SUMB[6][4] ), .Z(n1104) );
  ND2 U1619 ( .A(\CARRYB[6][3] ), .B(n345), .Z(n1105) );
  ND2 U1620 ( .A(\SUMB[6][4] ), .B(n345), .Z(n1106) );
  EO U1621 ( .A(\SUMB[21][4] ), .B(n1317), .Z(n1107) );
  EOP U1622 ( .A(\CARRYB[21][3] ), .B(n1107), .Z(\SUMB[22][3] ) );
  ND2P U1623 ( .A(\CARRYB[21][3] ), .B(\SUMB[21][4] ), .Z(n1108) );
  ND2P U1624 ( .A(\CARRYB[21][3] ), .B(n1317), .Z(n1109) );
  ND2 U1625 ( .A(\SUMB[21][4] ), .B(n1317), .Z(n1110) );
  ND3P U1626 ( .A(n1108), .B(n1109), .C(n1110), .Z(\CARRYB[22][3] ) );
  IV U1627 ( .A(n1444), .Z(n1442) );
  IV U1628 ( .A(n1444), .Z(n1441) );
  IV U1629 ( .A(n1444), .Z(n1440) );
  EOP U1630 ( .A(\SUMB[4][40] ), .B(n384), .Z(n1113) );
  EOP U1631 ( .A(\CARRYB[4][39] ), .B(n1113), .Z(\SUMB[5][39] ) );
  ND2 U1632 ( .A(\CARRYB[4][39] ), .B(\SUMB[4][40] ), .Z(n1114) );
  ND2 U1633 ( .A(\CARRYB[4][39] ), .B(n384), .Z(n1115) );
  ND2 U1634 ( .A(\SUMB[4][40] ), .B(n384), .Z(n1116) );
  ND2 U1635 ( .A(\SUMB[36][37] ), .B(\ab[37][36] ), .Z(n1120) );
  EOP U1636 ( .A(\SUMB[36][3] ), .B(n309), .Z(n1121) );
  ND2 U1637 ( .A(\SUMB[36][3] ), .B(n309), .Z(n1124) );
  EO3P U1638 ( .A(\CARRYB[26][4] ), .B(n356), .C(\SUMB[26][5] ), .Z(
        \SUMB[27][4] ) );
  ND2 U1639 ( .A(\CARRYB[26][4] ), .B(\SUMB[26][5] ), .Z(n1125) );
  ND2 U1640 ( .A(\CARRYB[26][4] ), .B(n356), .Z(n1126) );
  ND2 U1641 ( .A(\SUMB[26][5] ), .B(n356), .Z(n1127) );
  EO3P U1642 ( .A(\CARRYB[22][30] ), .B(\ab[30][23] ), .C(\SUMB[22][31] ), .Z(
        \SUMB[23][30] ) );
  ND2 U1643 ( .A(\CARRYB[22][30] ), .B(\SUMB[22][31] ), .Z(n1128) );
  ND2 U1644 ( .A(\CARRYB[22][30] ), .B(\ab[30][23] ), .Z(n1129) );
  ND2 U1645 ( .A(\SUMB[22][31] ), .B(\ab[30][23] ), .Z(n1130) );
  ND3 U1646 ( .A(n1128), .B(n1129), .C(n1130), .Z(\CARRYB[23][30] ) );
  EOP U1647 ( .A(\SUMB[44][27] ), .B(\ab[45][26] ), .Z(n1131) );
  ND2 U1648 ( .A(\CARRYB[44][26] ), .B(\SUMB[44][27] ), .Z(n1132) );
  ND2 U1649 ( .A(\CARRYB[44][26] ), .B(\ab[45][26] ), .Z(n1133) );
  ND2 U1650 ( .A(\SUMB[44][27] ), .B(\ab[45][26] ), .Z(n1134) );
  ND2 U1651 ( .A(\CARRYB[34][4] ), .B(\SUMB[34][5] ), .Z(n1136) );
  ND2 U1652 ( .A(\CARRYB[34][4] ), .B(n368), .Z(n1137) );
  ND2 U1653 ( .A(\SUMB[34][5] ), .B(n368), .Z(n1138) );
  EOP U1654 ( .A(\SUMB[17][7] ), .B(n428), .Z(n1139) );
  EOP U1655 ( .A(\CARRYB[17][6] ), .B(n1139), .Z(\SUMB[18][6] ) );
  ND2P U1656 ( .A(\CARRYB[17][6] ), .B(\SUMB[17][7] ), .Z(n1140) );
  ND2 U1657 ( .A(\SUMB[17][7] ), .B(n428), .Z(n1142) );
  AN2P U1658 ( .A(A[41]), .B(\ab[1][1] ), .Z(n1144) );
  EO3P U1659 ( .A(\CARRYB[43][2] ), .B(n308), .C(\SUMB[43][3] ), .Z(
        \SUMB[44][2] ) );
  ND2 U1660 ( .A(\CARRYB[43][2] ), .B(\SUMB[43][3] ), .Z(n1145) );
  ND2 U1661 ( .A(\CARRYB[43][2] ), .B(n308), .Z(n1146) );
  ND2 U1662 ( .A(\SUMB[43][3] ), .B(n308), .Z(n1147) );
  ND3 U1663 ( .A(n1145), .B(n1146), .C(n1147), .Z(\CARRYB[44][2] ) );
  EO U1664 ( .A(\SUMB[17][2] ), .B(n1329), .Z(n1148) );
  ND2P U1665 ( .A(\CARRYB[17][1] ), .B(\SUMB[17][2] ), .Z(n1149) );
  ND2 U1666 ( .A(\SUMB[17][2] ), .B(n1329), .Z(n1151) );
  ND3P U1667 ( .A(n1149), .B(n1150), .C(n1151), .Z(\CARRYB[18][1] ) );
  EO U1668 ( .A(\SUMB[22][2] ), .B(n1420), .Z(n1152) );
  ND2 U1669 ( .A(\SUMB[22][2] ), .B(n1420), .Z(n1155) );
  EOP U1670 ( .A(\CARRYB[23][1] ), .B(n1250), .Z(\SUMB[24][1] ) );
  ND2 U1671 ( .A(\CARRYB[23][1] ), .B(n1360), .Z(n1252) );
  ND2 U1672 ( .A(\CARRYB[23][1] ), .B(\SUMB[23][2] ), .Z(n1251) );
  EO U1673 ( .A(\SUMB[21][8] ), .B(n416), .Z(n1156) );
  ND2 U1674 ( .A(\SUMB[21][8] ), .B(n416), .Z(n1159) );
  ND2 U1675 ( .A(\CARRYB[13][7] ), .B(\SUMB[13][8] ), .Z(n1161) );
  ND2 U1676 ( .A(\CARRYB[13][7] ), .B(n459), .Z(n1162) );
  ND2 U1677 ( .A(\SUMB[13][8] ), .B(n459), .Z(n1163) );
  EOP U1678 ( .A(\SUMB[14][35] ), .B(\ab[34][15] ), .Z(n1164) );
  ND2 U1679 ( .A(\CARRYB[14][34] ), .B(\SUMB[14][35] ), .Z(n1165) );
  ND2 U1680 ( .A(\CARRYB[14][34] ), .B(\ab[34][15] ), .Z(n1166) );
  ND2 U1681 ( .A(\SUMB[14][35] ), .B(\ab[34][15] ), .Z(n1167) );
  ND2 U1682 ( .A(\CARRYB[16][34] ), .B(\SUMB[16][35] ), .Z(n1168) );
  ND2 U1683 ( .A(\CARRYB[16][34] ), .B(\ab[34][17] ), .Z(n1169) );
  ND2 U1684 ( .A(\SUMB[16][35] ), .B(\ab[34][17] ), .Z(n1170) );
  ND3 U1685 ( .A(n1168), .B(n1169), .C(n1170), .Z(\CARRYB[17][34] ) );
  ND2 U1686 ( .A(\CARRYB[8][38] ), .B(\SUMB[8][39] ), .Z(n1172) );
  ND2 U1687 ( .A(\CARRYB[8][38] ), .B(n522), .Z(n1173) );
  ND2 U1688 ( .A(\SUMB[8][39] ), .B(n522), .Z(n1174) );
  ND3P U1689 ( .A(n1172), .B(n1173), .C(n1174), .Z(\CARRYB[9][38] ) );
  EOP U1690 ( .A(\SUMB[44][5] ), .B(n344), .Z(n1175) );
  EOP U1691 ( .A(n1175), .B(\CARRYB[44][4] ), .Z(\SUMB[45][4] ) );
  ND2 U1692 ( .A(\CARRYB[44][4] ), .B(\SUMB[44][5] ), .Z(n1176) );
  ND2 U1693 ( .A(\CARRYB[44][4] ), .B(n344), .Z(n1177) );
  ND2 U1694 ( .A(\SUMB[44][5] ), .B(n344), .Z(n1178) );
  EOP U1695 ( .A(\SUMB[4][6] ), .B(n1445), .Z(n1179) );
  EOP U1696 ( .A(\CARRYB[4][5] ), .B(n1179), .Z(\SUMB[5][5] ) );
  ND2 U1697 ( .A(\CARRYB[4][5] ), .B(\SUMB[4][6] ), .Z(n1180) );
  ND2 U1698 ( .A(\CARRYB[4][5] ), .B(n1445), .Z(n1181) );
  ND2 U1699 ( .A(\SUMB[4][6] ), .B(n1445), .Z(n1182) );
  EO U1700 ( .A(\CARRYB[39][36] ), .B(n1183), .Z(\SUMB[40][36] ) );
  ND2 U1701 ( .A(\CARRYB[39][36] ), .B(\SUMB[39][37] ), .Z(n1184) );
  ND2 U1702 ( .A(\CARRYB[39][36] ), .B(\ab[40][36] ), .Z(n1185) );
  ND3 U1703 ( .A(n1184), .B(n1185), .C(n1186), .Z(\CARRYB[40][36] ) );
  ND2 U1704 ( .A(\CARRYB[10][2] ), .B(\SUMB[10][3] ), .Z(n1188) );
  ND2 U1705 ( .A(\CARRYB[10][2] ), .B(n312), .Z(n1189) );
  EO U1706 ( .A(\SUMB[13][3] ), .B(n342), .Z(n1195) );
  EO U1707 ( .A(\CARRYB[13][2] ), .B(n1195), .Z(\SUMB[14][2] ) );
  EO U1708 ( .A(\SUMB[39][37] ), .B(\ab[40][36] ), .Z(n1183) );
  ND2 U1709 ( .A(\SUMB[39][37] ), .B(\ab[40][36] ), .Z(n1186) );
  ND2 U1710 ( .A(\SUMB[10][3] ), .B(n312), .Z(n1190) );
  EOP U1711 ( .A(\SUMB[19][3] ), .B(n1341), .Z(n1191) );
  EOP U1712 ( .A(\CARRYB[19][2] ), .B(n1191), .Z(\SUMB[20][2] ) );
  ND2 U1713 ( .A(\CARRYB[19][2] ), .B(\SUMB[19][3] ), .Z(n1192) );
  ND2 U1714 ( .A(\CARRYB[19][2] ), .B(n1341), .Z(n1193) );
  ND2 U1715 ( .A(\SUMB[19][3] ), .B(n1341), .Z(n1194) );
  ND3 U1716 ( .A(n1192), .B(n1193), .C(n1194), .Z(\CARRYB[20][2] ) );
  AN2P U1717 ( .A(\ab[20][20] ), .B(A[2]), .Z(n1341) );
  ND2P U1718 ( .A(\CARRYB[13][2] ), .B(\SUMB[13][3] ), .Z(n1196) );
  ND2 U1719 ( .A(\SUMB[13][3] ), .B(n342), .Z(n1198) );
  ND3P U1720 ( .A(n1196), .B(n1197), .C(n1198), .Z(\CARRYB[14][2] ) );
  ND2 U1721 ( .A(\CARRYB[3][35] ), .B(\SUMB[3][36] ), .Z(n1199) );
  ND2 U1722 ( .A(\CARRYB[3][35] ), .B(n368), .Z(n1200) );
  ND2 U1723 ( .A(\SUMB[3][36] ), .B(n368), .Z(n1201) );
  ND3 U1724 ( .A(n1199), .B(n1200), .C(n1201), .Z(\CARRYB[4][35] ) );
  EO U1725 ( .A(\SUMB[37][4] ), .B(n343), .Z(n1202) );
  ND2 U1726 ( .A(\SUMB[37][4] ), .B(n343), .Z(n1205) );
  ND3P U1727 ( .A(n1203), .B(n1204), .C(n1205), .Z(\CARRYB[38][3] ) );
  ND3P U1728 ( .A(n1207), .B(n1208), .C(n1209), .Z(\CARRYB[40][0] ) );
  EO U1729 ( .A(\SUMB[39][1] ), .B(n1352), .Z(n1206) );
  EO U1730 ( .A(\CARRYB[39][0] ), .B(n1206), .Z(\A1[38] ) );
  ND2 U1731 ( .A(\CARRYB[39][0] ), .B(\SUMB[39][1] ), .Z(n1207) );
  ND2 U1732 ( .A(\CARRYB[39][0] ), .B(n1352), .Z(n1208) );
  ND2 U1733 ( .A(\SUMB[39][1] ), .B(n1352), .Z(n1209) );
  AN2P U1734 ( .A(\ab[40][40] ), .B(\B[0] ), .Z(n1352) );
  EO3P U1735 ( .A(n716), .B(\CARRYB[35][0] ), .C(\SUMB[35][1] ), .Z(\A1[34] )
         );
  ND2 U1736 ( .A(n1363), .B(\SUMB[35][1] ), .Z(n1211) );
  ND3P U1737 ( .A(n1210), .B(n1211), .C(n1212), .Z(\CARRYB[36][0] ) );
  EO U1738 ( .A(n1364), .B(\SUMB[36][1] ), .Z(n1213) );
  EO U1739 ( .A(n1213), .B(\CARRYB[36][0] ), .Z(\A1[35] ) );
  ND2P U1740 ( .A(\SUMB[36][1] ), .B(\CARRYB[36][0] ), .Z(n1216) );
  ND3P U1741 ( .A(n1214), .B(n1215), .C(n1216), .Z(\CARRYB[37][0] ) );
  EO U1742 ( .A(\SUMB[27][1] ), .B(n1335), .Z(n1217) );
  EO U1743 ( .A(\CARRYB[27][0] ), .B(n1217), .Z(\A1[26] ) );
  ND2 U1744 ( .A(\CARRYB[27][0] ), .B(\SUMB[27][1] ), .Z(n1218) );
  ND2 U1745 ( .A(\CARRYB[27][0] ), .B(n1335), .Z(n1219) );
  ND2 U1746 ( .A(\SUMB[27][1] ), .B(n1335), .Z(n1220) );
  AN2P U1747 ( .A(A[28]), .B(\B[0] ), .Z(n1335) );
  EO3P U1748 ( .A(n1319), .B(\CARRYB[39][2] ), .C(\SUMB[39][3] ), .Z(
        \SUMB[40][2] ) );
  ND2 U1749 ( .A(n1319), .B(\SUMB[39][3] ), .Z(n1222) );
  ND3P U1750 ( .A(n1221), .B(n1222), .C(n1223), .Z(\CARRYB[40][2] ) );
  EO3 U1751 ( .A(\CARRYB[33][3] ), .B(n305), .C(\SUMB[33][4] ), .Z(
        \SUMB[34][3] ) );
  ND2 U1752 ( .A(\CARRYB[33][3] ), .B(\SUMB[33][4] ), .Z(n1228) );
  ND2 U1753 ( .A(\CARRYB[33][3] ), .B(n305), .Z(n1229) );
  ND2 U1754 ( .A(\SUMB[33][4] ), .B(n305), .Z(n1230) );
  EO U1755 ( .A(\SUMB[44][4] ), .B(n285), .Z(n1242) );
  ND3P U1756 ( .A(n1259), .B(n1260), .C(n1261), .Z(\CARRYB[25][1] ) );
  ND3 U1757 ( .A(n1232), .B(n1233), .C(n1234), .Z(\CARRYB[20][4] ) );
  AN2P U1758 ( .A(A[37]), .B(\B[0] ), .Z(n1364) );
  AN2P U1759 ( .A(A[41]), .B(\B[0] ), .Z(n1373) );
  ND2 U1760 ( .A(\B[0] ), .B(\ab[1][1] ), .Z(n1249) );
  ND2 U1761 ( .A(\CARRYB[19][4] ), .B(\SUMB[19][5] ), .Z(n1232) );
  ND2 U1762 ( .A(\CARRYB[19][4] ), .B(n349), .Z(n1233) );
  ND2 U1763 ( .A(\SUMB[19][5] ), .B(n349), .Z(n1234) );
  EO3 U1764 ( .A(n358), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .Z(\SUMB[3][4] )
         );
  ND2 U1765 ( .A(n358), .B(\CARRYB[2][4] ), .Z(n1235) );
  ND2 U1766 ( .A(n358), .B(\SUMB[2][5] ), .Z(n1236) );
  ND2 U1767 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Z(n1237) );
  ND3 U1768 ( .A(n1235), .B(n1236), .C(n1237), .Z(\CARRYB[3][4] ) );
  EOP U1769 ( .A(n1440), .B(\SUMB[3][5] ), .Z(n1238) );
  EOP U1770 ( .A(n1238), .B(\CARRYB[3][4] ), .Z(\SUMB[4][4] ) );
  ND2 U1771 ( .A(n1440), .B(\CARRYB[3][4] ), .Z(n1240) );
  ND2P U1772 ( .A(\SUMB[3][5] ), .B(\CARRYB[3][4] ), .Z(n1241) );
  ND2 U1773 ( .A(\CARRYB[44][3] ), .B(\SUMB[44][4] ), .Z(n1243) );
  ND2 U1774 ( .A(\CARRYB[44][3] ), .B(n285), .Z(n1244) );
  ND2 U1775 ( .A(\SUMB[44][4] ), .B(n285), .Z(n1245) );
  EO3 U1776 ( .A(\CARRYB[17][4] ), .B(n350), .C(\SUMB[17][5] ), .Z(
        \SUMB[18][4] ) );
  ND2 U1777 ( .A(\CARRYB[17][4] ), .B(\SUMB[17][5] ), .Z(n1246) );
  ND2 U1778 ( .A(\CARRYB[17][4] ), .B(n350), .Z(n1247) );
  ND2 U1779 ( .A(\SUMB[17][5] ), .B(n350), .Z(n1248) );
  ND3 U1780 ( .A(n1246), .B(n1247), .C(n1248), .Z(\CARRYB[18][4] ) );
  EOP U1781 ( .A(\CARRYB[47][17] ), .B(\SUMB[47][18] ), .Z(\A1[63] ) );
  ND2 U1782 ( .A(\CARRYB[24][1] ), .B(n1413), .Z(n1260) );
  EOP U1783 ( .A(\SUMB[23][2] ), .B(n1360), .Z(n1250) );
  ND2 U1784 ( .A(\SUMB[23][2] ), .B(n1360), .Z(n1253) );
  ND3P U1785 ( .A(n1251), .B(n1252), .C(n1253), .Z(\CARRYB[24][1] ) );
  ND2 U1786 ( .A(\CARRYB[24][1] ), .B(\SUMB[24][2] ), .Z(n1259) );
  EO U1787 ( .A(\CARRYB[47][33] ), .B(\SUMB[47][34] ), .Z(\A1[79] ) );
  EO U1788 ( .A(\CARRYB[47][1] ), .B(\SUMB[47][2] ), .Z(\A1[47] ) );
  AN2P U1789 ( .A(A[38]), .B(A[2]), .Z(n1312) );
  AN2P U1790 ( .A(A[45]), .B(A[2]), .Z(n1314) );
  AN2P U1791 ( .A(A[21]), .B(A[2]), .Z(n1305) );
  AN2P U1792 ( .A(A[43]), .B(A[3]), .Z(n1320) );
  AN2P U1793 ( .A(\ab[16][16] ), .B(n1436), .Z(n1321) );
  AN2 U1794 ( .A(n1465), .B(n1441), .Z(n1278) );
  AN2P U1795 ( .A(n1470), .B(n1441), .Z(n1277) );
  EO U1796 ( .A(n1392), .B(n1383), .Z(\SUMB[1][6] ) );
  EO U1797 ( .A(n1375), .B(n1344), .Z(\SUMB[1][19] ) );
  EO U1798 ( .A(\CARRYB[42][1] ), .B(n1266), .Z(\SUMB[43][1] ) );
  ND2 U1799 ( .A(\CARRYB[42][1] ), .B(\SUMB[42][2] ), .Z(n1267) );
  ND2 U1800 ( .A(\CARRYB[42][1] ), .B(n1422), .Z(n1268) );
  ND2 U1801 ( .A(\CARRYB[34][1] ), .B(\SUMB[34][2] ), .Z(n1263) );
  ND2 U1802 ( .A(\CARRYB[34][1] ), .B(n743), .Z(n1264) );
  EO U1803 ( .A(\CARRYB[38][1] ), .B(n1254), .Z(\SUMB[39][1] ) );
  ND2 U1804 ( .A(\CARRYB[38][1] ), .B(\SUMB[38][2] ), .Z(n1255) );
  ND2 U1805 ( .A(\CARRYB[38][1] ), .B(n1347), .Z(n1256) );
  AN2P U1806 ( .A(\ab[6][6] ), .B(\B[0] ), .Z(n1387) );
  AN2P U1807 ( .A(A[4]), .B(\B[0] ), .Z(n1388) );
  IVP U1808 ( .A(\ab[5][5] ), .Z(n1448) );
  AN2P U1809 ( .A(A[39]), .B(\B[0] ), .Z(n1365) );
  AN2P U1810 ( .A(A[35]), .B(\B[0] ), .Z(n1362) );
  AN2P U1811 ( .A(\ab[31][31] ), .B(A[2]), .Z(n1340) );
  AN2P U1812 ( .A(A[29]), .B(\B[0] ), .Z(n1366) );
  AN2P U1813 ( .A(\ab[18][18] ), .B(A[2]), .Z(n1339) );
  AN2P U1814 ( .A(\ab[18][18] ), .B(n1436), .Z(n1391) );
  EO U1815 ( .A(\SUMB[38][2] ), .B(n1347), .Z(n1254) );
  ND2 U1816 ( .A(\SUMB[38][2] ), .B(n1347), .Z(n1257) );
  EO U1817 ( .A(\SUMB[24][2] ), .B(n1413), .Z(n1258) );
  ND2 U1818 ( .A(\SUMB[24][2] ), .B(n1413), .Z(n1261) );
  EO U1819 ( .A(\SUMB[34][2] ), .B(n743), .Z(n1262) );
  ND2 U1820 ( .A(\SUMB[34][2] ), .B(n743), .Z(n1265) );
  ND2 U1821 ( .A(\SUMB[42][2] ), .B(n1422), .Z(n1269) );
  EOP U1822 ( .A(\CARRYB[47][24] ), .B(\SUMB[47][25] ), .Z(\A1[70] ) );
  EOP U1823 ( .A(\CARRYB[47][27] ), .B(\SUMB[47][28] ), .Z(\A1[73] ) );
  EOP U1824 ( .A(\CARRYB[47][15] ), .B(\SUMB[47][16] ), .Z(\A1[61] ) );
  EOP U1825 ( .A(\CARRYB[47][35] ), .B(\SUMB[47][36] ), .Z(\A1[81] ) );
  EOP U1826 ( .A(\CARRYB[47][21] ), .B(\SUMB[47][22] ), .Z(\A1[67] ) );
  EOP U1827 ( .A(\CARRYB[47][10] ), .B(\SUMB[47][11] ), .Z(\A1[56] ) );
  ND2 U1828 ( .A(\CARRYB[28][5] ), .B(\SUMB[28][6] ), .Z(n1295) );
  ND2 U1829 ( .A(\CARRYB[28][5] ), .B(n1276), .Z(n1296) );
  AN2 U1830 ( .A(A[39]), .B(A[2]), .Z(n1313) );
  AN2P U1831 ( .A(n1491), .B(n1442), .Z(n1271) );
  AN2 U1832 ( .A(n1479), .B(n1441), .Z(n1272) );
  AN2P U1833 ( .A(A[38]), .B(n1447), .Z(n1273) );
  AN2P U1834 ( .A(n1505), .B(n1442), .Z(n1274) );
  AN2P U1835 ( .A(n1479), .B(n1446), .Z(n1275) );
  AN2P U1836 ( .A(n1491), .B(n1447), .Z(n1276) );
  AN2P U1837 ( .A(A[29]), .B(n1451), .Z(n1279) );
  AN2P U1838 ( .A(A[38]), .B(n1451), .Z(n1280) );
  AN2P U1839 ( .A(n1505), .B(n1447), .Z(n1281) );
  AN2P U1840 ( .A(n1479), .B(n1450), .Z(n1282) );
  AN2P U1841 ( .A(n1470), .B(n1446), .Z(n1283) );
  AN2P U1842 ( .A(n1465), .B(n1446), .Z(n1284) );
  AN2P U1843 ( .A(n1479), .B(n1454), .Z(n1285) );
  AN2P U1844 ( .A(n1505), .B(n1451), .Z(n1286) );
  AN2P U1845 ( .A(A[29]), .B(n1455), .Z(n1287) );
  AN2 U1846 ( .A(A[38]), .B(n1455), .Z(n1288) );
  AN2P U1847 ( .A(n1525), .B(n1453), .Z(\ab[7][46] ) );
  AN2P U1848 ( .A(n1470), .B(n1450), .Z(n1289) );
  AN2P U1849 ( .A(A[29]), .B(A[8]), .Z(n1290) );
  AN2P U1850 ( .A(n1479), .B(A[8]), .Z(n1291) );
  AN2P U1851 ( .A(n1465), .B(n1450), .Z(n1292) );
  AN2P U1852 ( .A(A[38]), .B(A[8]), .Z(n1293) );
  EOP U1853 ( .A(n1399), .B(n1360), .Z(\SUMB[1][24] ) );
  AN2 U1854 ( .A(n1369), .B(n1365), .Z(\CARRYB[1][38] ) );
  IV U1855 ( .A(n1439), .Z(n1437) );
  AN2 U1856 ( .A(n1323), .B(n1326), .Z(\CARRYB[1][32] ) );
  IV U1857 ( .A(n1439), .Z(n1436) );
  AN2 U1858 ( .A(n1422), .B(n306), .Z(\CARRYB[1][43] ) );
  IV U1859 ( .A(n1527), .Z(n1525) );
  IVP U1860 ( .A(n1448), .Z(n1447) );
  IVP U1861 ( .A(n1448), .Z(n1446) );
  AN2 U1862 ( .A(A[5]), .B(\B[0] ), .Z(n1389) );
  AN2 U1863 ( .A(\ab[2][2] ), .B(\B[0] ), .Z(n1390) );
  AN2 U1864 ( .A(\ab[19][19] ), .B(\B[0] ), .Z(n1334) );
  AN2 U1865 ( .A(A[23]), .B(\B[0] ), .Z(n1338) );
  AN2 U1866 ( .A(\ab[20][20] ), .B(\B[0] ), .Z(n1375) );
  AN2 U1867 ( .A(A[10]), .B(\B[0] ), .Z(n1385) );
  IVP U1868 ( .A(\ab[17][17] ), .Z(n1467) );
  ND2 U1869 ( .A(\SUMB[28][6] ), .B(n1276), .Z(n1297) );
  EO U1870 ( .A(\CARRYB[47][44] ), .B(\SUMB[47][45] ), .Z(\A1[90] ) );
  EO U1871 ( .A(\CARRYB[47][39] ), .B(\SUMB[47][40] ), .Z(\A1[85] ) );
  EO U1872 ( .A(\CARRYB[47][40] ), .B(\SUMB[47][41] ), .Z(\A1[86] ) );
  AN2P U1873 ( .A(\ab[16][16] ), .B(A[2]), .Z(n1299) );
  AN2P U1874 ( .A(\ab[24][24] ), .B(A[2]), .Z(n1300) );
  AN2P U1875 ( .A(A[22]), .B(A[2]), .Z(n1301) );
  AN2P U1876 ( .A(A[29]), .B(A[2]), .Z(n1303) );
  AN2P U1877 ( .A(A[15]), .B(A[2]), .Z(n1304) );
  AN2P U1878 ( .A(A[33]), .B(A[2]), .Z(n1306) );
  AN2P U1879 ( .A(\ab[34][34] ), .B(A[2]), .Z(n1307) );
  AN2P U1880 ( .A(A[46]), .B(A[2]), .Z(n1308) );
  AN2P U1881 ( .A(A[28]), .B(A[2]), .Z(n1309) );
  AN2P U1882 ( .A(A[27]), .B(A[2]), .Z(n1310) );
  AN2P U1883 ( .A(A[41]), .B(A[2]), .Z(n1311) );
  AN2P U1884 ( .A(A[32]), .B(A[2]), .Z(n1315) );
  AN2P U1885 ( .A(A[35]), .B(n1433), .Z(n1316) );
  AN2P U1886 ( .A(n1476), .B(n1436), .Z(n1317) );
  AN2P U1887 ( .A(A[15]), .B(n1436), .Z(n1318) );
  AN2P U1888 ( .A(A[40]), .B(A[2]), .Z(n1319) );
  EO U1889 ( .A(\CARRYB[47][0] ), .B(\SUMB[47][1] ), .Z(\A1[46] ) );
  EO U1890 ( .A(\CARRYB[47][46] ), .B(A[47]), .Z(\A1[92] ) );
  EO U1891 ( .A(n1334), .B(n1329), .Z(\SUMB[1][18] ) );
  EO U1892 ( .A(n1326), .B(n1323), .Z(\SUMB[1][32] ) );
  EO U1893 ( .A(n1335), .B(n1330), .Z(\SUMB[1][27] ) );
  EO U1894 ( .A(n310), .B(n268), .Z(\SUMB[1][21] ) );
  EO U1895 ( .A(n1429), .B(n1427), .Z(\SUMB[1][16] ) );
  EO U1896 ( .A(n1365), .B(n1369), .Z(\SUMB[1][38] ) );
  EO U1897 ( .A(n1373), .B(n1348), .Z(\SUMB[1][40] ) );
  EO U1898 ( .A(n1395), .B(n267), .Z(\SUMB[1][15] ) );
  EO U1899 ( .A(n1336), .B(n304), .Z(\SUMB[1][45] ) );
  EO U1900 ( .A(n1417), .B(n1333), .Z(\SUMB[1][42] ) );
  EO U1901 ( .A(n1431), .B(n1376), .Z(\SUMB[1][14] ) );
  IVP U1902 ( .A(n1467), .Z(n1466) );
  IVP U1903 ( .A(n1471), .Z(n1469) );
  EO U1904 ( .A(n1352), .B(n1347), .Z(\SUMB[1][39] ) );
  EO U1905 ( .A(n1384), .B(n1382), .Z(\SUMB[1][11] ) );
  IVP U1906 ( .A(n1471), .Z(n1468) );
  IV U1907 ( .A(n1481), .Z(n1480) );
  IV U1908 ( .A(n1492), .Z(n1491) );
  IVP U1909 ( .A(n1467), .Z(n1464) );
  EO U1910 ( .A(n1368), .B(n1353), .Z(\SUMB[1][8] ) );
  EO U1911 ( .A(n1389), .B(n1532), .Z(\SUMB[1][4] ) );
  EO U1912 ( .A(n1387), .B(n1377), .Z(\SUMB[1][5] ) );
  EO U1913 ( .A(n1388), .B(n1528), .Z(\SUMB[1][3] ) );
  IV U1914 ( .A(n1439), .Z(n1435) );
  IVP U1915 ( .A(n1452), .Z(n1449) );
  IVP U1916 ( .A(n1452), .Z(n1450) );
  IVP U1917 ( .A(n1452), .Z(n1451) );
  IVP U1918 ( .A(n1456), .Z(n1453) );
  IVP U1919 ( .A(n1456), .Z(n1454) );
  IVP U1920 ( .A(n1456), .Z(n1455) );
  IVDA U1921 ( .A(n1524), .Y(n1523) );
  IVDA U1922 ( .A(n1522), .Y(n1520) );
  IVDA U1923 ( .A(n1513), .Y(n1510) );
  NR2 U1924 ( .A(n1472), .B(n1458), .Z(n1322) );
  IVDA U1925 ( .A(n1463), .Y(n1462) );
  IVDA U1926 ( .A(n1477), .Y(n1476) );
  IVDA U1927 ( .A(n1490), .Y(n1489) );
  IVP U1928 ( .A(n1497), .Z(n1495) );
  IVDA U1929 ( .A(n1460), .Y(n1459) );
  IVP U1930 ( .A(n1519), .Z(n1517) );
  IVDA U1931 ( .A(n1513), .Y(n1512) );
  IVDA U1932 ( .A(n1477), .Y(n1474) );
  IVDA U1933 ( .A(n1477), .Y(n1475) );
  IVDA U1934 ( .A(n1490), .Y(n1488) );
  IVP U1935 ( .A(n1497), .Z(n1494) );
  IVDA U1936 ( .A(n1522), .Y(n1521) );
  IVP U1937 ( .A(n1519), .Z(n1516) );
  IVDA U1938 ( .A(n1513), .Y(n1511) );
  IVDA U1939 ( .A(n1527), .Y(n1526) );
  IVDA U1940 ( .A(n1490), .Y(n1487) );
  IVP U1941 ( .A(n1497), .Z(n1493) );
  AN2P U1942 ( .A(A[32]), .B(\ab[1][1] ), .Z(n1323) );
  AN2P U1943 ( .A(\ab[29][29] ), .B(\ab[1][1] ), .Z(n1324) );
  AN2P U1944 ( .A(\B[0] ), .B(\ab[47][47] ), .Z(n1327) );
  AN2P U1945 ( .A(\ab[42][42] ), .B(A[2]), .Z(n1328) );
  AN2P U1946 ( .A(\ab[18][18] ), .B(\ab[1][1] ), .Z(n1329) );
  AN2P U1947 ( .A(A[27]), .B(\ab[1][1] ), .Z(n1330) );
  AN2P U1948 ( .A(A[28]), .B(\ab[1][1] ), .Z(n1331) );
  AN2P U1949 ( .A(\ab[46][46] ), .B(\ab[1][1] ), .Z(n1332) );
  AN2P U1950 ( .A(\ab[42][42] ), .B(\ab[1][1] ), .Z(n1333) );
  NR2 U1951 ( .A(n1522), .B(n872), .Z(n1417) );
  AN2P U1952 ( .A(A[46]), .B(\B[0] ), .Z(n1336) );
  AN2P U1953 ( .A(\ab[1][1] ), .B(A[47]), .Z(n1343) );
  AN2P U1954 ( .A(A[19]), .B(\ab[1][1] ), .Z(n1344) );
  AN2P U1955 ( .A(\ab[37][37] ), .B(\ab[1][1] ), .Z(n1345) );
  AN2P U1956 ( .A(\ab[10][10] ), .B(\ab[1][1] ), .Z(n1346) );
  AN2P U1957 ( .A(\ab[39][39] ), .B(\ab[1][1] ), .Z(n1347) );
  AN2P U1958 ( .A(A[40]), .B(\ab[1][1] ), .Z(n1348) );
  AN2P U1959 ( .A(\ab[14][14] ), .B(\B[0] ), .Z(n1351) );
  AN2P U1960 ( .A(A[8]), .B(\ab[1][1] ), .Z(n1353) );
  AN2P U1961 ( .A(\ab[12][12] ), .B(\ab[1][1] ), .Z(n1354) );
  AN2P U1962 ( .A(A[35]), .B(\ab[1][1] ), .Z(n1355) );
  AN2P U1963 ( .A(\ab[44][44] ), .B(\ab[1][1] ), .Z(n1357) );
  AN2P U1964 ( .A(\ab[13][13] ), .B(\B[0] ), .Z(n1358) );
  AN2P U1965 ( .A(\ab[34][34] ), .B(\ab[1][1] ), .Z(n1359) );
  AN2P U1966 ( .A(A[24]), .B(\ab[1][1] ), .Z(n1360) );
  NR2 U1967 ( .A(n1524), .B(n872), .Z(n1415) );
  AN2P U1968 ( .A(\ab[31][31] ), .B(\ab[1][1] ), .Z(n1361) );
  AN2P U1969 ( .A(A[9]), .B(\B[0] ), .Z(n1368) );
  AN2P U1970 ( .A(A[38]), .B(\ab[1][1] ), .Z(n1369) );
  AN2P U1971 ( .A(A[13]), .B(\ab[1][1] ), .Z(n1370) );
  AN2P U1972 ( .A(\ab[11][11] ), .B(\B[0] ), .Z(n1371) );
  AN2P U1973 ( .A(A[33]), .B(\ab[1][1] ), .Z(n1372) );
  AN2P U1974 ( .A(A[14]), .B(\ab[1][1] ), .Z(n1376) );
  AN2P U1975 ( .A(\ab[5][5] ), .B(\ab[1][1] ), .Z(n1377) );
  AN2P U1976 ( .A(\ab[9][9] ), .B(\ab[1][1] ), .Z(n1378) );
  AN2P U1977 ( .A(\ab[20][20] ), .B(n1436), .Z(n1379) );
  AN2P U1978 ( .A(\ab[42][42] ), .B(A[3]), .Z(n1380) );
  AN2P U1979 ( .A(\ab[7][7] ), .B(\ab[1][1] ), .Z(n1381) );
  AN2P U1980 ( .A(A[11]), .B(\ab[1][1] ), .Z(n1382) );
  AN2P U1981 ( .A(\ab[6][6] ), .B(\ab[1][1] ), .Z(n1383) );
  AN2P U1982 ( .A(A[12]), .B(\B[0] ), .Z(n1384) );
  AN2P U1983 ( .A(\ab[7][7] ), .B(\B[0] ), .Z(n1392) );
  EO U1984 ( .A(n1530), .B(n1534), .Z(\SUMB[1][2] ) );
  IVP U1985 ( .A(\ab[42][42] ), .Z(n1519) );
  IVP U1986 ( .A(\ab[31][31] ), .Z(n1497) );
  AN2P U1987 ( .A(\CARRYB[47][3] ), .B(\SUMB[47][4] ), .Z(\A2[50] ) );
  EOP U1988 ( .A(\CARRYB[47][3] ), .B(\SUMB[47][4] ), .Z(\A1[49] ) );
  AN2P U1989 ( .A(\CARRYB[47][13] ), .B(\SUMB[47][14] ), .Z(\A2[60] ) );
  EOP U1990 ( .A(\SUMB[47][14] ), .B(\CARRYB[47][13] ), .Z(\A1[59] ) );
  AN2P U1991 ( .A(\CARRYB[47][14] ), .B(\SUMB[47][15] ), .Z(\A2[61] ) );
  EOP U1992 ( .A(\CARRYB[47][14] ), .B(\SUMB[47][15] ), .Z(\A1[60] ) );
  AN2P U1993 ( .A(\CARRYB[47][18] ), .B(\SUMB[47][19] ), .Z(\A2[65] ) );
  AN2P U1994 ( .A(\CARRYB[47][19] ), .B(\SUMB[47][20] ), .Z(\A2[66] ) );
  EOP U1995 ( .A(\CARRYB[47][19] ), .B(\SUMB[47][20] ), .Z(\A1[65] ) );
  AN2P U1996 ( .A(\CARRYB[47][20] ), .B(\SUMB[47][21] ), .Z(\A2[67] ) );
  AN2P U1997 ( .A(\CARRYB[47][29] ), .B(\SUMB[47][30] ), .Z(\A2[76] ) );
  AN2P U1998 ( .A(\CARRYB[47][31] ), .B(\SUMB[47][32] ), .Z(\A2[78] ) );
  EOP U1999 ( .A(\CARRYB[47][31] ), .B(\SUMB[47][32] ), .Z(\A1[77] ) );
  AN2P U2000 ( .A(\CARRYB[47][35] ), .B(\SUMB[47][36] ), .Z(\A2[82] ) );
  AN2P U2001 ( .A(\CARRYB[47][36] ), .B(\SUMB[47][37] ), .Z(\A2[83] ) );
  EOP U2002 ( .A(\CARRYB[47][36] ), .B(\SUMB[47][37] ), .Z(\A1[82] ) );
  AN2P U2003 ( .A(\CARRYB[47][37] ), .B(\SUMB[47][38] ), .Z(\A2[84] ) );
  EOP U2004 ( .A(\CARRYB[47][37] ), .B(\SUMB[47][38] ), .Z(\A1[83] ) );
  AN2P U2005 ( .A(\CARRYB[47][38] ), .B(\SUMB[47][39] ), .Z(\A2[85] ) );
  EOP U2006 ( .A(\CARRYB[47][38] ), .B(\SUMB[47][39] ), .Z(\A1[84] ) );
  AN2P U2007 ( .A(\CARRYB[47][42] ), .B(\SUMB[47][43] ), .Z(\A2[89] ) );
  AN2P U2008 ( .A(\CARRYB[47][43] ), .B(\SUMB[47][44] ), .Z(\A2[90] ) );
  EOP U2009 ( .A(\CARRYB[47][43] ), .B(\SUMB[47][44] ), .Z(\A1[89] ) );
  AN2P U2010 ( .A(\CARRYB[47][44] ), .B(\SUMB[47][45] ), .Z(\A2[91] ) );
  AN2P U2011 ( .A(\CARRYB[47][45] ), .B(\CARRYB[46][46] ), .Z(\A2[92] ) );
  EOP U2012 ( .A(\CARRYB[47][45] ), .B(\CARRYB[46][46] ), .Z(\A1[91] ) );
  AN2P U2013 ( .A(n1528), .B(n1388), .Z(\CARRYB[1][3] ) );
  AN2P U2014 ( .A(n1532), .B(n1389), .Z(\CARRYB[1][4] ) );
  AN2P U2015 ( .A(n1377), .B(n1387), .Z(\CARRYB[1][5] ) );
  AN2P U2016 ( .A(n1383), .B(n1392), .Z(\CARRYB[1][6] ) );
  AN2P U2017 ( .A(n1381), .B(n1386), .Z(\CARRYB[1][7] ) );
  AN2P U2018 ( .A(n1378), .B(n1385), .Z(\CARRYB[1][9] ) );
  AN2P U2019 ( .A(n1382), .B(n1384), .Z(\CARRYB[1][11] ) );
  AN2P U2020 ( .A(n1354), .B(n1358), .Z(\CARRYB[1][12] ) );
  AN2P U2021 ( .A(n1426), .B(n1428), .Z(\CARRYB[1][17] ) );
  EOP U2022 ( .A(n1428), .B(n1426), .Z(\SUMB[1][17] ) );
  EOP U2023 ( .A(n1337), .B(n1412), .Z(\SUMB[1][25] ) );
  AN2P U2024 ( .A(n1403), .B(n1364), .Z(\CARRYB[1][36] ) );
  EOP U2025 ( .A(n1364), .B(n1403), .Z(\SUMB[1][36] ) );
  AN2P U2026 ( .A(\CARRYB[47][34] ), .B(\SUMB[47][35] ), .Z(\A2[81] ) );
  AN2P U2027 ( .A(\CARRYB[47][12] ), .B(\SUMB[47][13] ), .Z(\A2[59] ) );
  EOP U2028 ( .A(\CARRYB[47][12] ), .B(\SUMB[47][13] ), .Z(\A1[58] ) );
  AN2P U2029 ( .A(\CARRYB[47][10] ), .B(\SUMB[47][11] ), .Z(\A2[57] ) );
  AN2P U2030 ( .A(\CARRYB[47][8] ), .B(\SUMB[47][9] ), .Z(\A2[55] ) );
  EOP U2031 ( .A(\CARRYB[47][8] ), .B(\SUMB[47][9] ), .Z(\A1[54] ) );
  AN2P U2032 ( .A(\CARRYB[47][27] ), .B(\SUMB[47][28] ), .Z(\A2[74] ) );
  AN2P U2033 ( .A(\CARRYB[47][22] ), .B(\SUMB[47][23] ), .Z(\A2[69] ) );
  EOP U2034 ( .A(\CARRYB[47][22] ), .B(\SUMB[47][23] ), .Z(\A1[68] ) );
  AN2P U2035 ( .A(\CARRYB[47][30] ), .B(\SUMB[47][31] ), .Z(\A2[77] ) );
  EOP U2036 ( .A(\CARRYB[47][30] ), .B(\SUMB[47][31] ), .Z(\A1[76] ) );
  AN2P U2037 ( .A(\CARRYB[47][39] ), .B(\SUMB[47][40] ), .Z(\A2[86] ) );
  AN2P U2038 ( .A(n1353), .B(n1368), .Z(\CARRYB[1][8] ) );
  AN2P U2039 ( .A(\CARRYB[47][46] ), .B(A[47]), .Z(\A2[93] ) );
  AN2P U2040 ( .A(\CARRYB[47][23] ), .B(\SUMB[47][24] ), .Z(\A2[70] ) );
  EOP U2041 ( .A(\CARRYB[47][23] ), .B(\SUMB[47][24] ), .Z(\A1[69] ) );
  AN2P U2042 ( .A(\CARRYB[47][17] ), .B(\SUMB[47][18] ), .Z(\A2[64] ) );
  AN2P U2043 ( .A(\CARRYB[47][41] ), .B(\SUMB[47][42] ), .Z(\A2[88] ) );
  AN2P U2044 ( .A(n1346), .B(n1371), .Z(\CARRYB[1][10] ) );
  AN2P U2045 ( .A(\CARRYB[47][6] ), .B(\SUMB[47][7] ), .Z(\A2[53] ) );
  AN2P U2046 ( .A(\CARRYB[47][24] ), .B(\SUMB[47][25] ), .Z(\A2[71] ) );
  AN2P U2047 ( .A(\CARRYB[47][28] ), .B(\SUMB[47][29] ), .Z(\A2[75] ) );
  AN2P U2048 ( .A(\CARRYB[47][16] ), .B(\SUMB[47][17] ), .Z(\A2[63] ) );
  EOP U2049 ( .A(\CARRYB[47][16] ), .B(\SUMB[47][17] ), .Z(\A1[62] ) );
  AN2P U2050 ( .A(\CARRYB[47][5] ), .B(\SUMB[47][6] ), .Z(\A2[52] ) );
  EOP U2051 ( .A(\CARRYB[47][5] ), .B(\SUMB[47][6] ), .Z(\A1[51] ) );
  AN2P U2052 ( .A(\CARRYB[47][2] ), .B(\SUMB[47][3] ), .Z(\A2[49] ) );
  AN2P U2053 ( .A(\CARRYB[47][4] ), .B(\SUMB[47][5] ), .Z(\A2[51] ) );
  EOP U2054 ( .A(\CARRYB[47][4] ), .B(\SUMB[47][5] ), .Z(\A1[50] ) );
  AN2P U2055 ( .A(\CARRYB[47][11] ), .B(\SUMB[47][12] ), .Z(\A2[58] ) );
  EOP U2056 ( .A(\CARRYB[47][11] ), .B(\SUMB[47][12] ), .Z(\A1[57] ) );
  AN2P U2057 ( .A(\CARRYB[47][9] ), .B(\SUMB[47][10] ), .Z(\A2[56] ) );
  AN2P U2058 ( .A(\CARRYB[47][15] ), .B(\SUMB[47][16] ), .Z(\A2[62] ) );
  AN2P U2059 ( .A(\CARRYB[47][7] ), .B(\SUMB[47][8] ), .Z(\A2[54] ) );
  AN2P U2060 ( .A(n1414), .B(n1398), .Z(\CARRYB[1][20] ) );
  AN2P U2061 ( .A(n1370), .B(n1351), .Z(\CARRYB[1][13] ) );
  AN2P U2062 ( .A(\CARRYB[47][21] ), .B(\SUMB[47][22] ), .Z(\A2[68] ) );
  AN2P U2063 ( .A(\CARRYB[47][40] ), .B(\SUMB[47][41] ), .Z(\A2[87] ) );
  AN2P U2064 ( .A(\CARRYB[47][25] ), .B(\SUMB[47][26] ), .Z(\A2[72] ) );
  EOP U2065 ( .A(\CARRYB[47][25] ), .B(\SUMB[47][26] ), .Z(\A1[71] ) );
  AN2P U2066 ( .A(n1329), .B(n1334), .Z(\CARRYB[1][18] ) );
  AN2P U2067 ( .A(n1405), .B(n1342), .Z(\CARRYB[1][30] ) );
  AN2P U2068 ( .A(n1359), .B(n1362), .Z(\CARRYB[1][34] ) );
  AN2P U2069 ( .A(n1427), .B(n1429), .Z(\CARRYB[1][16] ) );
  AN2P U2070 ( .A(\CARRYB[47][26] ), .B(\SUMB[47][27] ), .Z(\A2[73] ) );
  EOP U2071 ( .A(\CARRYB[47][26] ), .B(\SUMB[47][27] ), .Z(\A1[72] ) );
  AN2P U2072 ( .A(n1355), .B(n1363), .Z(\CARRYB[1][35] ) );
  AN2P U2073 ( .A(n1348), .B(n1373), .Z(\CARRYB[1][40] ) );
  AN2P U2074 ( .A(n1344), .B(n1375), .Z(\CARRYB[1][19] ) );
  AN2P U2075 ( .A(n1331), .B(n1366), .Z(\CARRYB[1][28] ) );
  AN2P U2076 ( .A(n1333), .B(n1417), .Z(\CARRYB[1][42] ) );
  AN2P U2077 ( .A(n1330), .B(n1335), .Z(\CARRYB[1][27] ) );
  AN2P U2078 ( .A(\CARRYB[47][32] ), .B(\SUMB[47][33] ), .Z(\A2[79] ) );
  EOP U2079 ( .A(\CARRYB[47][32] ), .B(\SUMB[47][33] ), .Z(\A1[78] ) );
  AN2P U2080 ( .A(n1419), .B(n1325), .Z(\CARRYB[1][23] ) );
  IVDA U2081 ( .A(n1503), .Y(n1501) );
  IVDA U2082 ( .A(n1503), .Y(n1500) );
  IVDA U2083 ( .A(n1486), .Y(n1485) );
  IVDA U2084 ( .A(n1486), .Y(n1484) );
  IVDA U2085 ( .A(n1486), .Y(n1483) );
  NR2P U2086 ( .A(n1482), .B(n1411), .Z(n1412) );
  AN2P U2087 ( .A(\ab[43][43] ), .B(A[1]), .Z(n1422) );
  AN2P U2088 ( .A(A[22]), .B(\ab[1][1] ), .Z(n1393) );
  NR2P U2089 ( .A(n720), .B(n1397), .Z(n1396) );
  B4IP U2090 ( .A(\B[0] ), .Z(n1397) );
  NR2P U2091 ( .A(n736), .B(n1397), .Z(n1399) );
  NR2P U2092 ( .A(n1472), .B(n1400), .Z(n1414) );
  AN2P U2093 ( .A(A[16]), .B(A[1]), .Z(n1427) );
  IVP U2094 ( .A(n1497), .Z(n1496) );
  AN2P U2095 ( .A(\ab[36][36] ), .B(\ab[1][1] ), .Z(n1404) );
  NR2P U2096 ( .A(n719), .B(n807), .Z(n1405) );
  AN2P U2097 ( .A(A[26]), .B(\ab[1][1] ), .Z(n1408) );
  AN2P U2098 ( .A(\ab[26][26] ), .B(\ab[1][1] ), .Z(n1409) );
  AN2 U2099 ( .A(A[25]), .B(\ab[1][1] ), .Z(n1413) );
  IVP U2100 ( .A(n1519), .Z(n1518) );
  AN2P U2101 ( .A(A[45]), .B(\B[0] ), .Z(n1416) );
  AN2P U2102 ( .A(n1521), .B(\B[0] ), .Z(n1418) );
  AN2 U2103 ( .A(A[23]), .B(\ab[1][1] ), .Z(n1420) );
  IVDA U2104 ( .A(n1519), .Y(n1515) );
  IVA U2105 ( .A(n1471), .Z(n1470) );
  IVA U2106 ( .A(n1481), .Z(n1479) );
  IVA U2107 ( .A(n1467), .Z(n1465) );
  AN2 U2108 ( .A(\ab[17][17] ), .B(\ab[1][1] ), .Z(n1426) );
  AN2 U2109 ( .A(n1465), .B(\ab[1][1] ), .Z(n1430) );
  AN2 U2110 ( .A(\ab[18][18] ), .B(\B[0] ), .Z(n1428) );
  AN2P U2111 ( .A(A[17]), .B(\B[0] ), .Z(n1429) );
  AN2 U2112 ( .A(A[15]), .B(\B[0] ), .Z(n1431) );
  AN2 U2113 ( .A(n1461), .B(\B[0] ), .Z(n1432) );
  B4IP U2114 ( .A(\ab[25][25] ), .Z(n1482) );
  IVA U2115 ( .A(n1439), .Z(n1438) );
  IV U2116 ( .A(n1444), .Z(n1443) );
  AN2P U2117 ( .A(n1443), .B(\ab[1][1] ), .Z(n1532) );
  AN2P U2118 ( .A(n1438), .B(\ab[1][1] ), .Z(n1528) );
  AN2P U2119 ( .A(n1438), .B(\B[0] ), .Z(n1530) );
  AN2P U2120 ( .A(n1433), .B(\ab[1][1] ), .Z(n1534) );
  AN2P U2121 ( .A(A[2]), .B(\ab[1][1] ), .Z(n1535) );
  AN2P U2122 ( .A(\ab[1][1] ), .B(\B[0] ), .Z(\ab[1][0] ) );
  AN2P U2123 ( .A(n1435), .B(\ab[1][1] ), .Z(n1529) );
  AN2P U2124 ( .A(n1435), .B(\B[0] ), .Z(n1531) );
  AN2P U2125 ( .A(n1440), .B(\ab[1][1] ), .Z(n1533) );
  AN2 U2127 ( .A(A[47]), .B(A[9]), .Z(\ab[9][47] ) );
  AN2 U2128 ( .A(A[47]), .B(A[8]), .Z(\ab[8][47] ) );
  AN2 U2129 ( .A(A[47]), .B(n1453), .Z(\ab[7][47] ) );
  AN2 U2130 ( .A(A[47]), .B(n1449), .Z(\ab[6][47] ) );
  AN2 U2131 ( .A(n1525), .B(A[9]), .Z(\ab[9][46] ) );
  AN2 U2132 ( .A(n1525), .B(A[8]), .Z(\ab[8][46] ) );
  AN2 U2133 ( .A(n1525), .B(A[47]), .Z(\CARRYB[47][46] ) );
  AN2 U2134 ( .A(n1523), .B(A[9]), .Z(\ab[9][45] ) );
  AN2 U2135 ( .A(n1523), .B(A[8]), .Z(\ab[8][45] ) );
  AN2 U2136 ( .A(n1523), .B(A[47]), .Z(\ab[47][45] ) );
  AN2 U2137 ( .A(n1523), .B(n1525), .Z(\ab[46][45] ) );
  AN2 U2138 ( .A(A[44]), .B(A[9]), .Z(\ab[9][44] ) );
  AN2 U2139 ( .A(A[44]), .B(A[8]), .Z(\ab[8][44] ) );
  AN2 U2140 ( .A(A[44]), .B(A[47]), .Z(\ab[47][44] ) );
  AN2 U2141 ( .A(A[44]), .B(n1525), .Z(\ab[46][44] ) );
  AN2 U2142 ( .A(A[44]), .B(n1523), .Z(\ab[45][44] ) );
  AN2 U2143 ( .A(n1520), .B(A[9]), .Z(\ab[9][43] ) );
  AN2 U2144 ( .A(n1520), .B(A[47]), .Z(\ab[47][43] ) );
  AN2 U2145 ( .A(n1520), .B(n1525), .Z(\ab[46][43] ) );
  AN2 U2146 ( .A(n1520), .B(n1523), .Z(\ab[45][43] ) );
  AN2 U2147 ( .A(n1520), .B(A[44]), .Z(\ab[44][43] ) );
  AN2 U2148 ( .A(n1515), .B(A[9]), .Z(\ab[9][42] ) );
  AN2 U2149 ( .A(n1515), .B(A[47]), .Z(\ab[47][42] ) );
  AN2 U2150 ( .A(n1515), .B(n1525), .Z(\ab[46][42] ) );
  AN2 U2151 ( .A(n1515), .B(n1523), .Z(\ab[45][42] ) );
  AN2 U2152 ( .A(n1515), .B(A[44]), .Z(\ab[44][42] ) );
  AN2 U2153 ( .A(n1515), .B(n1520), .Z(\ab[43][42] ) );
  AN2 U2154 ( .A(A[41]), .B(A[9]), .Z(\ab[9][41] ) );
  AN2 U2155 ( .A(A[41]), .B(A[47]), .Z(\ab[47][41] ) );
  AN2 U2156 ( .A(A[41]), .B(n1525), .Z(\ab[46][41] ) );
  AN2 U2157 ( .A(A[41]), .B(n1523), .Z(\ab[45][41] ) );
  AN2 U2158 ( .A(A[41]), .B(A[44]), .Z(\ab[44][41] ) );
  AN2 U2159 ( .A(A[41]), .B(n1520), .Z(\ab[43][41] ) );
  AN2 U2160 ( .A(A[41]), .B(n1515), .Z(\ab[42][41] ) );
  AN2 U2161 ( .A(n1510), .B(A[9]), .Z(\ab[9][40] ) );
  AN2 U2162 ( .A(n1510), .B(A[47]), .Z(\ab[47][40] ) );
  AN2 U2163 ( .A(n1510), .B(n1525), .Z(\ab[46][40] ) );
  AN2 U2164 ( .A(n1510), .B(n1523), .Z(\ab[45][40] ) );
  AN2 U2165 ( .A(n1510), .B(A[44]), .Z(\ab[44][40] ) );
  AN2 U2166 ( .A(n1510), .B(n1520), .Z(\ab[43][40] ) );
  AN2 U2167 ( .A(n1510), .B(n1515), .Z(\ab[42][40] ) );
  AN2 U2168 ( .A(n1510), .B(A[41]), .Z(\ab[41][40] ) );
  AN2 U2169 ( .A(n1507), .B(A[47]), .Z(\ab[47][39] ) );
  AN2 U2170 ( .A(n1507), .B(n1525), .Z(\ab[46][39] ) );
  AN2 U2171 ( .A(n1507), .B(n1523), .Z(\ab[45][39] ) );
  AN2 U2172 ( .A(n1507), .B(A[44]), .Z(\ab[44][39] ) );
  AN2 U2173 ( .A(n1507), .B(n1520), .Z(\ab[43][39] ) );
  AN2 U2174 ( .A(n1507), .B(n1515), .Z(\ab[42][39] ) );
  AN2 U2175 ( .A(n1507), .B(A[41]), .Z(\ab[41][39] ) );
  AN2 U2176 ( .A(n1507), .B(n1510), .Z(\ab[40][39] ) );
  AN2 U2177 ( .A(A[38]), .B(A[47]), .Z(\ab[47][38] ) );
  AN2 U2178 ( .A(A[38]), .B(n1526), .Z(\ab[46][38] ) );
  AN2 U2179 ( .A(A[38]), .B(n1523), .Z(\ab[45][38] ) );
  AN2 U2180 ( .A(A[38]), .B(A[44]), .Z(\ab[44][38] ) );
  AN2 U2181 ( .A(A[38]), .B(n1520), .Z(\ab[43][38] ) );
  AN2 U2182 ( .A(A[38]), .B(n1515), .Z(\ab[42][38] ) );
  AN2 U2183 ( .A(A[38]), .B(A[41]), .Z(\ab[41][38] ) );
  AN2 U2184 ( .A(A[38]), .B(n1510), .Z(\ab[40][38] ) );
  AN2 U2185 ( .A(A[38]), .B(n1507), .Z(\ab[39][38] ) );
  AN2 U2186 ( .A(n1505), .B(A[47]), .Z(\ab[47][37] ) );
  AN2 U2187 ( .A(n1505), .B(n1526), .Z(\ab[46][37] ) );
  AN2 U2188 ( .A(n1505), .B(A[45]), .Z(\ab[45][37] ) );
  AN2 U2189 ( .A(n1505), .B(A[44]), .Z(\ab[44][37] ) );
  AN2 U2190 ( .A(n1505), .B(n1520), .Z(\ab[43][37] ) );
  AN2 U2191 ( .A(n1505), .B(n1515), .Z(\ab[42][37] ) );
  AN2 U2192 ( .A(n1505), .B(A[41]), .Z(\ab[41][37] ) );
  AN2 U2193 ( .A(n1505), .B(n1510), .Z(\ab[40][37] ) );
  AN2 U2194 ( .A(n1505), .B(n1507), .Z(\ab[39][37] ) );
  AN2 U2195 ( .A(n1505), .B(A[38]), .Z(\ab[38][37] ) );
  AN2 U2196 ( .A(\ab[36][36] ), .B(A[47]), .Z(\ab[47][36] ) );
  AN2 U2197 ( .A(\ab[36][36] ), .B(n1526), .Z(\ab[46][36] ) );
  AN2 U2198 ( .A(\ab[36][36] ), .B(A[45]), .Z(\ab[45][36] ) );
  AN2 U2199 ( .A(\ab[36][36] ), .B(A[44]), .Z(\ab[44][36] ) );
  AN2 U2200 ( .A(\ab[36][36] ), .B(n1521), .Z(\ab[43][36] ) );
  AN2 U2201 ( .A(\ab[36][36] ), .B(n1516), .Z(\ab[42][36] ) );
  AN2 U2202 ( .A(\ab[36][36] ), .B(A[41]), .Z(\ab[41][36] ) );
  AN2 U2203 ( .A(\ab[36][36] ), .B(n1511), .Z(\ab[40][36] ) );
  AN2 U2204 ( .A(\ab[36][36] ), .B(n1507), .Z(\ab[39][36] ) );
  AN2 U2205 ( .A(\ab[36][36] ), .B(A[38]), .Z(\ab[38][36] ) );
  AN2 U2206 ( .A(\ab[36][36] ), .B(n1505), .Z(\ab[37][36] ) );
  AN2 U2207 ( .A(n1500), .B(A[47]), .Z(\ab[47][35] ) );
  AN2 U2208 ( .A(n1500), .B(n1526), .Z(\ab[46][35] ) );
  AN2 U2209 ( .A(n1500), .B(A[45]), .Z(\ab[45][35] ) );
  AN2 U2210 ( .A(n1500), .B(A[44]), .Z(\ab[44][35] ) );
  AN2 U2211 ( .A(n1500), .B(n1521), .Z(\ab[43][35] ) );
  AN2 U2212 ( .A(n1500), .B(n1516), .Z(\ab[42][35] ) );
  AN2 U2213 ( .A(n1500), .B(A[41]), .Z(\ab[41][35] ) );
  AN2 U2214 ( .A(n1500), .B(n1511), .Z(\ab[40][35] ) );
  AN2 U2215 ( .A(n1500), .B(n1508), .Z(\ab[39][35] ) );
  AN2 U2216 ( .A(n1500), .B(A[38]), .Z(\ab[38][35] ) );
  AN2 U2217 ( .A(n1500), .B(A[37]), .Z(\ab[37][35] ) );
  AN2 U2218 ( .A(n1501), .B(\ab[36][36] ), .Z(\ab[36][35] ) );
  AN2 U2219 ( .A(\ab[34][34] ), .B(A[47]), .Z(\ab[47][34] ) );
  AN2 U2220 ( .A(\ab[34][34] ), .B(n1526), .Z(\ab[46][34] ) );
  AN2 U2221 ( .A(\ab[34][34] ), .B(A[45]), .Z(\ab[45][34] ) );
  AN2 U2222 ( .A(\ab[34][34] ), .B(A[44]), .Z(\ab[44][34] ) );
  AN2 U2223 ( .A(\ab[34][34] ), .B(n1521), .Z(\ab[43][34] ) );
  AN2 U2224 ( .A(\ab[34][34] ), .B(n1516), .Z(\ab[42][34] ) );
  AN2 U2225 ( .A(\ab[34][34] ), .B(A[41]), .Z(\ab[41][34] ) );
  AN2 U2226 ( .A(\ab[34][34] ), .B(n1511), .Z(\ab[40][34] ) );
  AN2 U2227 ( .A(\ab[34][34] ), .B(n1508), .Z(\ab[39][34] ) );
  AN2 U2228 ( .A(\ab[34][34] ), .B(A[38]), .Z(\ab[38][34] ) );
  AN2 U2229 ( .A(\ab[34][34] ), .B(A[37]), .Z(\ab[37][34] ) );
  AN2 U2230 ( .A(\ab[34][34] ), .B(\ab[36][36] ), .Z(\ab[36][34] ) );
  AN2 U2231 ( .A(\ab[34][34] ), .B(n1501), .Z(\ab[35][34] ) );
  AN2 U2232 ( .A(A[33]), .B(A[47]), .Z(\ab[47][33] ) );
  AN2 U2233 ( .A(A[33]), .B(n1526), .Z(\ab[46][33] ) );
  AN2 U2234 ( .A(A[33]), .B(A[45]), .Z(\ab[45][33] ) );
  AN2 U2235 ( .A(A[33]), .B(A[44]), .Z(\ab[44][33] ) );
  AN2 U2236 ( .A(A[33]), .B(n1521), .Z(\ab[43][33] ) );
  AN2 U2237 ( .A(A[33]), .B(n1516), .Z(\ab[42][33] ) );
  AN2 U2238 ( .A(A[33]), .B(A[41]), .Z(\ab[41][33] ) );
  AN2 U2239 ( .A(A[33]), .B(n1511), .Z(\ab[40][33] ) );
  AN2 U2240 ( .A(A[33]), .B(n1508), .Z(\ab[39][33] ) );
  AN2 U2241 ( .A(A[33]), .B(A[38]), .Z(\ab[38][33] ) );
  AN2 U2242 ( .A(A[33]), .B(n1505), .Z(\ab[37][33] ) );
  AN2 U2243 ( .A(A[33]), .B(\ab[36][36] ), .Z(\ab[36][33] ) );
  AN2 U2244 ( .A(A[33]), .B(n1501), .Z(\ab[35][33] ) );
  AN2 U2245 ( .A(A[33]), .B(\ab[34][34] ), .Z(\ab[34][33] ) );
  AN2 U2246 ( .A(A[32]), .B(A[47]), .Z(\ab[47][32] ) );
  AN2 U2247 ( .A(A[32]), .B(n1526), .Z(\ab[46][32] ) );
  AN2 U2248 ( .A(A[32]), .B(A[45]), .Z(\ab[45][32] ) );
  AN2 U2249 ( .A(A[32]), .B(A[44]), .Z(\ab[44][32] ) );
  AN2 U2250 ( .A(A[32]), .B(n1521), .Z(\ab[43][32] ) );
  AN2 U2251 ( .A(A[32]), .B(n1516), .Z(\ab[42][32] ) );
  AN2 U2252 ( .A(A[32]), .B(A[41]), .Z(\ab[41][32] ) );
  AN2 U2253 ( .A(A[32]), .B(n1511), .Z(\ab[40][32] ) );
  AN2 U2254 ( .A(A[32]), .B(n1508), .Z(\ab[39][32] ) );
  AN2 U2255 ( .A(A[32]), .B(A[38]), .Z(\ab[38][32] ) );
  AN2 U2256 ( .A(A[32]), .B(n1505), .Z(\ab[37][32] ) );
  AN2 U2257 ( .A(A[32]), .B(\ab[36][36] ), .Z(\ab[36][32] ) );
  AN2 U2258 ( .A(A[32]), .B(n1501), .Z(\ab[35][32] ) );
  AN2 U2259 ( .A(A[32]), .B(\ab[34][34] ), .Z(\ab[34][32] ) );
  AN2 U2260 ( .A(A[32]), .B(A[33]), .Z(\ab[33][32] ) );
  AN2 U2261 ( .A(n1493), .B(A[47]), .Z(\ab[47][31] ) );
  AN2 U2262 ( .A(n1493), .B(n1526), .Z(\ab[46][31] ) );
  AN2 U2263 ( .A(n1493), .B(A[45]), .Z(\ab[45][31] ) );
  AN2 U2264 ( .A(n1493), .B(A[44]), .Z(\ab[44][31] ) );
  AN2 U2265 ( .A(n1493), .B(n1521), .Z(\ab[43][31] ) );
  AN2 U2266 ( .A(n1493), .B(n1516), .Z(\ab[42][31] ) );
  AN2 U2267 ( .A(n1493), .B(A[41]), .Z(\ab[41][31] ) );
  AN2 U2268 ( .A(n1493), .B(n1511), .Z(\ab[40][31] ) );
  AN2 U2269 ( .A(n1493), .B(n1508), .Z(\ab[39][31] ) );
  AN2 U2270 ( .A(n1493), .B(A[38]), .Z(\ab[38][31] ) );
  AN2 U2271 ( .A(n1493), .B(n1505), .Z(\ab[37][31] ) );
  AN2 U2272 ( .A(n1494), .B(\ab[36][36] ), .Z(\ab[36][31] ) );
  AN2 U2273 ( .A(n1494), .B(n1501), .Z(\ab[35][31] ) );
  AN2 U2274 ( .A(n1494), .B(\ab[34][34] ), .Z(\ab[34][31] ) );
  AN2 U2275 ( .A(n1494), .B(A[33]), .Z(\ab[33][31] ) );
  AN2 U2276 ( .A(n1494), .B(A[32]), .Z(\ab[32][31] ) );
  AN2 U2277 ( .A(A[30]), .B(A[47]), .Z(\ab[47][30] ) );
  AN2 U2278 ( .A(A[30]), .B(n1526), .Z(\ab[46][30] ) );
  AN2 U2279 ( .A(A[30]), .B(A[45]), .Z(\ab[45][30] ) );
  AN2 U2280 ( .A(A[30]), .B(A[44]), .Z(\ab[44][30] ) );
  AN2 U2281 ( .A(A[30]), .B(n1521), .Z(\ab[43][30] ) );
  AN2 U2282 ( .A(A[30]), .B(n1516), .Z(\ab[42][30] ) );
  AN2 U2283 ( .A(A[30]), .B(A[41]), .Z(\ab[41][30] ) );
  AN2 U2284 ( .A(A[30]), .B(n1511), .Z(\ab[40][30] ) );
  AN2 U2285 ( .A(A[30]), .B(n1508), .Z(\ab[39][30] ) );
  AN2 U2286 ( .A(A[30]), .B(A[38]), .Z(\ab[38][30] ) );
  AN2 U2287 ( .A(A[30]), .B(n1505), .Z(\ab[37][30] ) );
  AN2 U2288 ( .A(A[30]), .B(\ab[36][36] ), .Z(\ab[36][30] ) );
  AN2 U2289 ( .A(A[30]), .B(n1501), .Z(\ab[35][30] ) );
  AN2 U2290 ( .A(A[30]), .B(\ab[34][34] ), .Z(\ab[34][30] ) );
  AN2 U2291 ( .A(A[30]), .B(A[33]), .Z(\ab[33][30] ) );
  AN2 U2292 ( .A(A[30]), .B(A[32]), .Z(\ab[32][30] ) );
  AN2 U2293 ( .A(A[30]), .B(n1494), .Z(\ab[31][30] ) );
  AN2 U2294 ( .A(A[29]), .B(A[47]), .Z(\ab[47][29] ) );
  AN2 U2295 ( .A(A[29]), .B(n1526), .Z(\ab[46][29] ) );
  AN2 U2296 ( .A(A[29]), .B(A[45]), .Z(\ab[45][29] ) );
  AN2 U2297 ( .A(A[29]), .B(A[44]), .Z(\ab[44][29] ) );
  AN2 U2298 ( .A(A[29]), .B(n1521), .Z(\ab[43][29] ) );
  AN2 U2299 ( .A(A[29]), .B(n1516), .Z(\ab[42][29] ) );
  AN2 U2300 ( .A(A[29]), .B(A[41]), .Z(\ab[41][29] ) );
  AN2 U2301 ( .A(A[29]), .B(n1511), .Z(\ab[40][29] ) );
  AN2 U2302 ( .A(A[29]), .B(n1508), .Z(\ab[39][29] ) );
  AN2 U2303 ( .A(A[29]), .B(A[38]), .Z(\ab[38][29] ) );
  AN2 U2304 ( .A(A[29]), .B(n1505), .Z(\ab[37][29] ) );
  AN2 U2305 ( .A(n1491), .B(\ab[36][36] ), .Z(\ab[36][29] ) );
  AN2 U2306 ( .A(n1491), .B(n1501), .Z(\ab[35][29] ) );
  AN2 U2307 ( .A(n1491), .B(\ab[34][34] ), .Z(\ab[34][29] ) );
  AN2 U2308 ( .A(n1491), .B(A[33]), .Z(\ab[33][29] ) );
  AN2 U2309 ( .A(n1491), .B(A[32]), .Z(\ab[32][29] ) );
  AN2 U2310 ( .A(n1491), .B(n1494), .Z(\ab[31][29] ) );
  AN2 U2311 ( .A(n1491), .B(A[30]), .Z(\ab[30][29] ) );
  AN2 U2312 ( .A(n1487), .B(A[47]), .Z(\ab[47][28] ) );
  AN2 U2313 ( .A(n1487), .B(n1526), .Z(\ab[46][28] ) );
  AN2 U2314 ( .A(n1487), .B(A[45]), .Z(\ab[45][28] ) );
  AN2 U2315 ( .A(n1487), .B(A[44]), .Z(\ab[44][28] ) );
  AN2 U2316 ( .A(n1487), .B(n1521), .Z(\ab[43][28] ) );
  AN2 U2317 ( .A(n1487), .B(n1516), .Z(\ab[42][28] ) );
  AN2 U2318 ( .A(n1487), .B(A[41]), .Z(\ab[41][28] ) );
  AN2 U2319 ( .A(n1487), .B(n1511), .Z(\ab[40][28] ) );
  AN2 U2320 ( .A(n1487), .B(n1508), .Z(\ab[39][28] ) );
  AN2 U2321 ( .A(n1487), .B(A[38]), .Z(\ab[38][28] ) );
  AN2 U2322 ( .A(n1487), .B(n1505), .Z(\ab[37][28] ) );
  AN2 U2323 ( .A(n1488), .B(\ab[36][36] ), .Z(\ab[36][28] ) );
  AN2 U2324 ( .A(n1488), .B(n1501), .Z(\ab[35][28] ) );
  AN2 U2325 ( .A(n1488), .B(\ab[34][34] ), .Z(\ab[34][28] ) );
  AN2 U2326 ( .A(n1488), .B(A[33]), .Z(\ab[33][28] ) );
  AN2 U2327 ( .A(n1488), .B(A[32]), .Z(\ab[32][28] ) );
  AN2 U2328 ( .A(n1488), .B(n1494), .Z(\ab[31][28] ) );
  AN2 U2329 ( .A(n1488), .B(A[30]), .Z(\ab[30][28] ) );
  AN2 U2330 ( .A(n1488), .B(n1491), .Z(\ab[29][28] ) );
  AN2 U2331 ( .A(n1483), .B(A[47]), .Z(\ab[47][27] ) );
  AN2 U2332 ( .A(n1483), .B(n1526), .Z(\ab[46][27] ) );
  AN2 U2333 ( .A(n1483), .B(A[45]), .Z(\ab[45][27] ) );
  AN2 U2334 ( .A(n1483), .B(A[44]), .Z(\ab[44][27] ) );
  AN2 U2335 ( .A(n1483), .B(n1521), .Z(\ab[43][27] ) );
  AN2 U2336 ( .A(n1483), .B(n1516), .Z(\ab[42][27] ) );
  AN2 U2337 ( .A(n1483), .B(A[41]), .Z(\ab[41][27] ) );
  AN2 U2338 ( .A(n1483), .B(n1511), .Z(\ab[40][27] ) );
  AN2 U2339 ( .A(n1483), .B(n1508), .Z(\ab[39][27] ) );
  AN2 U2340 ( .A(n1483), .B(A[38]), .Z(\ab[38][27] ) );
  AN2 U2341 ( .A(n1483), .B(n1505), .Z(\ab[37][27] ) );
  AN2 U2342 ( .A(n1484), .B(\ab[36][36] ), .Z(\ab[36][27] ) );
  AN2 U2343 ( .A(n1484), .B(n1501), .Z(\ab[35][27] ) );
  AN2 U2344 ( .A(n1484), .B(\ab[34][34] ), .Z(\ab[34][27] ) );
  AN2 U2345 ( .A(n1484), .B(A[33]), .Z(\ab[33][27] ) );
  AN2 U2346 ( .A(n1484), .B(A[32]), .Z(\ab[32][27] ) );
  AN2 U2347 ( .A(n1484), .B(n1494), .Z(\ab[31][27] ) );
  AN2 U2348 ( .A(n1484), .B(A[30]), .Z(\ab[30][27] ) );
  AN2 U2349 ( .A(n1484), .B(n1491), .Z(\ab[29][27] ) );
  AN2 U2350 ( .A(n1484), .B(n1488), .Z(\ab[28][27] ) );
  AN2 U2351 ( .A(\ab[26][26] ), .B(A[47]), .Z(\ab[47][26] ) );
  AN2 U2352 ( .A(\ab[26][26] ), .B(A[46]), .Z(\ab[46][26] ) );
  AN2 U2353 ( .A(\ab[26][26] ), .B(A[45]), .Z(\ab[45][26] ) );
  AN2 U2354 ( .A(\ab[26][26] ), .B(A[44]), .Z(\ab[44][26] ) );
  AN2 U2355 ( .A(\ab[26][26] ), .B(n1521), .Z(\ab[43][26] ) );
  AN2 U2356 ( .A(\ab[26][26] ), .B(n1516), .Z(\ab[42][26] ) );
  AN2 U2357 ( .A(\ab[26][26] ), .B(A[41]), .Z(\ab[41][26] ) );
  AN2 U2358 ( .A(\ab[26][26] ), .B(n1511), .Z(\ab[40][26] ) );
  AN2 U2359 ( .A(\ab[26][26] ), .B(n1508), .Z(\ab[39][26] ) );
  AN2 U2360 ( .A(\ab[26][26] ), .B(A[38]), .Z(\ab[38][26] ) );
  AN2 U2361 ( .A(\ab[26][26] ), .B(n1505), .Z(\ab[37][26] ) );
  AN2 U2362 ( .A(\ab[26][26] ), .B(\ab[36][36] ), .Z(\ab[36][26] ) );
  AN2 U2363 ( .A(\ab[26][26] ), .B(n1501), .Z(\ab[35][26] ) );
  AN2 U2364 ( .A(\ab[26][26] ), .B(\ab[34][34] ), .Z(\ab[34][26] ) );
  AN2 U2365 ( .A(\ab[26][26] ), .B(A[33]), .Z(\ab[33][26] ) );
  AN2 U2366 ( .A(\ab[26][26] ), .B(A[32]), .Z(\ab[32][26] ) );
  AN2 U2367 ( .A(\ab[26][26] ), .B(n1494), .Z(\ab[31][26] ) );
  AN2 U2368 ( .A(\ab[26][26] ), .B(A[30]), .Z(\ab[30][26] ) );
  AN2 U2369 ( .A(\ab[26][26] ), .B(n1491), .Z(\ab[29][26] ) );
  AN2 U2370 ( .A(\ab[26][26] ), .B(n1488), .Z(\ab[28][26] ) );
  AN2 U2371 ( .A(\ab[26][26] ), .B(n1484), .Z(\ab[27][26] ) );
  AN2 U2372 ( .A(A[25]), .B(A[47]), .Z(\ab[47][25] ) );
  AN2 U2373 ( .A(A[25]), .B(A[46]), .Z(\ab[46][25] ) );
  AN2 U2374 ( .A(A[25]), .B(A[45]), .Z(\ab[45][25] ) );
  AN2 U2375 ( .A(A[25]), .B(A[44]), .Z(\ab[44][25] ) );
  AN2 U2376 ( .A(A[25]), .B(n1521), .Z(\ab[43][25] ) );
  AN2 U2377 ( .A(A[25]), .B(n1516), .Z(\ab[42][25] ) );
  AN2 U2378 ( .A(A[25]), .B(A[41]), .Z(\ab[41][25] ) );
  AN2 U2379 ( .A(A[25]), .B(n1511), .Z(\ab[40][25] ) );
  AN2 U2380 ( .A(A[25]), .B(n1508), .Z(\ab[39][25] ) );
  AN2 U2381 ( .A(A[25]), .B(A[38]), .Z(\ab[38][25] ) );
  AN2 U2382 ( .A(A[25]), .B(n1505), .Z(\ab[37][25] ) );
  AN2 U2383 ( .A(A[25]), .B(\ab[36][36] ), .Z(\ab[36][25] ) );
  AN2 U2384 ( .A(A[25]), .B(n1501), .Z(\ab[35][25] ) );
  AN2 U2385 ( .A(A[25]), .B(\ab[34][34] ), .Z(\ab[34][25] ) );
  AN2 U2386 ( .A(A[25]), .B(A[33]), .Z(\ab[33][25] ) );
  AN2 U2387 ( .A(A[25]), .B(A[32]), .Z(\ab[32][25] ) );
  AN2 U2388 ( .A(A[25]), .B(n1494), .Z(\ab[31][25] ) );
  AN2 U2389 ( .A(A[25]), .B(A[30]), .Z(\ab[30][25] ) );
  AN2 U2390 ( .A(A[25]), .B(n1491), .Z(\ab[29][25] ) );
  AN2 U2391 ( .A(A[25]), .B(n1488), .Z(\ab[28][25] ) );
  AN2 U2392 ( .A(A[25]), .B(n1484), .Z(\ab[27][25] ) );
  AN2 U2393 ( .A(A[25]), .B(\ab[26][26] ), .Z(\ab[26][25] ) );
  AN2 U2394 ( .A(n1479), .B(A[47]), .Z(\ab[47][24] ) );
  AN2 U2395 ( .A(n1479), .B(A[46]), .Z(\ab[46][24] ) );
  AN2 U2396 ( .A(n1479), .B(A[45]), .Z(\ab[45][24] ) );
  AN2 U2397 ( .A(n1479), .B(A[44]), .Z(\ab[44][24] ) );
  AN2 U2398 ( .A(n1479), .B(A[43]), .Z(\ab[43][24] ) );
  AN2 U2399 ( .A(n1479), .B(n1517), .Z(\ab[42][24] ) );
  AN2 U2400 ( .A(n1479), .B(A[41]), .Z(\ab[41][24] ) );
  AN2 U2401 ( .A(n1479), .B(n1512), .Z(\ab[40][24] ) );
  AN2 U2402 ( .A(n1479), .B(n1508), .Z(\ab[39][24] ) );
  AN2 U2403 ( .A(n1479), .B(A[38]), .Z(\ab[38][24] ) );
  AN2 U2404 ( .A(n1479), .B(n1505), .Z(\ab[37][24] ) );
  AN2 U2405 ( .A(n1480), .B(\ab[36][36] ), .Z(\ab[36][24] ) );
  AN2 U2406 ( .A(n1480), .B(n1501), .Z(\ab[35][24] ) );
  AN2 U2407 ( .A(n1480), .B(\ab[34][34] ), .Z(\ab[34][24] ) );
  AN2 U2408 ( .A(n1480), .B(A[33]), .Z(\ab[33][24] ) );
  AN2 U2409 ( .A(n1480), .B(A[32]), .Z(\ab[32][24] ) );
  AN2 U2410 ( .A(n1480), .B(n1494), .Z(\ab[31][24] ) );
  AN2 U2411 ( .A(n1480), .B(A[30]), .Z(\ab[30][24] ) );
  AN2 U2412 ( .A(n1480), .B(n1491), .Z(\ab[29][24] ) );
  AN2 U2413 ( .A(n1480), .B(n1488), .Z(\ab[28][24] ) );
  AN2 U2414 ( .A(n1480), .B(n1484), .Z(\ab[27][24] ) );
  AN2 U2415 ( .A(n1480), .B(\ab[26][26] ), .Z(\ab[26][24] ) );
  AN2 U2416 ( .A(n1480), .B(A[25]), .Z(\ab[25][24] ) );
  AN2 U2417 ( .A(A[23]), .B(A[47]), .Z(\ab[47][23] ) );
  AN2 U2418 ( .A(A[23]), .B(A[46]), .Z(\ab[46][23] ) );
  AN2 U2419 ( .A(A[23]), .B(A[45]), .Z(\ab[45][23] ) );
  AN2 U2420 ( .A(A[23]), .B(A[44]), .Z(\ab[44][23] ) );
  AN2 U2421 ( .A(A[23]), .B(n1521), .Z(\ab[43][23] ) );
  AN2 U2422 ( .A(A[23]), .B(n1517), .Z(\ab[42][23] ) );
  AN2 U2423 ( .A(A[23]), .B(A[41]), .Z(\ab[41][23] ) );
  AN2 U2424 ( .A(A[23]), .B(n1512), .Z(\ab[40][23] ) );
  AN2 U2425 ( .A(A[23]), .B(n1508), .Z(\ab[39][23] ) );
  AN2 U2426 ( .A(A[23]), .B(A[38]), .Z(\ab[38][23] ) );
  AN2 U2427 ( .A(A[23]), .B(n1505), .Z(\ab[37][23] ) );
  AN2 U2428 ( .A(A[23]), .B(\ab[36][36] ), .Z(\ab[36][23] ) );
  AN2 U2429 ( .A(A[23]), .B(n1502), .Z(\ab[35][23] ) );
  AN2 U2430 ( .A(A[23]), .B(\ab[34][34] ), .Z(\ab[34][23] ) );
  AN2 U2431 ( .A(A[23]), .B(A[33]), .Z(\ab[33][23] ) );
  AN2 U2432 ( .A(A[23]), .B(A[32]), .Z(\ab[32][23] ) );
  AN2 U2433 ( .A(A[23]), .B(n1495), .Z(\ab[31][23] ) );
  AN2 U2434 ( .A(A[23]), .B(A[30]), .Z(\ab[30][23] ) );
  AN2 U2435 ( .A(A[23]), .B(A[29]), .Z(\ab[29][23] ) );
  AN2 U2436 ( .A(A[23]), .B(n1489), .Z(\ab[28][23] ) );
  AN2 U2437 ( .A(A[23]), .B(n1485), .Z(\ab[27][23] ) );
  AN2 U2438 ( .A(A[23]), .B(\ab[26][26] ), .Z(\ab[26][23] ) );
  AN2 U2439 ( .A(A[23]), .B(A[25]), .Z(\ab[25][23] ) );
  AN2 U2440 ( .A(A[23]), .B(n1479), .Z(\ab[24][23] ) );
  AN2 U2441 ( .A(n1474), .B(A[47]), .Z(\ab[47][22] ) );
  AN2 U2442 ( .A(n1474), .B(n1526), .Z(\ab[46][22] ) );
  AN2 U2443 ( .A(n1474), .B(A[45]), .Z(\ab[45][22] ) );
  AN2 U2444 ( .A(n1474), .B(A[44]), .Z(\ab[44][22] ) );
  AN2 U2445 ( .A(n1474), .B(n1521), .Z(\ab[43][22] ) );
  AN2 U2446 ( .A(n1474), .B(n1517), .Z(\ab[42][22] ) );
  AN2 U2447 ( .A(n1474), .B(A[41]), .Z(\ab[41][22] ) );
  AN2 U2448 ( .A(n1474), .B(n1512), .Z(\ab[40][22] ) );
  AN2 U2449 ( .A(n1474), .B(n1508), .Z(\ab[39][22] ) );
  AN2 U2450 ( .A(n1474), .B(A[38]), .Z(\ab[38][22] ) );
  AN2 U2451 ( .A(n1474), .B(n1505), .Z(\ab[37][22] ) );
  AN2 U2452 ( .A(n1475), .B(\ab[36][36] ), .Z(\ab[36][22] ) );
  AN2 U2453 ( .A(n1475), .B(n1502), .Z(\ab[35][22] ) );
  AN2 U2454 ( .A(n1475), .B(\ab[34][34] ), .Z(\ab[34][22] ) );
  AN2 U2455 ( .A(n1475), .B(A[33]), .Z(\ab[33][22] ) );
  AN2 U2456 ( .A(n1475), .B(A[32]), .Z(\ab[32][22] ) );
  AN2 U2457 ( .A(n1475), .B(n1495), .Z(\ab[31][22] ) );
  AN2 U2458 ( .A(n1475), .B(A[30]), .Z(\ab[30][22] ) );
  AN2 U2459 ( .A(n1475), .B(A[29]), .Z(\ab[29][22] ) );
  AN2 U2460 ( .A(n1475), .B(n1489), .Z(\ab[28][22] ) );
  AN2 U2461 ( .A(n1475), .B(n1485), .Z(\ab[27][22] ) );
  AN2 U2462 ( .A(n1475), .B(\ab[26][26] ), .Z(\ab[26][22] ) );
  AN2 U2463 ( .A(n1475), .B(A[25]), .Z(\ab[25][22] ) );
  AN2 U2464 ( .A(n1476), .B(n1479), .Z(\ab[24][22] ) );
  AN2 U2465 ( .A(n1476), .B(A[23]), .Z(\ab[23][22] ) );
  AN2 U2466 ( .A(A[21]), .B(A[47]), .Z(\ab[47][21] ) );
  AN2 U2467 ( .A(A[21]), .B(n1526), .Z(\ab[46][21] ) );
  AN2 U2468 ( .A(A[21]), .B(A[45]), .Z(\ab[45][21] ) );
  AN2 U2469 ( .A(A[21]), .B(A[44]), .Z(\ab[44][21] ) );
  AN2 U2470 ( .A(A[21]), .B(n1521), .Z(\ab[43][21] ) );
  AN2 U2471 ( .A(A[21]), .B(n1517), .Z(\ab[42][21] ) );
  AN2 U2472 ( .A(A[21]), .B(A[41]), .Z(\ab[41][21] ) );
  AN2 U2473 ( .A(A[21]), .B(n1512), .Z(\ab[40][21] ) );
  AN2 U2474 ( .A(A[21]), .B(n1508), .Z(\ab[39][21] ) );
  AN2 U2475 ( .A(A[21]), .B(A[38]), .Z(\ab[38][21] ) );
  AN2 U2476 ( .A(A[21]), .B(n1505), .Z(\ab[37][21] ) );
  AN2 U2477 ( .A(A[21]), .B(\ab[36][36] ), .Z(\ab[36][21] ) );
  AN2 U2478 ( .A(A[21]), .B(n1502), .Z(\ab[35][21] ) );
  AN2 U2479 ( .A(A[21]), .B(\ab[34][34] ), .Z(\ab[34][21] ) );
  AN2 U2480 ( .A(A[21]), .B(A[33]), .Z(\ab[33][21] ) );
  AN2 U2481 ( .A(A[21]), .B(A[32]), .Z(\ab[32][21] ) );
  AN2 U2482 ( .A(A[21]), .B(n1495), .Z(\ab[31][21] ) );
  AN2 U2483 ( .A(A[21]), .B(A[30]), .Z(\ab[30][21] ) );
  AN2 U2484 ( .A(A[21]), .B(A[29]), .Z(\ab[29][21] ) );
  AN2 U2485 ( .A(A[21]), .B(n1489), .Z(\ab[28][21] ) );
  AN2 U2486 ( .A(A[21]), .B(n1485), .Z(\ab[27][21] ) );
  AN2 U2487 ( .A(A[21]), .B(\ab[26][26] ), .Z(\ab[26][21] ) );
  AN2 U2488 ( .A(A[21]), .B(A[25]), .Z(\ab[25][21] ) );
  AN2 U2489 ( .A(A[21]), .B(n1479), .Z(\ab[24][21] ) );
  AN2 U2490 ( .A(A[21]), .B(A[23]), .Z(\ab[23][21] ) );
  AN2 U2491 ( .A(A[21]), .B(n1476), .Z(\ab[22][21] ) );
  AN2 U2492 ( .A(A[20]), .B(A[47]), .Z(\ab[47][20] ) );
  AN2 U2493 ( .A(A[20]), .B(n1526), .Z(\ab[46][20] ) );
  AN2 U2494 ( .A(A[20]), .B(A[45]), .Z(\ab[45][20] ) );
  AN2 U2495 ( .A(A[20]), .B(A[44]), .Z(\ab[44][20] ) );
  AN2 U2496 ( .A(A[20]), .B(n1521), .Z(\ab[43][20] ) );
  AN2 U2497 ( .A(A[20]), .B(n1517), .Z(\ab[42][20] ) );
  AN2 U2498 ( .A(A[20]), .B(A[41]), .Z(\ab[41][20] ) );
  AN2 U2499 ( .A(A[20]), .B(n1512), .Z(\ab[40][20] ) );
  AN2 U2500 ( .A(A[20]), .B(n1508), .Z(\ab[39][20] ) );
  AN2 U2501 ( .A(A[20]), .B(A[38]), .Z(\ab[38][20] ) );
  AN2 U2502 ( .A(A[20]), .B(n1505), .Z(\ab[37][20] ) );
  AN2 U2503 ( .A(A[20]), .B(\ab[36][36] ), .Z(\ab[36][20] ) );
  AN2 U2504 ( .A(A[20]), .B(n1502), .Z(\ab[35][20] ) );
  AN2 U2505 ( .A(A[20]), .B(\ab[34][34] ), .Z(\ab[34][20] ) );
  AN2 U2506 ( .A(A[20]), .B(A[33]), .Z(\ab[33][20] ) );
  AN2 U2507 ( .A(A[20]), .B(A[32]), .Z(\ab[32][20] ) );
  AN2 U2508 ( .A(A[20]), .B(n1495), .Z(\ab[31][20] ) );
  AN2 U2509 ( .A(A[20]), .B(A[30]), .Z(\ab[30][20] ) );
  AN2 U2510 ( .A(A[20]), .B(A[29]), .Z(\ab[29][20] ) );
  AN2 U2511 ( .A(A[20]), .B(n1489), .Z(\ab[28][20] ) );
  AN2 U2512 ( .A(A[20]), .B(n1485), .Z(\ab[27][20] ) );
  AN2 U2513 ( .A(A[20]), .B(\ab[26][26] ), .Z(\ab[26][20] ) );
  AN2 U2514 ( .A(A[20]), .B(A[25]), .Z(\ab[25][20] ) );
  AN2 U2515 ( .A(A[20]), .B(n1479), .Z(\ab[24][20] ) );
  AN2 U2516 ( .A(A[20]), .B(A[23]), .Z(\ab[23][20] ) );
  AN2 U2517 ( .A(A[20]), .B(n1476), .Z(\ab[22][20] ) );
  AN2 U2518 ( .A(A[20]), .B(A[21]), .Z(\ab[21][20] ) );
  AN2 U2519 ( .A(n1468), .B(A[47]), .Z(\ab[47][19] ) );
  AN2 U2520 ( .A(n1468), .B(n1526), .Z(\ab[46][19] ) );
  AN2 U2521 ( .A(n1468), .B(A[45]), .Z(\ab[45][19] ) );
  AN2 U2522 ( .A(n1468), .B(A[44]), .Z(\ab[44][19] ) );
  AN2 U2523 ( .A(n1468), .B(n1521), .Z(\ab[43][19] ) );
  AN2 U2524 ( .A(n1468), .B(n1517), .Z(\ab[42][19] ) );
  AN2 U2525 ( .A(n1468), .B(A[41]), .Z(\ab[41][19] ) );
  AN2 U2526 ( .A(n1468), .B(n1512), .Z(\ab[40][19] ) );
  AN2 U2527 ( .A(n1468), .B(n1508), .Z(\ab[39][19] ) );
  AN2 U2528 ( .A(n1468), .B(A[38]), .Z(\ab[38][19] ) );
  AN2 U2529 ( .A(n1468), .B(n1505), .Z(\ab[37][19] ) );
  AN2 U2530 ( .A(n1469), .B(\ab[36][36] ), .Z(\ab[36][19] ) );
  AN2 U2531 ( .A(n1469), .B(n1502), .Z(\ab[35][19] ) );
  AN2 U2532 ( .A(n1469), .B(\ab[34][34] ), .Z(\ab[34][19] ) );
  AN2 U2533 ( .A(n1469), .B(A[33]), .Z(\ab[33][19] ) );
  AN2 U2534 ( .A(n1469), .B(A[32]), .Z(\ab[32][19] ) );
  AN2 U2535 ( .A(n1469), .B(n1495), .Z(\ab[31][19] ) );
  AN2 U2536 ( .A(n1469), .B(A[30]), .Z(\ab[30][19] ) );
  AN2 U2537 ( .A(n1469), .B(A[29]), .Z(\ab[29][19] ) );
  AN2 U2538 ( .A(n1469), .B(n1489), .Z(\ab[28][19] ) );
  AN2 U2539 ( .A(n1469), .B(n1485), .Z(\ab[27][19] ) );
  AN2 U2540 ( .A(n1469), .B(\ab[26][26] ), .Z(\ab[26][19] ) );
  AN2 U2541 ( .A(n1469), .B(A[25]), .Z(\ab[25][19] ) );
  AN2 U2542 ( .A(n1470), .B(n1479), .Z(\ab[24][19] ) );
  AN2 U2543 ( .A(n1470), .B(A[23]), .Z(\ab[23][19] ) );
  AN2 U2544 ( .A(n1470), .B(n1476), .Z(\ab[22][19] ) );
  AN2 U2545 ( .A(n1470), .B(A[21]), .Z(\ab[21][19] ) );
  AN2 U2546 ( .A(n1470), .B(A[20]), .Z(\ab[20][19] ) );
  AN2 U2547 ( .A(\ab[18][18] ), .B(A[47]), .Z(\ab[47][18] ) );
  AN2 U2548 ( .A(\ab[18][18] ), .B(n1526), .Z(\ab[46][18] ) );
  AN2 U2549 ( .A(\ab[18][18] ), .B(A[45]), .Z(\ab[45][18] ) );
  AN2 U2550 ( .A(\ab[18][18] ), .B(A[44]), .Z(\ab[44][18] ) );
  AN2 U2551 ( .A(\ab[18][18] ), .B(n1521), .Z(\ab[43][18] ) );
  AN2 U2552 ( .A(\ab[18][18] ), .B(n1517), .Z(\ab[42][18] ) );
  AN2 U2553 ( .A(\ab[18][18] ), .B(A[41]), .Z(\ab[41][18] ) );
  AN2 U2554 ( .A(\ab[18][18] ), .B(n1512), .Z(\ab[40][18] ) );
  AN2 U2555 ( .A(\ab[18][18] ), .B(n1508), .Z(\ab[39][18] ) );
  AN2 U2556 ( .A(\ab[18][18] ), .B(A[38]), .Z(\ab[38][18] ) );
  AN2 U2557 ( .A(\ab[18][18] ), .B(n1505), .Z(\ab[37][18] ) );
  AN2 U2558 ( .A(\ab[18][18] ), .B(\ab[36][36] ), .Z(\ab[36][18] ) );
  AN2 U2559 ( .A(\ab[18][18] ), .B(n1502), .Z(\ab[35][18] ) );
  AN2 U2560 ( .A(\ab[18][18] ), .B(\ab[34][34] ), .Z(\ab[34][18] ) );
  AN2 U2561 ( .A(\ab[18][18] ), .B(A[33]), .Z(\ab[33][18] ) );
  AN2 U2562 ( .A(\ab[18][18] ), .B(A[32]), .Z(\ab[32][18] ) );
  AN2 U2563 ( .A(\ab[18][18] ), .B(n1495), .Z(\ab[31][18] ) );
  AN2 U2564 ( .A(\ab[18][18] ), .B(A[30]), .Z(\ab[30][18] ) );
  AN2 U2565 ( .A(\ab[18][18] ), .B(A[29]), .Z(\ab[29][18] ) );
  AN2 U2566 ( .A(\ab[18][18] ), .B(n1489), .Z(\ab[28][18] ) );
  AN2 U2567 ( .A(\ab[18][18] ), .B(n1485), .Z(\ab[27][18] ) );
  AN2 U2568 ( .A(\ab[18][18] ), .B(\ab[26][26] ), .Z(\ab[26][18] ) );
  AN2 U2569 ( .A(\ab[18][18] ), .B(A[25]), .Z(\ab[25][18] ) );
  AN2 U2570 ( .A(\ab[18][18] ), .B(n1479), .Z(\ab[24][18] ) );
  AN2 U2571 ( .A(\ab[18][18] ), .B(A[23]), .Z(\ab[23][18] ) );
  AN2 U2572 ( .A(\ab[18][18] ), .B(n1476), .Z(\ab[22][18] ) );
  AN2 U2573 ( .A(\ab[18][18] ), .B(A[21]), .Z(\ab[21][18] ) );
  AN2 U2574 ( .A(\ab[18][18] ), .B(A[20]), .Z(\ab[20][18] ) );
  AN2 U2575 ( .A(\ab[18][18] ), .B(n1470), .Z(\ab[19][18] ) );
  AN2 U2576 ( .A(n1464), .B(A[47]), .Z(\ab[47][17] ) );
  AN2 U2577 ( .A(n1464), .B(n1526), .Z(\ab[46][17] ) );
  AN2 U2578 ( .A(n1464), .B(n1523), .Z(\ab[45][17] ) );
  AN2 U2579 ( .A(n1464), .B(A[44]), .Z(\ab[44][17] ) );
  AN2 U2580 ( .A(n1464), .B(n1521), .Z(\ab[43][17] ) );
  AN2 U2581 ( .A(n1464), .B(n1517), .Z(\ab[42][17] ) );
  AN2 U2582 ( .A(n1464), .B(A[41]), .Z(\ab[41][17] ) );
  AN2 U2583 ( .A(n1464), .B(n1512), .Z(\ab[40][17] ) );
  AN2 U2584 ( .A(n1464), .B(n1508), .Z(\ab[39][17] ) );
  AN2 U2585 ( .A(n1464), .B(A[38]), .Z(\ab[38][17] ) );
  AN2 U2586 ( .A(n1464), .B(n1505), .Z(\ab[37][17] ) );
  AN2 U2587 ( .A(n1465), .B(\ab[36][36] ), .Z(\ab[36][17] ) );
  AN2 U2588 ( .A(n1465), .B(n1502), .Z(\ab[35][17] ) );
  AN2 U2589 ( .A(n1465), .B(\ab[34][34] ), .Z(\ab[34][17] ) );
  AN2 U2590 ( .A(n1465), .B(A[33]), .Z(\ab[33][17] ) );
  AN2 U2591 ( .A(n1465), .B(A[32]), .Z(\ab[32][17] ) );
  AN2 U2592 ( .A(n1465), .B(n1495), .Z(\ab[31][17] ) );
  AN2 U2593 ( .A(n1465), .B(A[30]), .Z(\ab[30][17] ) );
  AN2 U2594 ( .A(n1465), .B(A[29]), .Z(\ab[29][17] ) );
  AN2 U2595 ( .A(n1465), .B(n1489), .Z(\ab[28][17] ) );
  AN2 U2596 ( .A(n1465), .B(n1485), .Z(\ab[27][17] ) );
  AN2 U2597 ( .A(n1465), .B(\ab[26][26] ), .Z(\ab[26][17] ) );
  AN2 U2598 ( .A(n1465), .B(A[25]), .Z(\ab[25][17] ) );
  AN2 U2599 ( .A(n1466), .B(n1479), .Z(\ab[24][17] ) );
  AN2 U2600 ( .A(n1466), .B(A[23]), .Z(\ab[23][17] ) );
  AN2 U2601 ( .A(n1466), .B(n1476), .Z(\ab[22][17] ) );
  AN2 U2602 ( .A(n1466), .B(A[21]), .Z(\ab[21][17] ) );
  AN2 U2603 ( .A(n1466), .B(A[20]), .Z(\ab[20][17] ) );
  AN2 U2604 ( .A(n1466), .B(n1470), .Z(\ab[19][17] ) );
  AN2 U2605 ( .A(n1466), .B(\ab[18][18] ), .Z(\ab[18][17] ) );
  AN2 U2606 ( .A(A[16]), .B(A[47]), .Z(\ab[47][16] ) );
  AN2 U2607 ( .A(A[16]), .B(A[46]), .Z(\ab[46][16] ) );
  AN2 U2608 ( .A(A[16]), .B(n1523), .Z(\ab[45][16] ) );
  AN2 U2609 ( .A(A[16]), .B(A[44]), .Z(\ab[44][16] ) );
  AN2 U2610 ( .A(A[16]), .B(n1521), .Z(\ab[43][16] ) );
  AN2 U2611 ( .A(A[16]), .B(n1517), .Z(\ab[42][16] ) );
  AN2 U2612 ( .A(A[16]), .B(A[41]), .Z(\ab[41][16] ) );
  AN2 U2613 ( .A(A[16]), .B(n1512), .Z(\ab[40][16] ) );
  AN2 U2614 ( .A(A[16]), .B(n1508), .Z(\ab[39][16] ) );
  AN2 U2615 ( .A(A[16]), .B(A[38]), .Z(\ab[38][16] ) );
  AN2 U2616 ( .A(A[16]), .B(n1505), .Z(\ab[37][16] ) );
  AN2 U2617 ( .A(A[16]), .B(\ab[36][36] ), .Z(\ab[36][16] ) );
  AN2 U2618 ( .A(A[16]), .B(n1502), .Z(\ab[35][16] ) );
  AN2 U2619 ( .A(A[16]), .B(\ab[34][34] ), .Z(\ab[34][16] ) );
  AN2 U2620 ( .A(A[16]), .B(A[33]), .Z(\ab[33][16] ) );
  AN2 U2621 ( .A(A[16]), .B(A[32]), .Z(\ab[32][16] ) );
  AN2 U2622 ( .A(A[16]), .B(n1495), .Z(\ab[31][16] ) );
  AN2 U2623 ( .A(A[16]), .B(A[30]), .Z(\ab[30][16] ) );
  AN2 U2624 ( .A(A[16]), .B(A[29]), .Z(\ab[29][16] ) );
  AN2 U2625 ( .A(A[16]), .B(n1489), .Z(\ab[28][16] ) );
  AN2 U2626 ( .A(A[16]), .B(n1485), .Z(\ab[27][16] ) );
  AN2 U2627 ( .A(A[16]), .B(\ab[26][26] ), .Z(\ab[26][16] ) );
  AN2 U2628 ( .A(A[16]), .B(A[25]), .Z(\ab[25][16] ) );
  AN2 U2629 ( .A(A[16]), .B(n1479), .Z(\ab[24][16] ) );
  AN2 U2630 ( .A(A[16]), .B(A[23]), .Z(\ab[23][16] ) );
  AN2 U2631 ( .A(A[16]), .B(n1476), .Z(\ab[22][16] ) );
  AN2 U2632 ( .A(A[16]), .B(A[21]), .Z(\ab[21][16] ) );
  AN2 U2633 ( .A(A[16]), .B(A[20]), .Z(\ab[20][16] ) );
  AN2 U2634 ( .A(A[16]), .B(n1470), .Z(\ab[19][16] ) );
  AN2 U2635 ( .A(A[16]), .B(\ab[18][18] ), .Z(\ab[18][16] ) );
  AN2 U2636 ( .A(A[16]), .B(n1466), .Z(\ab[17][16] ) );
  AN2 U2637 ( .A(n1461), .B(A[47]), .Z(\ab[47][15] ) );
  AN2 U2638 ( .A(n1461), .B(A[46]), .Z(\ab[46][15] ) );
  AN2 U2639 ( .A(n1461), .B(A[45]), .Z(\ab[45][15] ) );
  AN2 U2640 ( .A(n1461), .B(A[44]), .Z(\ab[44][15] ) );
  AN2 U2641 ( .A(n1461), .B(n1521), .Z(\ab[43][15] ) );
  AN2 U2642 ( .A(n1461), .B(n1517), .Z(\ab[42][15] ) );
  AN2 U2643 ( .A(n1461), .B(A[41]), .Z(\ab[41][15] ) );
  AN2 U2644 ( .A(n1461), .B(n1512), .Z(\ab[40][15] ) );
  AN2 U2645 ( .A(n1461), .B(n1508), .Z(\ab[39][15] ) );
  AN2 U2646 ( .A(n1461), .B(A[38]), .Z(\ab[38][15] ) );
  AN2 U2647 ( .A(n1461), .B(n1505), .Z(\ab[37][15] ) );
  AN2 U2648 ( .A(A[15]), .B(\ab[36][36] ), .Z(\ab[36][15] ) );
  AN2 U2649 ( .A(A[15]), .B(n1502), .Z(\ab[35][15] ) );
  AN2 U2650 ( .A(A[15]), .B(\ab[34][34] ), .Z(\ab[34][15] ) );
  AN2 U2651 ( .A(A[15]), .B(A[33]), .Z(\ab[33][15] ) );
  AN2 U2652 ( .A(A[15]), .B(A[32]), .Z(\ab[32][15] ) );
  AN2 U2653 ( .A(A[15]), .B(n1495), .Z(\ab[31][15] ) );
  AN2 U2654 ( .A(A[15]), .B(A[30]), .Z(\ab[30][15] ) );
  AN2 U2655 ( .A(A[15]), .B(A[29]), .Z(\ab[29][15] ) );
  AN2 U2656 ( .A(A[15]), .B(n1489), .Z(\ab[28][15] ) );
  AN2 U2657 ( .A(A[15]), .B(n1485), .Z(\ab[27][15] ) );
  AN2 U2658 ( .A(A[15]), .B(\ab[26][26] ), .Z(\ab[26][15] ) );
  AN2 U2659 ( .A(A[15]), .B(A[25]), .Z(\ab[25][15] ) );
  AN2 U2660 ( .A(n1462), .B(n1479), .Z(\ab[24][15] ) );
  AN2 U2661 ( .A(n1462), .B(A[23]), .Z(\ab[23][15] ) );
  AN2 U2662 ( .A(n1462), .B(n1476), .Z(\ab[22][15] ) );
  AN2 U2663 ( .A(n1462), .B(A[21]), .Z(\ab[21][15] ) );
  AN2 U2664 ( .A(n1462), .B(A[20]), .Z(\ab[20][15] ) );
  AN2 U2665 ( .A(n1462), .B(n1470), .Z(\ab[19][15] ) );
  AN2 U2666 ( .A(n1462), .B(\ab[18][18] ), .Z(\ab[18][15] ) );
  AN2 U2667 ( .A(n1462), .B(n1466), .Z(\ab[17][15] ) );
  AN2 U2668 ( .A(n1462), .B(A[16]), .Z(\ab[16][15] ) );
  AN2 U2669 ( .A(n1459), .B(A[47]), .Z(\ab[47][14] ) );
  AN2 U2670 ( .A(n1459), .B(n1526), .Z(\ab[46][14] ) );
  AN2 U2671 ( .A(n1459), .B(A[45]), .Z(\ab[45][14] ) );
  AN2 U2672 ( .A(n1459), .B(A[44]), .Z(\ab[44][14] ) );
  AN2 U2673 ( .A(n1459), .B(A[43]), .Z(\ab[43][14] ) );
  AN2 U2674 ( .A(n1459), .B(n1517), .Z(\ab[42][14] ) );
  AN2 U2675 ( .A(n1459), .B(A[41]), .Z(\ab[41][14] ) );
  AN2 U2676 ( .A(n1459), .B(n1512), .Z(\ab[40][14] ) );
  AN2 U2677 ( .A(n1459), .B(n1508), .Z(\ab[39][14] ) );
  AN2 U2678 ( .A(n1459), .B(A[38]), .Z(\ab[38][14] ) );
  AN2 U2679 ( .A(n1459), .B(n1505), .Z(\ab[37][14] ) );
  AN2 U2680 ( .A(A[14]), .B(\ab[36][36] ), .Z(\ab[36][14] ) );
  AN2 U2681 ( .A(A[14]), .B(n1502), .Z(\ab[35][14] ) );
  AN2 U2682 ( .A(A[14]), .B(\ab[34][34] ), .Z(\ab[34][14] ) );
  AN2 U2683 ( .A(A[14]), .B(A[33]), .Z(\ab[33][14] ) );
  AN2 U2684 ( .A(A[14]), .B(A[32]), .Z(\ab[32][14] ) );
  AN2 U2685 ( .A(A[14]), .B(n1495), .Z(\ab[31][14] ) );
  AN2 U2686 ( .A(A[14]), .B(A[30]), .Z(\ab[30][14] ) );
  AN2 U2687 ( .A(A[14]), .B(A[29]), .Z(\ab[29][14] ) );
  AN2 U2688 ( .A(A[14]), .B(n1489), .Z(\ab[28][14] ) );
  AN2 U2689 ( .A(A[14]), .B(n1485), .Z(\ab[27][14] ) );
  AN2 U2690 ( .A(A[13]), .B(A[47]), .Z(\ab[47][13] ) );
  AN2 U2691 ( .A(A[13]), .B(n1525), .Z(\ab[46][13] ) );
  AN2 U2692 ( .A(A[13]), .B(n1523), .Z(\ab[45][13] ) );
  AN2 U2693 ( .A(A[13]), .B(A[44]), .Z(\ab[44][13] ) );
  AN2 U2694 ( .A(A[13]), .B(A[43]), .Z(\ab[43][13] ) );
  AN2 U2695 ( .A(A[13]), .B(n1517), .Z(\ab[42][13] ) );
  AN2 U2696 ( .A(A[13]), .B(A[41]), .Z(\ab[41][13] ) );
  AN2 U2697 ( .A(A[13]), .B(n1512), .Z(\ab[40][13] ) );
  AN2 U2698 ( .A(A[13]), .B(n1508), .Z(\ab[39][13] ) );
  AN2 U2699 ( .A(A[13]), .B(A[38]), .Z(\ab[38][13] ) );
  AN2 U2700 ( .A(A[13]), .B(n1505), .Z(\ab[37][13] ) );
  AN2 U2701 ( .A(A[13]), .B(\ab[36][36] ), .Z(\ab[36][13] ) );
  AN2 U2702 ( .A(A[13]), .B(n1502), .Z(\ab[35][13] ) );
  AN2 U2703 ( .A(A[13]), .B(\ab[34][34] ), .Z(\ab[34][13] ) );
  AN2 U2704 ( .A(A[13]), .B(A[33]), .Z(\ab[33][13] ) );
  AN2 U2705 ( .A(A[13]), .B(A[32]), .Z(\ab[32][13] ) );
  AN2 U2706 ( .A(A[13]), .B(n1495), .Z(\ab[31][13] ) );
  AN2 U2707 ( .A(A[12]), .B(A[47]), .Z(\ab[47][12] ) );
  AN2 U2708 ( .A(A[12]), .B(n1526), .Z(\ab[46][12] ) );
  AN2 U2709 ( .A(A[12]), .B(n1523), .Z(\ab[45][12] ) );
  AN2 U2710 ( .A(A[12]), .B(A[44]), .Z(\ab[44][12] ) );
  AN2 U2711 ( .A(A[12]), .B(n1521), .Z(\ab[43][12] ) );
  AN2 U2712 ( .A(A[12]), .B(n1518), .Z(\ab[42][12] ) );
  AN2 U2713 ( .A(A[12]), .B(A[41]), .Z(\ab[41][12] ) );
  AN2 U2714 ( .A(A[12]), .B(n1510), .Z(\ab[40][12] ) );
  AN2 U2715 ( .A(A[12]), .B(n1508), .Z(\ab[39][12] ) );
  AN2 U2716 ( .A(A[12]), .B(A[38]), .Z(\ab[38][12] ) );
  AN2 U2717 ( .A(A[12]), .B(n1505), .Z(\ab[37][12] ) );
  AN2 U2718 ( .A(A[12]), .B(\ab[36][36] ), .Z(\ab[36][12] ) );
  AN2 U2719 ( .A(A[12]), .B(n1502), .Z(\ab[35][12] ) );
  AN2 U2720 ( .A(A[12]), .B(\ab[34][34] ), .Z(\ab[34][12] ) );
  AN2 U2721 ( .A(A[12]), .B(A[33]), .Z(\ab[33][12] ) );
  AN2 U2722 ( .A(A[11]), .B(A[47]), .Z(\ab[47][11] ) );
  AN2 U2723 ( .A(A[11]), .B(n1526), .Z(\ab[46][11] ) );
  AN2 U2724 ( .A(A[11]), .B(n1523), .Z(\ab[45][11] ) );
  AN2 U2725 ( .A(A[11]), .B(A[44]), .Z(\ab[44][11] ) );
  AN2 U2726 ( .A(A[11]), .B(n1521), .Z(\ab[43][11] ) );
  AN2 U2727 ( .A(A[11]), .B(\ab[42][42] ), .Z(\ab[42][11] ) );
  AN2 U2728 ( .A(A[11]), .B(A[41]), .Z(\ab[41][11] ) );
  AN2 U2729 ( .A(A[11]), .B(n1510), .Z(\ab[40][11] ) );
  AN2 U2730 ( .A(A[11]), .B(n1507), .Z(\ab[39][11] ) );
  AN2 U2731 ( .A(A[11]), .B(A[38]), .Z(\ab[38][11] ) );
  AN2 U2732 ( .A(A[11]), .B(n1505), .Z(\ab[37][11] ) );
  AN2 U2733 ( .A(A[11]), .B(\ab[36][36] ), .Z(\ab[36][11] ) );
  AN2 U2734 ( .A(A[11]), .B(n1500), .Z(\ab[35][11] ) );
  AN2 U2735 ( .A(A[10]), .B(A[47]), .Z(\ab[47][10] ) );
  AN2 U2736 ( .A(A[10]), .B(n1526), .Z(\ab[46][10] ) );
  AN2 U2737 ( .A(A[10]), .B(n1523), .Z(\ab[45][10] ) );
  AN2 U2738 ( .A(A[10]), .B(A[44]), .Z(\ab[44][10] ) );
  AN2 U2739 ( .A(A[10]), .B(n1521), .Z(\ab[43][10] ) );
  AN2 U2740 ( .A(A[10]), .B(\ab[42][42] ), .Z(\ab[42][10] ) );
  AN2 U2741 ( .A(A[10]), .B(A[41]), .Z(\ab[41][10] ) );
  AN2 U2742 ( .A(A[10]), .B(n1510), .Z(\ab[40][10] ) );
  AN2 U2743 ( .A(A[10]), .B(n1507), .Z(\ab[39][10] ) );
  AN2 U2744 ( .A(A[10]), .B(A[38]), .Z(\ab[38][10] ) );
endmodule


module LOG_POLY ( clk, reset, LogIn, LogOut );
  input [47:0] LogIn;
  output [30:0] LogOut;
  input clk, reset;
  wire   N9, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N254, N255, N256, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, N277, N292, N293,
         N294, N295, N296, N297, N298, N284, N283, N282, N281, N280, N279,
         N278, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243,
         N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232,
         N231, N230, \add_1_root_sub_1_root_add_55_2/carry[6] ,
         \add_1_root_sub_1_root_add_55_2/carry[5] ,
         \add_1_root_sub_1_root_add_55_2/carry[4] ,
         \add_1_root_sub_1_root_add_55_2/carry[3] ,
         \add_1_root_sub_1_root_add_55_2/carry[2] ,
         \add_1_root_sub_1_root_add_55_2/carry[1] , n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388;
  wire   [95:0] LogInSquare;
  wire   [47:0] LogIn2;
  wire   [118:89] Term1;
  wire   [67:38] Term2;
  wire   [26:1] Term3;
  wire   [118:112] Term11;
  wire   [67:61] Term21;
  wire   [26:24] Term31;
  wire   [23:0] FractionBit;
  wire   [6:0] IntegerBits;
  wire   [22:0] LogPipe;
  wire   [29:0] Log;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136;
  assign LogOut[0] = 1'b0;

  LOG_POLY_DW02_mult_2 mult_44 ( .A({n356, n355, n354, n395, n389, n388, N171, 
        N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, 
        N184, N185, N186}), .B(LogIn2), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, N216, N215, N214, 
        N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, 
        N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, 
        N189, N188, N187, SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39}) );
  LOG_POLY_DW02_mult_1 mult_43 ( .A({n361, n360, n359, n358, n357, n406, n405, 
        n791, n397, n394, n392, N116, N117, N118, N119, N120, N121, N122, N123, 
        N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134}), 
        .B(LogInSquare), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N164, N163, N162, 
        N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, 
        N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137, N136, N135, SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135}) );
  LOG_POLY_DW01_sub_0 sub_0_root_sub_1_root_add_55_2 ( .A({N284, N283, N282, 
        N281, N280, N279, N278}), .B(Term21), .CI(1'b0), .DIFF({N298, N297, 
        N296, N295, N294, N293, N292}) );
  LOG_POLY_DW01_sub_1 sub_0_root_sub_0_root_add_52 ( .A({n792, N252, N251, 
        N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, 
        N238, N237, N236, N235, N234, N233, N232, N231, N230}), .B({1'b0, 
        Term2[60:38]}), .CI(1'b0), .DIFF({N277, N276, N275, N274, N273, N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254}) );
  LOG_POLY_DW02_mult_0 mult_39 ( .A(LogIn), .B(LogIn), .TC(1'b0), .PRODUCT({
        N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, 
        N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, 
        N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, 
        N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        SYNOPSYS_UNCONNECTED__136, N9}) );
  FD1 \LogInSquare_reg[61]  ( .D(n826), .CP(clk), .Q(LogInSquare[61]) );
  MUX21L \LogInSquare_reg[84]/U5  ( .A(LogInSquare[84]), .B(N93), .S(n5367), 
        .Z(n823) );
  FD1 \LogInSquare_reg[84]  ( .D(n824), .CP(clk), .Q(LogInSquare[84]) );
  MUX21L \LogInSquare_reg[83]/U5  ( .A(LogInSquare[83]), .B(N92), .S(n5366), 
        .Z(n821) );
  FD1 \LogInSquare_reg[83]  ( .D(n822), .CP(clk), .Q(LogInSquare[83]) );
  FD1 \LogInSquare_reg[69]  ( .D(n820), .CP(clk), .Q(LogInSquare[69]) );
  FD1 \LogInSquare_reg[81]  ( .D(n818), .CP(clk), .Q(LogInSquare[81]) );
  FD1 \LogInSquare_reg[65]  ( .D(n816), .CP(clk), .Q(LogInSquare[65]) );
  FD1 \LogInSquare_reg[77]  ( .D(n814), .CP(clk), .Q(LogInSquare[77]) );
  MUX21L \LogInSquare_reg[87]/U5  ( .A(LogInSquare[87]), .B(N96), .S(n5367), 
        .Z(n811) );
  FD1 \LogInSquare_reg[87]  ( .D(n812), .CP(clk), .Q(LogInSquare[87]) );
  MUX21L \LogInSquare_reg[85]/U5  ( .A(LogInSquare[85]), .B(N94), .S(n5367), 
        .Z(n809) );
  FD1 \LogInSquare_reg[85]  ( .D(n810), .CP(clk), .Q(LogInSquare[85]) );
  MUX21L \LogInSquare_reg[86]/U5  ( .A(LogInSquare[86]), .B(N95), .S(n5367), 
        .Z(n807) );
  FD1 \LogInSquare_reg[86]  ( .D(n808), .CP(clk), .Q(LogInSquare[86]) );
  FD1 \LogInSquare_reg[73]  ( .D(n806), .CP(clk), .Q(LogInSquare[73]) );
  FD1 \LogInSquare_reg[94]  ( .D(n804), .CP(clk), .Q(LogInSquare[94]) );
  FD1 \LogInSquare_reg[93]  ( .D(n802), .CP(clk), .Q(LogInSquare[93]) );
  FD1 \LogInSquare_reg[92]  ( .D(n800), .CP(clk), .Q(LogInSquare[92]) );
  FD1 \LogInSquare_reg[91]  ( .D(n798), .CP(clk), .Q(LogInSquare[91]) );
  FD1 \LogInSquare_reg[90]  ( .D(n796), .CP(clk), .Q(LogInSquare[90]) );
  FDS2L \Term1_reg[111]  ( .CR(1'b1), .D(N157), .LD(n5364), .CP(clk), .Q(
        Term1[111]), .QN(n793) );
  FDS2L \Term3_reg[23]  ( .CR(1'b1), .D(N220), .LD(n5363), .CP(clk), .Q(
        Term3[23]), .QN(n794) );
  FDS2L \LogInSquare_reg[1]  ( .CR(1'b1), .D(1'b0), .LD(n5362), .CP(clk), .Q(
        LogInSquare[1]) );
  FDS2L \LogInSquare_reg[0]  ( .CR(1'b1), .D(N9), .LD(n5388), .CP(clk), .Q(
        LogInSquare[0]) );
  FDS2L \LogIn2_reg[47]  ( .CR(1'b1), .D(LogIn[47]), .LD(n5388), .CP(clk), .Q(
        LogIn2[47]), .QN(n353) );
  FDS2L \LogIn2_reg[46]  ( .CR(1'b1), .D(LogIn[46]), .LD(n5388), .CP(clk), .Q(
        LogIn2[46]), .QN(n351) );
  FDS2L \LogIn2_reg[45]  ( .CR(1'b1), .D(LogIn[45]), .LD(n5388), .CP(clk), .Q(
        LogIn2[45]), .QN(n4269) );
  FDS2L \LogIn2_reg[44]  ( .CR(1'b1), .D(LogIn[44]), .LD(n5388), .CP(clk), .Q(
        LogIn2[44]), .QN(n350) );
  FDS2L \LogIn2_reg[43]  ( .CR(1'b1), .D(LogIn[43]), .LD(n5388), .CP(clk), .Q(
        LogIn2[43]) );
  FDS2L \LogIn2_reg[42]  ( .CR(1'b1), .D(LogIn[42]), .LD(n5388), .CP(clk), .Q(
        LogIn2[42]) );
  FDS2L \LogIn2_reg[41]  ( .CR(1'b1), .D(LogIn[41]), .LD(n5388), .CP(clk), .Q(
        LogIn2[41]) );
  FDS2L \LogIn2_reg[40]  ( .CR(1'b1), .D(LogIn[40]), .LD(n5388), .CP(clk), .Q(
        LogIn2[40]), .QN(n352) );
  FDS2L \Term31_reg[26]  ( .CR(1'b1), .D(Term3[26]), .LD(n5388), .CP(clk), .Q(
        Term31[26]) );
  FDS2L \Term31_reg[25]  ( .CR(1'b1), .D(Term3[25]), .LD(n5388), .CP(clk), .Q(
        Term31[25]) );
  FDS2L \Term31_reg[24]  ( .CR(1'b1), .D(Term3[24]), .LD(n5388), .CP(clk), .Q(
        Term31[24]) );
  FDS2L \Term21_reg[67]  ( .CR(1'b1), .D(Term2[67]), .LD(n5388), .CP(clk), .Q(
        Term21[67]) );
  FDS2L \Term21_reg[66]  ( .CR(1'b1), .D(Term2[66]), .LD(n5388), .CP(clk), .Q(
        Term21[66]) );
  FDS2L \Term21_reg[65]  ( .CR(1'b1), .D(Term2[65]), .LD(n5388), .CP(clk), .Q(
        Term21[65]) );
  FDS2L \Term21_reg[64]  ( .CR(1'b1), .D(Term2[64]), .LD(n5388), .CP(clk), .Q(
        Term21[64]) );
  FDS2L \Term21_reg[63]  ( .CR(1'b1), .D(Term2[63]), .LD(n5388), .CP(clk), .Q(
        Term21[63]) );
  FDS2L \Term21_reg[62]  ( .CR(1'b1), .D(Term2[62]), .LD(n5388), .CP(clk), .Q(
        Term21[62]) );
  FDS2L \Term21_reg[61]  ( .CR(1'b1), .D(Term2[61]), .LD(n5388), .CP(clk), .Q(
        Term21[61]) );
  FDS2L \Term11_reg[118]  ( .CR(1'b1), .D(Term1[118]), .LD(n5388), .CP(clk), 
        .Q(Term11[118]) );
  FDS2L \Term11_reg[117]  ( .CR(1'b1), .D(Term1[117]), .LD(n5388), .CP(clk), 
        .Q(Term11[117]) );
  FDS2L \Term11_reg[116]  ( .CR(1'b1), .D(Term1[116]), .LD(n5388), .CP(clk), 
        .Q(Term11[116]) );
  FDS2L \Term11_reg[115]  ( .CR(1'b1), .D(Term1[115]), .LD(n5388), .CP(clk), 
        .Q(Term11[115]) );
  FDS2L \Term11_reg[114]  ( .CR(1'b1), .D(Term1[114]), .LD(n5388), .CP(clk), 
        .Q(Term11[114]) );
  FDS2L \Term11_reg[113]  ( .CR(1'b1), .D(Term1[113]), .LD(n5388), .CP(clk), 
        .Q(Term11[113]) );
  FDS2L \Term11_reg[112]  ( .CR(1'b1), .D(Term1[112]), .LD(n5388), .CP(clk), 
        .Q(Term11[112]) );
  FDS2L \Log_reg[29]  ( .CR(1'b1), .D(IntegerBits[6]), .LD(n5388), .CP(clk), 
        .Q(Log[29]) );
  FDS2L \Log_reg[28]  ( .CR(1'b1), .D(IntegerBits[5]), .LD(n5388), .CP(clk), 
        .Q(Log[28]) );
  FDS2L \Log_reg[27]  ( .CR(1'b1), .D(IntegerBits[4]), .LD(n5388), .CP(clk), 
        .Q(Log[27]) );
  FDS2L \Log_reg[26]  ( .CR(1'b1), .D(IntegerBits[3]), .LD(n5388), .CP(clk), 
        .Q(Log[26]) );
  FDS2L \Log_reg[25]  ( .CR(1'b1), .D(IntegerBits[2]), .LD(n5388), .CP(clk), 
        .Q(Log[25]) );
  FDS2L \Log_reg[24]  ( .CR(1'b1), .D(IntegerBits[1]), .LD(n5388), .CP(clk), 
        .Q(Log[24]) );
  FDS2L \Log_reg[23]  ( .CR(1'b1), .D(IntegerBits[0]), .LD(n5388), .CP(clk), 
        .Q(Log[23]) );
  FDS2L \Log_reg[22]  ( .CR(1'b1), .D(LogPipe[22]), .LD(n5388), .CP(clk), .Q(
        Log[22]) );
  FDS2L \Log_reg[21]  ( .CR(1'b1), .D(LogPipe[21]), .LD(n5388), .CP(clk), .Q(
        Log[21]) );
  FDS2L \Log_reg[20]  ( .CR(1'b1), .D(LogPipe[20]), .LD(n5388), .CP(clk), .Q(
        Log[20]) );
  FDS2L \Log_reg[19]  ( .CR(1'b1), .D(LogPipe[19]), .LD(n5388), .CP(clk), .Q(
        Log[19]) );
  FDS2L \Log_reg[18]  ( .CR(1'b1), .D(LogPipe[18]), .LD(n5388), .CP(clk), .Q(
        Log[18]) );
  FDS2L \Log_reg[17]  ( .CR(1'b1), .D(LogPipe[17]), .LD(n5388), .CP(clk), .Q(
        Log[17]) );
  FDS2L \Log_reg[16]  ( .CR(1'b1), .D(LogPipe[16]), .LD(n5388), .CP(clk), .Q(
        Log[16]) );
  FDS2L \Log_reg[15]  ( .CR(1'b1), .D(LogPipe[15]), .LD(n5388), .CP(clk), .Q(
        Log[15]) );
  FDS2L \Log_reg[14]  ( .CR(1'b1), .D(LogPipe[14]), .LD(n5388), .CP(clk), .Q(
        Log[14]) );
  FDS2L \Log_reg[13]  ( .CR(1'b1), .D(LogPipe[13]), .LD(n5388), .CP(clk), .Q(
        Log[13]) );
  FDS2L \Log_reg[12]  ( .CR(1'b1), .D(LogPipe[12]), .LD(n5388), .CP(clk), .Q(
        Log[12]) );
  FDS2L \Log_reg[11]  ( .CR(1'b1), .D(LogPipe[11]), .LD(n5388), .CP(clk), .Q(
        Log[11]) );
  FDS2L \Log_reg[10]  ( .CR(1'b1), .D(LogPipe[10]), .LD(n5388), .CP(clk), .Q(
        Log[10]) );
  FDS2L \Log_reg[9]  ( .CR(1'b1), .D(LogPipe[9]), .LD(n5388), .CP(clk), .Q(
        Log[9]) );
  FDS2L \Log_reg[8]  ( .CR(1'b1), .D(LogPipe[8]), .LD(n5388), .CP(clk), .Q(
        Log[8]) );
  FDS2L \Log_reg[7]  ( .CR(1'b1), .D(LogPipe[7]), .LD(n5388), .CP(clk), .Q(
        Log[7]) );
  FDS2L \Log_reg[6]  ( .CR(1'b1), .D(LogPipe[6]), .LD(n5388), .CP(clk), .Q(
        Log[6]) );
  FDS2L \Log_reg[5]  ( .CR(1'b1), .D(LogPipe[5]), .LD(n5388), .CP(clk), .Q(
        Log[5]) );
  FDS2L \Log_reg[4]  ( .CR(1'b1), .D(LogPipe[4]), .LD(n5388), .CP(clk), .Q(
        Log[4]) );
  FDS2L \Log_reg[3]  ( .CR(1'b1), .D(LogPipe[3]), .LD(n5388), .CP(clk), .Q(
        Log[3]) );
  FDS2L \Log_reg[2]  ( .CR(1'b1), .D(LogPipe[2]), .LD(n5388), .CP(clk), .Q(
        Log[2]) );
  FDS2L \Log_reg[1]  ( .CR(1'b1), .D(LogPipe[1]), .LD(n5388), .CP(clk), .Q(
        Log[1]) );
  FDS2L \Log_reg[0]  ( .CR(1'b1), .D(LogPipe[0]), .LD(n5388), .CP(clk), .Q(
        Log[0]) );
  FDS2L \LogPipe_reg[22]  ( .CR(1'b1), .D(FractionBit[22]), .LD(n5388), .CP(
        clk), .Q(LogPipe[22]) );
  FDS2L \LogPipe_reg[21]  ( .CR(1'b1), .D(FractionBit[21]), .LD(n5388), .CP(
        clk), .Q(LogPipe[21]) );
  FDS2L \LogPipe_reg[20]  ( .CR(1'b1), .D(FractionBit[20]), .LD(n5388), .CP(
        clk), .Q(LogPipe[20]) );
  FDS2L \LogPipe_reg[19]  ( .CR(1'b1), .D(FractionBit[19]), .LD(n5388), .CP(
        clk), .Q(LogPipe[19]) );
  FDS2L \LogPipe_reg[18]  ( .CR(1'b1), .D(FractionBit[18]), .LD(n5388), .CP(
        clk), .Q(LogPipe[18]) );
  FDS2L \LogPipe_reg[17]  ( .CR(1'b1), .D(FractionBit[17]), .LD(n5388), .CP(
        clk), .Q(LogPipe[17]) );
  FDS2L \LogPipe_reg[16]  ( .CR(1'b1), .D(FractionBit[16]), .LD(n5388), .CP(
        clk), .Q(LogPipe[16]) );
  FDS2L \LogPipe_reg[15]  ( .CR(1'b1), .D(FractionBit[15]), .LD(n5388), .CP(
        clk), .Q(LogPipe[15]) );
  FDS2L \LogPipe_reg[14]  ( .CR(1'b1), .D(FractionBit[14]), .LD(n5388), .CP(
        clk), .Q(LogPipe[14]) );
  FDS2L \LogPipe_reg[13]  ( .CR(1'b1), .D(FractionBit[13]), .LD(n5388), .CP(
        clk), .Q(LogPipe[13]) );
  FDS2L \LogPipe_reg[12]  ( .CR(1'b1), .D(FractionBit[12]), .LD(n5388), .CP(
        clk), .Q(LogPipe[12]) );
  FDS2L \LogPipe_reg[11]  ( .CR(1'b1), .D(FractionBit[11]), .LD(n5388), .CP(
        clk), .Q(LogPipe[11]) );
  FDS2L \LogPipe_reg[10]  ( .CR(1'b1), .D(FractionBit[10]), .LD(n5388), .CP(
        clk), .Q(LogPipe[10]) );
  FDS2L \LogPipe_reg[9]  ( .CR(1'b1), .D(FractionBit[9]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[9]) );
  FDS2L \LogPipe_reg[8]  ( .CR(1'b1), .D(FractionBit[8]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[8]) );
  FDS2L \LogPipe_reg[7]  ( .CR(1'b1), .D(FractionBit[7]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[7]) );
  FDS2L \LogPipe_reg[6]  ( .CR(1'b1), .D(FractionBit[6]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[6]) );
  FDS2L \LogPipe_reg[5]  ( .CR(1'b1), .D(FractionBit[5]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[5]) );
  FDS2L \LogPipe_reg[4]  ( .CR(1'b1), .D(FractionBit[4]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[4]) );
  FDS2L \LogPipe_reg[3]  ( .CR(1'b1), .D(FractionBit[3]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[3]) );
  FDS2L \LogPipe_reg[2]  ( .CR(1'b1), .D(FractionBit[2]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[2]) );
  FDS2L \LogPipe_reg[1]  ( .CR(1'b1), .D(FractionBit[1]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[1]) );
  FDS2L \LogPipe_reg[0]  ( .CR(1'b1), .D(FractionBit[0]), .LD(n5388), .CP(clk), 
        .Q(LogPipe[0]) );
  FDS2L \LogOut_reg[30]  ( .CR(1'b1), .D(Log[29]), .LD(n5388), .CP(clk), .Q(
        LogOut[30]) );
  FDS2L \LogOut_reg[29]  ( .CR(1'b1), .D(Log[28]), .LD(n5388), .CP(clk), .Q(
        LogOut[29]) );
  FDS2L \LogOut_reg[28]  ( .CR(1'b1), .D(Log[27]), .LD(n5388), .CP(clk), .Q(
        LogOut[28]) );
  FDS2L \LogOut_reg[27]  ( .CR(1'b1), .D(Log[26]), .LD(n5388), .CP(clk), .Q(
        LogOut[27]) );
  FDS2L \LogOut_reg[26]  ( .CR(1'b1), .D(Log[25]), .LD(n5388), .CP(clk), .Q(
        LogOut[26]) );
  FDS2L \LogOut_reg[25]  ( .CR(1'b1), .D(Log[24]), .LD(n5388), .CP(clk), .Q(
        LogOut[25]) );
  FDS2L \LogOut_reg[24]  ( .CR(1'b1), .D(Log[23]), .LD(n5388), .CP(clk), .Q(
        LogOut[24]) );
  FDS2L \LogOut_reg[23]  ( .CR(1'b1), .D(Log[22]), .LD(n5388), .CP(clk), .Q(
        LogOut[23]) );
  FDS2L \LogOut_reg[22]  ( .CR(1'b1), .D(Log[21]), .LD(n5388), .CP(clk), .Q(
        LogOut[22]) );
  FDS2L \LogOut_reg[21]  ( .CR(1'b1), .D(Log[20]), .LD(n5388), .CP(clk), .Q(
        LogOut[21]) );
  FDS2L \LogOut_reg[20]  ( .CR(1'b1), .D(Log[19]), .LD(n5388), .CP(clk), .Q(
        LogOut[20]) );
  FDS2L \LogOut_reg[19]  ( .CR(1'b1), .D(Log[18]), .LD(n5388), .CP(clk), .Q(
        LogOut[19]) );
  FDS2L \LogOut_reg[18]  ( .CR(1'b1), .D(Log[17]), .LD(n5388), .CP(clk), .Q(
        LogOut[18]) );
  FDS2L \LogOut_reg[17]  ( .CR(1'b1), .D(Log[16]), .LD(n5388), .CP(clk), .Q(
        LogOut[17]) );
  FDS2L \LogOut_reg[16]  ( .CR(1'b1), .D(Log[15]), .LD(n5388), .CP(clk), .Q(
        LogOut[16]) );
  FDS2L \LogOut_reg[15]  ( .CR(1'b1), .D(Log[14]), .LD(n5388), .CP(clk), .Q(
        LogOut[15]) );
  FDS2L \LogOut_reg[14]  ( .CR(1'b1), .D(Log[13]), .LD(n5388), .CP(clk), .Q(
        LogOut[14]) );
  FDS2L \LogOut_reg[13]  ( .CR(1'b1), .D(Log[12]), .LD(n5388), .CP(clk), .Q(
        LogOut[13]) );
  FDS2L \LogOut_reg[12]  ( .CR(1'b1), .D(Log[11]), .LD(n5388), .CP(clk), .Q(
        LogOut[12]) );
  FDS2L \LogOut_reg[11]  ( .CR(1'b1), .D(Log[10]), .LD(n5388), .CP(clk), .Q(
        LogOut[11]) );
  FDS2L \LogOut_reg[10]  ( .CR(1'b1), .D(Log[9]), .LD(n5388), .CP(clk), .Q(
        LogOut[10]) );
  FDS2L \LogOut_reg[9]  ( .CR(1'b1), .D(Log[8]), .LD(n5388), .CP(clk), .Q(
        LogOut[9]) );
  FDS2L \LogOut_reg[8]  ( .CR(1'b1), .D(Log[7]), .LD(n5388), .CP(clk), .Q(
        LogOut[8]) );
  FDS2L \LogOut_reg[7]  ( .CR(1'b1), .D(Log[6]), .LD(n5388), .CP(clk), .Q(
        LogOut[7]) );
  FDS2L \LogOut_reg[6]  ( .CR(1'b1), .D(Log[5]), .LD(n5388), .CP(clk), .Q(
        LogOut[6]) );
  FDS2L \LogOut_reg[5]  ( .CR(1'b1), .D(Log[4]), .LD(n5388), .CP(clk), .Q(
        LogOut[5]) );
  FDS2L \LogOut_reg[4]  ( .CR(1'b1), .D(Log[3]), .LD(n5388), .CP(clk), .Q(
        LogOut[4]) );
  FDS2L \LogOut_reg[3]  ( .CR(1'b1), .D(Log[2]), .LD(n5388), .CP(clk), .Q(
        LogOut[3]) );
  FDS2L \LogOut_reg[2]  ( .CR(1'b1), .D(Log[1]), .LD(n5388), .CP(clk), .Q(
        LogOut[2]) );
  FDS2L \LogOut_reg[1]  ( .CR(1'b1), .D(Log[0]), .LD(n5388), .CP(clk), .Q(
        LogOut[1]) );
  FDS2L \LogIn2_reg[39]  ( .CR(1'b1), .D(LogIn[39]), .LD(n5388), .CP(clk), .Q(
        LogIn2[39]) );
  FDS2L \LogIn2_reg[38]  ( .CR(1'b1), .D(LogIn[38]), .LD(n5388), .CP(clk), .Q(
        LogIn2[38]) );
  FDS2L \LogIn2_reg[37]  ( .CR(1'b1), .D(LogIn[37]), .LD(n5388), .CP(clk), .Q(
        LogIn2[37]) );
  FDS2L \LogIn2_reg[36]  ( .CR(1'b1), .D(LogIn[36]), .LD(n5388), .CP(clk), .Q(
        LogIn2[36]) );
  FDS2L \LogIn2_reg[35]  ( .CR(1'b1), .D(LogIn[35]), .LD(n5388), .CP(clk), .Q(
        LogIn2[35]) );
  FDS2L \LogIn2_reg[34]  ( .CR(1'b1), .D(LogIn[34]), .LD(n5388), .CP(clk), .Q(
        LogIn2[34]) );
  FDS2L \LogIn2_reg[33]  ( .CR(1'b1), .D(LogIn[33]), .LD(n5388), .CP(clk), .Q(
        LogIn2[33]) );
  FDS2L \LogIn2_reg[32]  ( .CR(1'b1), .D(LogIn[32]), .LD(n5388), .CP(clk), .Q(
        LogIn2[32]) );
  FDS2L \LogIn2_reg[31]  ( .CR(1'b1), .D(LogIn[31]), .LD(n5388), .CP(clk), .Q(
        LogIn2[31]) );
  FDS2L \LogIn2_reg[30]  ( .CR(1'b1), .D(LogIn[30]), .LD(n5388), .CP(clk), .Q(
        LogIn2[30]) );
  FDS2L \LogIn2_reg[29]  ( .CR(1'b1), .D(LogIn[29]), .LD(n5388), .CP(clk), .Q(
        LogIn2[29]) );
  FDS2L \LogIn2_reg[28]  ( .CR(1'b1), .D(LogIn[28]), .LD(n5388), .CP(clk), .Q(
        LogIn2[28]) );
  FDS2L \LogIn2_reg[27]  ( .CR(1'b1), .D(LogIn[27]), .LD(n5388), .CP(clk), .Q(
        LogIn2[27]) );
  FDS2L \LogIn2_reg[26]  ( .CR(1'b1), .D(LogIn[26]), .LD(n5388), .CP(clk), .Q(
        LogIn2[26]) );
  FDS2L \LogIn2_reg[25]  ( .CR(1'b1), .D(LogIn[25]), .LD(n5388), .CP(clk), .Q(
        LogIn2[25]) );
  FDS2L \LogIn2_reg[24]  ( .CR(1'b1), .D(LogIn[24]), .LD(n5388), .CP(clk), .Q(
        LogIn2[24]) );
  FDS2L \LogIn2_reg[23]  ( .CR(1'b1), .D(LogIn[23]), .LD(n5388), .CP(clk), .Q(
        LogIn2[23]) );
  FDS2L \LogIn2_reg[22]  ( .CR(1'b1), .D(LogIn[22]), .LD(n5388), .CP(clk), .Q(
        LogIn2[22]) );
  FDS2L \LogIn2_reg[21]  ( .CR(1'b1), .D(LogIn[21]), .LD(n5388), .CP(clk), .Q(
        LogIn2[21]) );
  FDS2L \LogIn2_reg[20]  ( .CR(1'b1), .D(LogIn[20]), .LD(n5388), .CP(clk), .Q(
        LogIn2[20]) );
  FDS2L \LogIn2_reg[19]  ( .CR(1'b1), .D(LogIn[19]), .LD(n5388), .CP(clk), .Q(
        LogIn2[19]) );
  FDS2L \LogIn2_reg[18]  ( .CR(1'b1), .D(LogIn[18]), .LD(n5388), .CP(clk), .Q(
        LogIn2[18]) );
  FDS2L \LogIn2_reg[17]  ( .CR(1'b1), .D(LogIn[17]), .LD(n5388), .CP(clk), .Q(
        LogIn2[17]) );
  FDS2L \LogIn2_reg[16]  ( .CR(1'b1), .D(LogIn[16]), .LD(n5388), .CP(clk), .Q(
        LogIn2[16]) );
  FDS2L \LogIn2_reg[15]  ( .CR(1'b1), .D(LogIn[15]), .LD(n5388), .CP(clk), .Q(
        LogIn2[15]) );
  FDS2L \LogIn2_reg[14]  ( .CR(1'b1), .D(LogIn[14]), .LD(n5388), .CP(clk), .Q(
        LogIn2[14]) );
  FDS2L \LogIn2_reg[13]  ( .CR(1'b1), .D(LogIn[13]), .LD(n5388), .CP(clk), .Q(
        LogIn2[13]) );
  FDS2L \LogIn2_reg[12]  ( .CR(1'b1), .D(LogIn[12]), .LD(n5388), .CP(clk), .Q(
        LogIn2[12]) );
  FDS2L \LogIn2_reg[11]  ( .CR(1'b1), .D(LogIn[11]), .LD(n5388), .CP(clk), .Q(
        LogIn2[11]) );
  FDS2L \LogIn2_reg[10]  ( .CR(1'b1), .D(LogIn[10]), .LD(n5388), .CP(clk), .Q(
        LogIn2[10]) );
  FDS2L \LogIn2_reg[9]  ( .CR(1'b1), .D(LogIn[9]), .LD(n5388), .CP(clk), .Q(
        LogIn2[9]) );
  FDS2L \LogIn2_reg[8]  ( .CR(1'b1), .D(LogIn[8]), .LD(n5388), .CP(clk), .Q(
        LogIn2[8]) );
  FDS2L \LogIn2_reg[7]  ( .CR(1'b1), .D(LogIn[7]), .LD(n5388), .CP(clk), .Q(
        LogIn2[7]) );
  FDS2L \LogIn2_reg[6]  ( .CR(1'b1), .D(LogIn[6]), .LD(n5388), .CP(clk), .Q(
        LogIn2[6]) );
  FDS2L \LogIn2_reg[5]  ( .CR(1'b1), .D(LogIn[5]), .LD(n5388), .CP(clk), .Q(
        LogIn2[5]) );
  FDS2L \LogIn2_reg[4]  ( .CR(1'b1), .D(LogIn[4]), .LD(n5388), .CP(clk), .Q(
        LogIn2[4]) );
  FDS2L \LogIn2_reg[3]  ( .CR(1'b1), .D(LogIn[3]), .LD(n5388), .CP(clk), .Q(
        LogIn2[3]) );
  FDS2L \LogIn2_reg[2]  ( .CR(1'b1), .D(LogIn[2]), .LD(n5388), .CP(clk), .Q(
        LogIn2[2]) );
  FDS2L \LogIn2_reg[1]  ( .CR(1'b1), .D(LogIn[1]), .LD(n5388), .CP(clk), .Q(
        LogIn2[1]) );
  FDS2L \LogIn2_reg[0]  ( .CR(1'b1), .D(LogIn[0]), .LD(n5388), .CP(clk), .Q(
        LogIn2[0]) );
  FDS2L \LogInSquare_reg[2]  ( .CR(1'b1), .D(N11), .LD(n5388), .CP(clk), .Q(
        LogInSquare[2]) );
  FDS2L \FractionBit_reg[0]  ( .CR(1'b1), .D(N254), .LD(n5388), .CP(clk), .Q(
        FractionBit[0]) );
  FDS2L \FractionBit_reg[1]  ( .CR(1'b1), .D(N255), .LD(n5388), .CP(clk), .Q(
        FractionBit[1]) );
  FDS2L \IntegerBits_reg[0]  ( .CR(1'b1), .D(N292), .LD(n5388), .CP(clk), .Q(
        IntegerBits[0]) );
  FDS2L \FractionBit_reg[2]  ( .CR(1'b1), .D(N256), .LD(n5388), .CP(clk), .Q(
        FractionBit[2]) );
  FDS2L \LogInSquare_reg[3]  ( .CR(1'b1), .D(N12), .LD(n5388), .CP(clk), .Q(
        LogInSquare[3]) );
  FDS2L \FractionBit_reg[3]  ( .CR(1'b1), .D(N257), .LD(n5388), .CP(clk), .Q(
        FractionBit[3]) );
  FDS2L \IntegerBits_reg[1]  ( .CR(1'b1), .D(N293), .LD(n5388), .CP(clk), .Q(
        IntegerBits[1]) );
  FDS2L \FractionBit_reg[4]  ( .CR(1'b1), .D(N258), .LD(n5388), .CP(clk), .Q(
        FractionBit[4]) );
  FDS2L \LogInSquare_reg[4]  ( .CR(1'b1), .D(N13), .LD(n5388), .CP(clk), .Q(
        LogInSquare[4]) );
  FDS2L \IntegerBits_reg[2]  ( .CR(1'b1), .D(N294), .LD(n5388), .CP(clk), .Q(
        IntegerBits[2]) );
  FDS2L \FractionBit_reg[5]  ( .CR(1'b1), .D(N259), .LD(n5388), .CP(clk), .Q(
        FractionBit[5]) );
  FDS2L \Term3_reg[26]  ( .CR(1'b1), .D(n423), .LD(n5388), .CP(clk), .Q(
        Term3[26]) );
  FDS2L \IntegerBits_reg[3]  ( .CR(1'b1), .D(N295), .LD(n5388), .CP(clk), .Q(
        IntegerBits[3]) );
  FDS2L \FractionBit_reg[6]  ( .CR(1'b1), .D(N260), .LD(n5388), .CP(clk), .Q(
        FractionBit[6]) );
  FDS2L \LogInSquare_reg[5]  ( .CR(1'b1), .D(N14), .LD(n5388), .CP(clk), .Q(
        LogInSquare[5]) );
  FDS2L \IntegerBits_reg[4]  ( .CR(1'b1), .D(N296), .LD(n5388), .CP(clk), .Q(
        IntegerBits[4]) );
  FDS2L \Term3_reg[25]  ( .CR(1'b1), .D(N218), .LD(n5388), .CP(clk), .Q(
        Term3[25]) );
  FDS2L \FractionBit_reg[7]  ( .CR(1'b1), .D(N261), .LD(n5388), .CP(clk), .Q(
        FractionBit[7]) );
  FDS2L \Term3_reg[21]  ( .CR(1'b1), .D(N222), .LD(n5388), .CP(clk), .Q(
        Term3[21]) );
  FDS2L \Term3_reg[20]  ( .CR(1'b1), .D(N223), .LD(n5388), .CP(clk), .Q(
        Term3[20]) );
  FDS2L \Term3_reg[18]  ( .CR(1'b1), .D(N225), .LD(n5388), .CP(clk), .Q(
        Term3[18]) );
  FDS2L \Term3_reg[17]  ( .CR(1'b1), .D(N226), .LD(n5388), .CP(clk), .Q(
        Term3[17]) );
  FDS2L \Term3_reg[19]  ( .CR(1'b1), .D(N224), .LD(n5388), .CP(clk), .Q(
        Term3[19]) );
  FDS2L \IntegerBits_reg[5]  ( .CR(1'b1), .D(N297), .LD(n5388), .CP(clk), .Q(
        IntegerBits[5]) );
  FDS2L \Term3_reg[16]  ( .CR(1'b1), .D(N227), .LD(n5388), .CP(clk), .Q(
        Term3[16]) );
  FDS2L \Term3_reg[15]  ( .CR(1'b1), .D(N228), .LD(n5388), .CP(clk), .Q(
        Term3[15]) );
  FDS2L \FractionBit_reg[8]  ( .CR(1'b1), .D(N262), .LD(n5388), .CP(clk), .Q(
        FractionBit[8]) );
  FDS2L \LogInSquare_reg[6]  ( .CR(1'b1), .D(N15), .LD(n5388), .CP(clk), .Q(
        LogInSquare[6]) );
  FDS2L \Term3_reg[24]  ( .CR(1'b1), .D(N219), .LD(n5388), .CP(clk), .Q(
        Term3[24]) );
  FDS2L \Term3_reg[14]  ( .CR(1'b1), .D(N229), .LD(n5388), .CP(clk), .Q(
        Term3[14]) );
  FDS2L \Term3_reg[22]  ( .CR(1'b1), .D(N221), .LD(n5388), .CP(clk), .Q(
        Term3[22]) );
  FDS2L \FractionBit_reg[9]  ( .CR(1'b1), .D(N263), .LD(n5388), .CP(clk), .Q(
        FractionBit[9]) );
  FDS2L \IntegerBits_reg[6]  ( .CR(1'b1), .D(N298), .LD(n5388), .CP(clk), .Q(
        IntegerBits[6]) );
  FDS2L \FractionBit_reg[10]  ( .CR(1'b1), .D(N264), .LD(n5388), .CP(clk), .Q(
        FractionBit[10]) );
  FDS2L \LogInSquare_reg[7]  ( .CR(1'b1), .D(N16), .LD(n5388), .CP(clk), .Q(
        LogInSquare[7]) );
  FDS2L \FractionBit_reg[11]  ( .CR(1'b1), .D(N265), .LD(n5388), .CP(clk), .Q(
        FractionBit[11]) );
  FDS2L \FractionBit_reg[12]  ( .CR(1'b1), .D(N266), .LD(n5388), .CP(clk), .Q(
        FractionBit[12]) );
  FDS2L \LogInSquare_reg[8]  ( .CR(1'b1), .D(N17), .LD(n5388), .CP(clk), .Q(
        LogInSquare[8]) );
  FDS2L \FractionBit_reg[13]  ( .CR(1'b1), .D(N267), .LD(n5388), .CP(clk), .Q(
        FractionBit[13]) );
  FDS2L \LogInSquare_reg[9]  ( .CR(1'b1), .D(N18), .LD(n5388), .CP(clk), .Q(
        LogInSquare[9]) );
  FDS2L \FractionBit_reg[14]  ( .CR(1'b1), .D(N268), .LD(n5388), .CP(clk), .Q(
        FractionBit[14]) );
  FDS2L \FractionBit_reg[15]  ( .CR(1'b1), .D(N269), .LD(n5388), .CP(clk), .Q(
        FractionBit[15]) );
  FDS2L \LogInSquare_reg[10]  ( .CR(1'b1), .D(N19), .LD(n5388), .CP(clk), .Q(
        LogInSquare[10]) );
  FDS2L \FractionBit_reg[16]  ( .CR(1'b1), .D(N270), .LD(n5388), .CP(clk), .Q(
        FractionBit[16]) );
  FDS2L \FractionBit_reg[17]  ( .CR(1'b1), .D(N271), .LD(n5388), .CP(clk), .Q(
        FractionBit[17]) );
  FDS2L \LogInSquare_reg[11]  ( .CR(1'b1), .D(N20), .LD(n5388), .CP(clk), .Q(
        LogInSquare[11]) );
  FDS2L \FractionBit_reg[18]  ( .CR(1'b1), .D(N272), .LD(n5388), .CP(clk), .Q(
        FractionBit[18]) );
  FDS2L \FractionBit_reg[19]  ( .CR(1'b1), .D(N273), .LD(n5388), .CP(clk), .Q(
        FractionBit[19]) );
  FDS2L \LogInSquare_reg[12]  ( .CR(1'b1), .D(N21), .LD(n5388), .CP(clk), .Q(
        LogInSquare[12]) );
  FDS2L \FractionBit_reg[20]  ( .CR(1'b1), .D(N274), .LD(n5388), .CP(clk), .Q(
        FractionBit[20]) );
  FDS2L \FractionBit_reg[21]  ( .CR(1'b1), .D(N275), .LD(n5388), .CP(clk), .Q(
        FractionBit[21]) );
  FDS2L \LogInSquare_reg[13]  ( .CR(1'b1), .D(N22), .LD(n5388), .CP(clk), .Q(
        LogInSquare[13]) );
  FDS2L \FractionBit_reg[22]  ( .CR(1'b1), .D(N276), .LD(n5388), .CP(clk), .Q(
        FractionBit[22]) );
  FDS2L \FractionBit_reg[23]  ( .CR(1'b1), .D(N277), .LD(n5388), .CP(clk), .Q(
        FractionBit[23]) );
  FDS2L \LogInSquare_reg[14]  ( .CR(1'b1), .D(N23), .LD(n5388), .CP(clk), .Q(
        LogInSquare[14]) );
  FDS2L \LogInSquare_reg[15]  ( .CR(1'b1), .D(N24), .LD(n5388), .CP(clk), .Q(
        LogInSquare[15]) );
  FDS2L \LogInSquare_reg[16]  ( .CR(1'b1), .D(N25), .LD(n5388), .CP(clk), .Q(
        LogInSquare[16]) );
  FDS2L \LogInSquare_reg[17]  ( .CR(1'b1), .D(N26), .LD(n5388), .CP(clk), .Q(
        LogInSquare[17]) );
  FDS2L \LogInSquare_reg[18]  ( .CR(1'b1), .D(N27), .LD(n5388), .CP(clk), .Q(
        LogInSquare[18]) );
  FDS2L \LogInSquare_reg[19]  ( .CR(1'b1), .D(N28), .LD(n5388), .CP(clk), .Q(
        LogInSquare[19]) );
  FDS2L \LogInSquare_reg[20]  ( .CR(1'b1), .D(N29), .LD(n5388), .CP(clk), .Q(
        LogInSquare[20]) );
  FDS2L \LogInSquare_reg[21]  ( .CR(1'b1), .D(N30), .LD(n5388), .CP(clk), .Q(
        LogInSquare[21]) );
  FDS2L \LogInSquare_reg[22]  ( .CR(1'b1), .D(N31), .LD(n5388), .CP(clk), .Q(
        LogInSquare[22]) );
  FDS2L \LogInSquare_reg[23]  ( .CR(1'b1), .D(N32), .LD(n5388), .CP(clk), .Q(
        LogInSquare[23]) );
  FDS2L \LogInSquare_reg[24]  ( .CR(1'b1), .D(N33), .LD(n5388), .CP(clk), .Q(
        LogInSquare[24]) );
  FDS2L \LogInSquare_reg[25]  ( .CR(1'b1), .D(N34), .LD(n5388), .CP(clk), .Q(
        LogInSquare[25]) );
  FDS2L \LogInSquare_reg[26]  ( .CR(1'b1), .D(N35), .LD(n5388), .CP(clk), .Q(
        LogInSquare[26]) );
  FDS2L \LogInSquare_reg[27]  ( .CR(1'b1), .D(N36), .LD(n5388), .CP(clk), .Q(
        LogInSquare[27]) );
  FDS2L \LogInSquare_reg[28]  ( .CR(1'b1), .D(N37), .LD(n5388), .CP(clk), .Q(
        LogInSquare[28]) );
  FDS2L \LogInSquare_reg[29]  ( .CR(1'b1), .D(N38), .LD(n5388), .CP(clk), .Q(
        LogInSquare[29]) );
  FDS2L \LogInSquare_reg[30]  ( .CR(1'b1), .D(N39), .LD(n5388), .CP(clk), .Q(
        LogInSquare[30]) );
  FDS2L \LogInSquare_reg[31]  ( .CR(1'b1), .D(N40), .LD(n5388), .CP(clk), .Q(
        LogInSquare[31]) );
  FDS2L \LogInSquare_reg[32]  ( .CR(1'b1), .D(N41), .LD(n5388), .CP(clk), .Q(
        LogInSquare[32]) );
  FDS2L \LogInSquare_reg[33]  ( .CR(1'b1), .D(N42), .LD(n5388), .CP(clk), .Q(
        LogInSquare[33]) );
  FDS2L \LogInSquare_reg[34]  ( .CR(1'b1), .D(N43), .LD(n5388), .CP(clk), .Q(
        LogInSquare[34]) );
  FDS2L \LogInSquare_reg[35]  ( .CR(1'b1), .D(N44), .LD(n5388), .CP(clk), .Q(
        LogInSquare[35]) );
  FDS2L \LogInSquare_reg[36]  ( .CR(1'b1), .D(N45), .LD(n5388), .CP(clk), .Q(
        LogInSquare[36]) );
  FDS2L \LogInSquare_reg[37]  ( .CR(1'b1), .D(N46), .LD(n5388), .CP(clk), .Q(
        LogInSquare[37]) );
  FDS2L \LogInSquare_reg[38]  ( .CR(1'b1), .D(N47), .LD(n5388), .CP(clk), .Q(
        LogInSquare[38]) );
  FDS2L \LogInSquare_reg[39]  ( .CR(1'b1), .D(N48), .LD(n5388), .CP(clk), .Q(
        LogInSquare[39]) );
  FDS2L \LogInSquare_reg[40]  ( .CR(1'b1), .D(N49), .LD(n5388), .CP(clk), .Q(
        LogInSquare[40]) );
  FDS2L \LogInSquare_reg[41]  ( .CR(1'b1), .D(N50), .LD(n5388), .CP(clk), .Q(
        LogInSquare[41]) );
  FDS2L \LogInSquare_reg[42]  ( .CR(1'b1), .D(N51), .LD(n5388), .CP(clk), .Q(
        LogInSquare[42]) );
  FDS2L \Term2_reg[38]  ( .CR(1'b1), .D(N187), .LD(n5388), .CP(clk), .Q(
        Term2[38]) );
  FDS2L \Term2_reg[39]  ( .CR(1'b1), .D(N188), .LD(n5388), .CP(clk), .Q(
        Term2[39]) );
  FDS2L \Term2_reg[42]  ( .CR(1'b1), .D(N191), .LD(n5388), .CP(clk), .Q(
        Term2[42]) );
  FDS2L \LogInSquare_reg[43]  ( .CR(1'b1), .D(N52), .LD(n5388), .CP(clk), .Q(
        LogInSquare[43]) );
  FDS2L \Term2_reg[40]  ( .CR(1'b1), .D(N189), .LD(n5388), .CP(clk), .Q(
        Term2[40]) );
  FDS2L \Term2_reg[46]  ( .CR(1'b1), .D(N195), .LD(n5388), .CP(clk), .Q(
        Term2[46]) );
  FDS2L \Term2_reg[43]  ( .CR(1'b1), .D(N192), .LD(n5388), .CP(clk), .Q(
        Term2[43]) );
  FDS2L \Term2_reg[41]  ( .CR(1'b1), .D(N190), .LD(n5388), .CP(clk), .Q(
        Term2[41]) );
  FDS2L \Term2_reg[47]  ( .CR(1'b1), .D(N196), .LD(n5388), .CP(clk), .Q(
        Term2[47]) );
  FDS2L \Term2_reg[44]  ( .CR(1'b1), .D(N193), .LD(n5388), .CP(clk), .Q(
        Term2[44]) );
  FDS2L \LogInSquare_reg[44]  ( .CR(1'b1), .D(N53), .LD(n5388), .CP(clk), .Q(
        LogInSquare[44]) );
  FDS2L \Term2_reg[50]  ( .CR(1'b1), .D(N199), .LD(n5388), .CP(clk), .Q(
        Term2[50]) );
  FDS2L \Term2_reg[51]  ( .CR(1'b1), .D(N200), .LD(n5388), .CP(clk), .Q(
        Term2[51]) );
  FDS2L \Term2_reg[45]  ( .CR(1'b1), .D(N194), .LD(n5388), .CP(clk), .Q(
        Term2[45]) );
  FDS2L \Term2_reg[48]  ( .CR(1'b1), .D(N197), .LD(n5388), .CP(clk), .Q(
        Term2[48]) );
  FDS2L \LogInSquare_reg[45]  ( .CR(1'b1), .D(N54), .LD(n5388), .CP(clk), .Q(
        LogInSquare[45]) );
  FDS2L \Term2_reg[49]  ( .CR(1'b1), .D(N198), .LD(n5388), .CP(clk), .Q(
        Term2[49]) );
  FDS2L \Term2_reg[54]  ( .CR(1'b1), .D(N203), .LD(n5388), .CP(clk), .Q(
        Term2[54]) );
  FDS2L \Term2_reg[52]  ( .CR(1'b1), .D(N201), .LD(n5388), .CP(clk), .Q(
        Term2[52]) );
  FDS2L \Term2_reg[53]  ( .CR(1'b1), .D(N202), .LD(n5388), .CP(clk), .Q(
        Term2[53]) );
  FDS2L \LogInSquare_reg[46]  ( .CR(1'b1), .D(N55), .LD(n5388), .CP(clk), .Q(
        LogInSquare[46]) );
  FDS2L \Term2_reg[55]  ( .CR(1'b1), .D(N204), .LD(n5388), .CP(clk), .Q(
        Term2[55]) );
  FDS2L \Term2_reg[58]  ( .CR(1'b1), .D(N207), .LD(n5388), .CP(clk), .Q(
        Term2[58]) );
  FDS2L \Term2_reg[56]  ( .CR(1'b1), .D(N205), .LD(n5388), .CP(clk), .Q(
        Term2[56]) );
  FDS2L \Term2_reg[62]  ( .CR(1'b1), .D(N211), .LD(n5388), .CP(clk), .Q(
        Term2[62]) );
  FDS2L \LogInSquare_reg[47]  ( .CR(1'b1), .D(N56), .LD(n5388), .CP(clk), .Q(
        LogInSquare[47]) );
  FDS2L \Term2_reg[59]  ( .CR(1'b1), .D(N208), .LD(n5388), .CP(clk), .Q(
        Term2[59]) );
  FDS2L \Term2_reg[57]  ( .CR(1'b1), .D(N206), .LD(n5388), .CP(clk), .Q(
        Term2[57]) );
  FDS2L \LogInSquare_reg[48]  ( .CR(1'b1), .D(N57), .LD(n5388), .CP(clk), .Q(
        LogInSquare[48]) );
  FDS2L \Term2_reg[60]  ( .CR(1'b1), .D(N209), .LD(n5388), .CP(clk), .Q(
        Term2[60]) );
  FDS2L \Term1_reg[106]  ( .CR(1'b1), .D(N152), .LD(n5388), .CP(clk), .Q(
        Term1[106]) );
  FDS2L \Term1_reg[90]  ( .CR(1'b1), .D(N136), .LD(n5388), .CP(clk), .Q(N231)
         );
  FDS2L \Term1_reg[98]  ( .CR(1'b1), .D(N144), .LD(n5388), .CP(clk), .Q(N239)
         );
  FDS2L \Term2_reg[63]  ( .CR(1'b1), .D(N212), .LD(n5388), .CP(clk), .Q(
        Term2[63]) );
  FDS2L \Term2_reg[66]  ( .CR(1'b1), .D(N215), .LD(n5388), .CP(clk), .Q(
        Term2[66]) );
  FDS2L \Term1_reg[89]  ( .CR(1'b1), .D(N135), .LD(n5388), .CP(clk), .Q(N230)
         );
  FDS2L \Term2_reg[64]  ( .CR(1'b1), .D(N213), .LD(n5388), .CP(clk), .Q(
        Term2[64]) );
  FDS2L \Term1_reg[114]  ( .CR(1'b1), .D(N160), .LD(n5388), .CP(clk), .Q(
        Term1[114]) );
  FDS2L \Term1_reg[115]  ( .CR(1'b1), .D(N161), .LD(n5388), .CP(clk), .Q(
        Term1[115]) );
  FDS2L \Term1_reg[110]  ( .CR(1'b1), .D(N156), .LD(n5388), .CP(clk), .Q(
        Term1[110]) );
  FDS2L \Term1_reg[107]  ( .CR(1'b1), .D(N153), .LD(n5388), .CP(clk), .Q(
        Term1[107]) );
  FDS2L \Term1_reg[94]  ( .CR(1'b1), .D(N140), .LD(n5388), .CP(clk), .Q(N235)
         );
  FDS2L \Term1_reg[91]  ( .CR(1'b1), .D(N137), .LD(n5388), .CP(clk), .Q(N232)
         );
  FDS2L \Term1_reg[99]  ( .CR(1'b1), .D(N145), .LD(n5388), .CP(clk), .Q(N240)
         );
  FDS2L \LogInSquare_reg[49]  ( .CR(1'b1), .D(N58), .LD(n5388), .CP(clk), .Q(
        LogInSquare[49]) );
  FDS2L \Term2_reg[61]  ( .CR(1'b1), .D(N210), .LD(n5388), .CP(clk), .Q(
        Term2[61]) );
  FDS2L \Term1_reg[102]  ( .CR(1'b1), .D(N148), .LD(n5388), .CP(clk), .Q(
        Term1[102]) );
  FDS2L \Term2_reg[67]  ( .CR(1'b1), .D(N216), .LD(n5388), .CP(clk), .Q(
        Term2[67]) );
  FDS2L \Term2_reg[65]  ( .CR(1'b1), .D(N214), .LD(n5388), .CP(clk), .Q(
        Term2[65]) );
  FDS2L \LogInSquare_reg[50]  ( .CR(1'b1), .D(N59), .LD(n5388), .CP(clk), .Q(
        LogInSquare[50]) );
  FDS2L \Term1_reg[116]  ( .CR(1'b1), .D(N162), .LD(n5388), .CP(clk), .Q(
        Term1[116]) );
  FDS2L \Term1_reg[108]  ( .CR(1'b1), .D(N154), .LD(n5388), .CP(clk), .Q(
        Term1[108]) );
  FDS2L \Term1_reg[95]  ( .CR(1'b1), .D(N141), .LD(n5388), .CP(clk), .Q(N236)
         );
  FDS2L \Term1_reg[92]  ( .CR(1'b1), .D(N138), .LD(n5388), .CP(clk), .Q(N233)
         );
  FDS2L \Term1_reg[100]  ( .CR(1'b1), .D(N146), .LD(n5388), .CP(clk), .Q(N241)
         );
  FDS2L \Term1_reg[103]  ( .CR(1'b1), .D(N149), .LD(n5388), .CP(clk), .Q(
        Term1[103]) );
  FDS2L \Term1_reg[117]  ( .CR(1'b1), .D(N163), .LD(n5388), .CP(clk), .Q(
        Term1[117]) );
  FDS2L \LogInSquare_reg[51]  ( .CR(1'b1), .D(N60), .LD(n5388), .CP(clk), .Q(
        LogInSquare[51]) );
  FDS2L \Term1_reg[101]  ( .CR(1'b1), .D(N147), .LD(n5388), .CP(clk), .Q(N242)
         );
  FDS2L \Term1_reg[109]  ( .CR(1'b1), .D(N155), .LD(n5388), .CP(clk), .Q(
        Term1[109]) );
  FDS2L \Term1_reg[93]  ( .CR(1'b1), .D(N139), .LD(n5388), .CP(clk), .Q(N234)
         );
  FDS2L \Term1_reg[118]  ( .CR(1'b1), .D(N164), .LD(n5388), .CP(clk), .Q(
        Term1[118]) );
  FDS2L \Term1_reg[112]  ( .CR(1'b1), .D(N158), .LD(n5388), .CP(clk), .Q(
        Term1[112]) );
  FDS2L \Term1_reg[96]  ( .CR(1'b1), .D(N142), .LD(n5388), .CP(clk), .Q(N237)
         );
  FDS2L \Term1_reg[104]  ( .CR(1'b1), .D(N150), .LD(n5388), .CP(clk), .Q(
        Term1[104]) );
  FDS2L \LogInSquare_reg[54]  ( .CR(1'b1), .D(N63), .LD(n5388), .CP(clk), .Q(
        LogInSquare[54]) );
  FDS2L \LogInSquare_reg[52]  ( .CR(1'b1), .D(N61), .LD(n5388), .CP(clk), .Q(
        LogInSquare[52]) );
  FDS2L \Term1_reg[113]  ( .CR(1'b1), .D(N159), .LD(n5388), .CP(clk), .Q(
        Term1[113]) );
  FDS2L \Term1_reg[97]  ( .CR(1'b1), .D(N143), .LD(n5388), .CP(clk), .Q(N238)
         );
  FDS2L \LogInSquare_reg[58]  ( .CR(1'b1), .D(N67), .LD(n5388), .CP(clk), .Q(
        LogInSquare[58]) );
  FDS2L \Term1_reg[105]  ( .CR(1'b1), .D(N151), .LD(n5388), .CP(clk), .Q(
        Term1[105]) );
  FDS2L \LogInSquare_reg[53]  ( .CR(1'b1), .D(N62), .LD(n5388), .CP(clk), .Q(
        LogInSquare[53]) );
  FDS2L \LogInSquare_reg[55]  ( .CR(1'b1), .D(N64), .LD(n5388), .CP(clk), .Q(
        LogInSquare[55]) );
  FDS2L \LogInSquare_reg[67]  ( .CR(1'b1), .D(N76), .LD(n5388), .CP(clk), .Q(
        LogInSquare[67]) );
  FDS2L \LogInSquare_reg[71]  ( .CR(1'b1), .D(N80), .LD(n5388), .CP(clk), .Q(
        LogInSquare[71]) );
  FDS2L \LogInSquare_reg[62]  ( .CR(1'b1), .D(N71), .LD(n5388), .CP(clk), .Q(
        LogInSquare[62]) );
  FDS2L \LogInSquare_reg[70]  ( .CR(1'b1), .D(N79), .LD(n5388), .CP(clk), .Q(
        LogInSquare[70]) );
  FDS2L \LogInSquare_reg[66]  ( .CR(1'b1), .D(N75), .LD(n5388), .CP(clk), .Q(
        LogInSquare[66]) );
  FDS2L \LogInSquare_reg[63]  ( .CR(1'b1), .D(N72), .LD(n5388), .CP(clk), .Q(
        LogInSquare[63]) );
  FDS2L \LogInSquare_reg[59]  ( .CR(1'b1), .D(N68), .LD(n5388), .CP(clk), .Q(
        LogInSquare[59]) );
  FDS2L \LogInSquare_reg[82]  ( .CR(1'b1), .D(N91), .LD(n5388), .CP(clk), .Q(
        LogInSquare[82]) );
  FDS2L \LogInSquare_reg[79]  ( .CR(1'b1), .D(N88), .LD(n5388), .CP(clk), .Q(
        LogInSquare[79]) );
  FDS2L \LogInSquare_reg[78]  ( .CR(1'b1), .D(N87), .LD(n5388), .CP(clk), .Q(
        LogInSquare[78]) );
  FDS2L \LogInSquare_reg[75]  ( .CR(1'b1), .D(N84), .LD(n5388), .CP(clk), .Q(
        LogInSquare[75]) );
  FDS2L \LogInSquare_reg[74]  ( .CR(1'b1), .D(N83), .LD(n5388), .CP(clk), .Q(
        LogInSquare[74]) );
  FDS2L \LogInSquare_reg[60]  ( .CR(1'b1), .D(N69), .LD(n5388), .CP(clk), .Q(
        LogInSquare[60]) );
  FDS2L \LogInSquare_reg[76]  ( .CR(1'b1), .D(N85), .LD(n5388), .CP(clk), .Q(
        LogInSquare[76]) );
  FDS2L \LogInSquare_reg[56]  ( .CR(1'b1), .D(N65), .LD(n5388), .CP(clk), .Q(
        LogInSquare[56]) );
  FDS2L \LogInSquare_reg[72]  ( .CR(1'b1), .D(N81), .LD(n5388), .CP(clk), .Q(
        LogInSquare[72]) );
  FDS2L \LogInSquare_reg[89]  ( .CR(1'b1), .D(N98), .LD(n5388), .CP(clk), .Q(
        LogInSquare[89]) );
  FDS2L \LogInSquare_reg[68]  ( .CR(1'b1), .D(N77), .LD(n5388), .CP(clk), .Q(
        LogInSquare[68]) );
  FDS2L \LogInSquare_reg[80]  ( .CR(1'b1), .D(N89), .LD(n5388), .CP(clk), .Q(
        LogInSquare[80]) );
  FDS2L \LogInSquare_reg[64]  ( .CR(1'b1), .D(N73), .LD(n5388), .CP(clk), .Q(
        LogInSquare[64]) );
  FDS2L \LogInSquare_reg[95]  ( .CR(1'b1), .D(N104), .LD(n5388), .CP(clk), .Q(
        LogInSquare[95]) );
  FDS2L \LogInSquare_reg[57]  ( .CR(1'b1), .D(N66), .LD(n5388), .CP(clk), .Q(
        LogInSquare[57]) );
  FDS2L \LogInSquare_reg[88]  ( .CR(1'b1), .D(N97), .LD(n5367), .CP(clk), .Q(
        LogInSquare[88]) );
  B5I U17007 ( .A(n817), .Z(n818) );
  B5I U17008 ( .A(n795), .Z(n796) );
  B5I U17009 ( .A(n815), .Z(n816) );
  MUX21LP U17010 ( .A(LogInSquare[65]), .B(N74), .S(n5365), .Z(n815) );
  MUX21LP U17011 ( .A(LogInSquare[77]), .B(N86), .S(n5366), .Z(n813) );
  NR3 U17012 ( .A(n4352), .B(n784), .C(n4267), .Z(n3735) );
  NR3 U17013 ( .A(n4262), .B(n4339), .C(n782), .Z(n3988) );
  NR2 U17014 ( .A(n4336), .B(n783), .Z(n4118) );
  NR3 U17015 ( .A(n4335), .B(n788), .C(n4265), .Z(n3839) );
  NR2 U17016 ( .A(n4290), .B(n789), .Z(n3838) );
  NR2 U17017 ( .A(n4266), .B(n787), .Z(n3780) );
  NR2 U17018 ( .A(n4351), .B(n785), .Z(n3687) );
  NR2 U17019 ( .A(n4265), .B(n786), .Z(n3802) );
  NR3 U17020 ( .A(n790), .B(n4337), .C(n4292), .Z(n3927) );
  IVP U17021 ( .A(n797), .Z(n798) );
  IVP U17022 ( .A(n799), .Z(n800) );
  IVP U17023 ( .A(n801), .Z(n802) );
  IVP U17024 ( .A(n803), .Z(n804) );
  IVP U17025 ( .A(n813), .Z(n814) );
  IVP U17026 ( .A(n825), .Z(n826) );
  MUX21L U17027 ( .A(LogInSquare[61]), .B(N70), .S(n5365), .Z(n825) );
  AN3 U17028 ( .A(n4203), .B(n4212), .C(n400), .Z(n354) );
  AN3 U17029 ( .A(n4203), .B(n4212), .C(n402), .Z(n355) );
  AN3 U17030 ( .A(n4202), .B(n4211), .C(n403), .Z(n356) );
  AN3 U17031 ( .A(n4205), .B(n4211), .C(n407), .Z(n357) );
  AN3 U17032 ( .A(n4205), .B(n4211), .C(n408), .Z(n358) );
  AN3 U17033 ( .A(n4205), .B(n4215), .C(n409), .Z(n359) );
  AN3 U17034 ( .A(n4205), .B(n4215), .C(n410), .Z(n360) );
  AN3 U17035 ( .A(n4205), .B(n4214), .C(n411), .Z(n361) );
  AN2P U17036 ( .A(n2985), .B(n2984), .Z(n362) );
  AN2P U17037 ( .A(n2859), .B(n2858), .Z(n363) );
  AN2P U17038 ( .A(n3123), .B(n3122), .Z(n364) );
  AN2P U17039 ( .A(n2429), .B(n4528), .Z(n365) );
  AN2P U17040 ( .A(n2898), .B(n2897), .Z(n366) );
  MUX21H U17041 ( .A(n3014), .B(n3013), .S(n5239), .Z(n367) );
  MUX21H U17042 ( .A(n2518), .B(n4477), .S(n4904), .Z(n368) );
  MUX21H U17043 ( .A(n4632), .B(n2316), .S(n5261), .Z(n369) );
  AN2P U17044 ( .A(n2329), .B(n2328), .Z(n370) );
  AN2P U17045 ( .A(n2162), .B(n2161), .Z(n371) );
  AN2P U17046 ( .A(n2520), .B(n2519), .Z(n372) );
  AN2P U17047 ( .A(n2654), .B(n2653), .Z(n373) );
  MUX21H U17048 ( .A(n3093), .B(n3092), .S(n4581), .Z(n374) );
  AN3 U17049 ( .A(n2884), .B(n2883), .C(n2882), .Z(n375) );
  AN3 U17050 ( .A(n3487), .B(n3486), .C(n3485), .Z(n376) );
  AN2P U17051 ( .A(n3559), .B(n3558), .Z(n377) );
  AN2P U17052 ( .A(n2302), .B(n2301), .Z(n378) );
  AN2P U17053 ( .A(n2354), .B(n4534), .Z(n379) );
  AN2P U17054 ( .A(n2276), .B(n2275), .Z(n380) );
  MUX21H U17055 ( .A(n4874), .B(n2313), .S(n4631), .Z(n381) );
  AN3 U17056 ( .A(n3070), .B(n3069), .C(n3068), .Z(n382) );
  AN2P U17057 ( .A(n4534), .B(n4878), .Z(n383) );
  AN3 U17058 ( .A(n4266), .B(n3758), .C(n3757), .Z(n384) );
  AN2P U17059 ( .A(n3029), .B(n3028), .Z(n385) );
  MUX21H U17060 ( .A(n4817), .B(n3044), .S(n4550), .Z(n386) );
  AN2P U17061 ( .A(n3633), .B(n3632), .Z(n387) );
  AN3 U17062 ( .A(n4204), .B(n4214), .C(n1097), .Z(n388) );
  AN3 U17063 ( .A(n4203), .B(n4213), .C(n1094), .Z(n389) );
  AN2P U17064 ( .A(n3581), .B(n3580), .Z(n390) );
  MUX21H U17065 ( .A(n3498), .B(n3497), .S(n5245), .Z(n391) );
  AN3 U17066 ( .A(n4206), .B(n4217), .C(n1509), .Z(n392) );
  AN2P U17067 ( .A(n3560), .B(n4924), .Z(n393) );
  AN3 U17068 ( .A(n4206), .B(n4217), .C(n1504), .Z(n394) );
  AN3 U17069 ( .A(n4203), .B(n4213), .C(n1092), .Z(n395) );
  MUX21H U17070 ( .A(n4590), .B(n4783), .S(n5243), .Z(n396) );
  AN3 U17071 ( .A(n4206), .B(n4211), .C(n1501), .Z(n397) );
  MUX21H U17072 ( .A(n4591), .B(n3450), .S(n4919), .Z(n398) );
  MUX21H U17073 ( .A(n3562), .B(n3561), .S(n5248), .Z(n399) );
  AN4P U17074 ( .A(n1090), .B(n4233), .C(n4280), .D(n4316), .Z(n400) );
  MUX21H U17075 ( .A(n5119), .B(n4570), .S(n4921), .Z(n401) );
  AN4P U17076 ( .A(n1089), .B(n4231), .C(n4283), .D(n4317), .Z(n402) );
  AN4P U17077 ( .A(n1088), .B(n4232), .C(n4280), .D(n4317), .Z(n403) );
  AN4P U17078 ( .A(n4338), .B(n1498), .C(n4237), .D(n4281), .Z(n404) );
  AN3 U17079 ( .A(n4205), .B(n4216), .C(n1496), .Z(n405) );
  AN3 U17080 ( .A(n4205), .B(n4216), .C(n1494), .Z(n406) );
  AN4P U17081 ( .A(n1491), .B(n4236), .C(n4287), .D(n4319), .Z(n407) );
  AN4P U17082 ( .A(n1490), .B(n4235), .C(n4281), .D(n4319), .Z(n408) );
  AN4P U17083 ( .A(n1489), .B(n4235), .C(n4283), .D(n4319), .Z(n409) );
  AN4P U17084 ( .A(n1488), .B(n4234), .C(n4281), .D(n4318), .Z(n410) );
  AN4P U17085 ( .A(n1487), .B(n4234), .C(n4284), .D(n4318), .Z(n411) );
  AN2P U17086 ( .A(Term3[14]), .B(Term1[102]), .Z(n412) );
  AN4P U17087 ( .A(n4010), .B(n4009), .C(n4008), .D(n4007), .Z(n413) );
  AN2P U17088 ( .A(n2335), .B(n2334), .Z(n414) );
  AN2P U17089 ( .A(n3593), .B(n3592), .Z(n415) );
  AN4P U17090 ( .A(n4020), .B(n4019), .C(n4018), .D(n4017), .Z(n416) );
  MUX21H U17091 ( .A(n4926), .B(n4576), .S(n5249), .Z(n417) );
  AN2P U17092 ( .A(n2497), .B(n2496), .Z(n418) );
  MUX21H U17093 ( .A(n2660), .B(n4970), .S(n4625), .Z(n419) );
  AN3 U17094 ( .A(n2338), .B(n2337), .C(n2336), .Z(n420) );
  MUX21H U17095 ( .A(n2348), .B(n2347), .S(n5262), .Z(n421) );
  AN4P U17096 ( .A(n845), .B(n4245), .C(n4286), .D(n4327), .Z(n422) );
  AN3 U17097 ( .A(n4202), .B(n4211), .C(n827), .Z(n423) );
  IVP U17427 ( .A(n819), .Z(n820) );
  MUX21LP U17428 ( .A(LogInSquare[69]), .B(N78), .S(n5365), .Z(n819) );
  MUX21LP U17429 ( .A(LogInSquare[81]), .B(N90), .S(n5366), .Z(n817) );
  MUX21LP U17430 ( .A(LogInSquare[93]), .B(N102), .S(n5367), .Z(n801) );
  MUX21LP U17431 ( .A(LogInSquare[94]), .B(N103), .S(n5367), .Z(n803) );
  MUX21LP U17432 ( .A(LogInSquare[91]), .B(N100), .S(n5367), .Z(n797) );
  MUX21LP U17433 ( .A(LogInSquare[92]), .B(N101), .S(n5367), .Z(n799) );
  IVP U17434 ( .A(n805), .Z(n806) );
  MUX21LP U17435 ( .A(LogInSquare[73]), .B(N82), .S(n5366), .Z(n805) );
  MUX21LP U17436 ( .A(LogInSquare[90]), .B(N99), .S(n5367), .Z(n795) );
  ND2 U17437 ( .A(n2957), .B(n2956), .Z(n1979) );
  ND2 U17438 ( .A(n5286), .B(n4550), .Z(n2956) );
  EN U17439 ( .A(n4900), .B(n4548), .Z(n2957) );
  NR2 U17440 ( .A(n5283), .B(n4932), .Z(n2857) );
  EO U17441 ( .A(n5225), .B(n4610), .Z(n2021) );
  EN U17442 ( .A(n4903), .B(n4560), .Z(n2756) );
  ND2 U17443 ( .A(n5278), .B(n4560), .Z(n2755) );
  ND2 U17444 ( .A(n2028), .B(n2027), .Z(n1959) );
  EN U17445 ( .A(n4902), .B(n4628), .Z(n2028) );
  EN U17446 ( .A(n5227), .B(n4628), .Z(n2027) );
  ND2 U17447 ( .A(n2267), .B(n2266), .Z(n1965) );
  ND2 U17448 ( .A(n2263), .B(n5277), .Z(n2266) );
  MUX21L U17449 ( .A(n2264), .B(n2265), .S(n4628), .Z(n2267) );
  NR2 U17450 ( .A(n4963), .B(n4628), .Z(n2263) );
  NR2 U17451 ( .A(n5238), .B(n4580), .Z(n3086) );
  NR2 U17452 ( .A(n5259), .B(n4963), .Z(n2265) );
  EO U17453 ( .A(n5225), .B(n4917), .Z(n1430) );
  EN U17454 ( .A(n4899), .B(n4568), .Z(n1955) );
  EN U17455 ( .A(n5225), .B(n4584), .Z(n1950) );
  ND2 U17456 ( .A(n3594), .B(n4576), .Z(n2025) );
  EO U17457 ( .A(n5229), .B(n4926), .Z(n3594) );
  ND2 U17458 ( .A(n3458), .B(n3457), .Z(n2023) );
  EN U17459 ( .A(n5221), .B(n4591), .Z(n3458) );
  ND2 U17460 ( .A(n4919), .B(n4585), .Z(n3457) );
  ND2 U17461 ( .A(n3079), .B(n3078), .Z(n1475) );
  ND2 U17462 ( .A(n4941), .B(n4580), .Z(n3078) );
  MUX21L U17463 ( .A(n3077), .B(n4580), .S(n5235), .Z(n3079) );
  NR2 U17464 ( .A(n4941), .B(n4580), .Z(n3077) );
  ND2 U17465 ( .A(n2837), .B(n4564), .Z(n1471) );
  EO U17466 ( .A(n5230), .B(n4931), .Z(n2837) );
  ND2 U17467 ( .A(n2117), .B(n2116), .Z(n1455) );
  ND2 U17468 ( .A(n2113), .B(n5272), .Z(n2116) );
  MUX21L U17469 ( .A(n2114), .B(n2115), .S(n5272), .Z(n2117) );
  NR2 U17470 ( .A(n4912), .B(n4601), .Z(n2113) );
  ND2 U17471 ( .A(n2804), .B(n2803), .Z(n1437) );
  EN U17472 ( .A(n5222), .B(n4562), .Z(n2804) );
  EO U17473 ( .A(n4903), .B(n4562), .Z(n2803) );
  ND2 U17474 ( .A(n4914), .B(n4599), .Z(n2157) );
  ND2 U17475 ( .A(n2924), .B(n2923), .Z(n1947) );
  MUX21L U17476 ( .A(n2921), .B(n2922), .S(n5285), .Z(n2923) );
  MUX21L U17477 ( .A(n2919), .B(n2920), .S(n4969), .Z(n2924) );
  NR2 U17478 ( .A(n4968), .B(n4550), .Z(n2921) );
  ND2 U17479 ( .A(n3595), .B(n4926), .Z(n1957) );
  EO U17480 ( .A(n5228), .B(n4577), .Z(n3595) );
  MUX21L U17481 ( .A(n4636), .B(n5264), .S(n4977), .Z(n2002) );
  AO4 U17482 ( .A(n4973), .B(n4622), .C(n5290), .D(n4622), .Z(n1432) );
  NR2 U17483 ( .A(n4914), .B(n4615), .Z(n2432) );
  NR2 U17484 ( .A(n5276), .B(n4965), .Z(n1932) );
  EO U17485 ( .A(n5227), .B(n4908), .Z(n1928) );
  EO U17486 ( .A(n4899), .B(n4582), .Z(n3123) );
  ND3 U17487 ( .A(n3121), .B(n3120), .C(n3119), .Z(n1442) );
  ND2 U17488 ( .A(n4938), .B(n5239), .Z(n3121) );
  ND2 U17489 ( .A(n5239), .B(n4582), .Z(n3120) );
  ND2 U17490 ( .A(n4938), .B(n4582), .Z(n3119) );
  ND2 U17491 ( .A(n4914), .B(n4599), .Z(n2149) );
  ND2 U17492 ( .A(n4954), .B(n4588), .Z(n3212) );
  ND2 U17493 ( .A(n5244), .B(n3461), .Z(n1449) );
  ND2 U17494 ( .A(n4919), .B(n4568), .Z(n3461) );
  ND2 U17495 ( .A(n4620), .B(n2562), .Z(n1940) );
  ND2 U17496 ( .A(n5289), .B(n4974), .Z(n2562) );
  ND2 U17497 ( .A(n4944), .B(n4552), .Z(n3013) );
  ND2 U17498 ( .A(n3348), .B(n3347), .Z(n1414) );
  ND2 U17499 ( .A(n3344), .B(n5257), .Z(n3347) );
  MUX21L U17500 ( .A(n3345), .B(n3346), .S(n4606), .Z(n3348) );
  NR2 U17501 ( .A(n4935), .B(n4605), .Z(n3344) );
  AN2P U17502 ( .A(n4944), .B(n4553), .Z(n753) );
  MUX21L U17503 ( .A(n5260), .B(n4961), .S(n4631), .Z(n1460) );
  MUX21L U17504 ( .A(n4561), .B(n2784), .S(n4929), .Z(n1945) );
  ND2 U17505 ( .A(n5279), .B(n4561), .Z(n2784) );
  MUX21L U17506 ( .A(n4601), .B(n2112), .S(n5272), .Z(n1929) );
  ND2 U17507 ( .A(n4912), .B(n4601), .Z(n2112) );
  NR2 U17508 ( .A(n4917), .B(n4593), .Z(n2484) );
  NR2 U17509 ( .A(n5257), .B(n4935), .Z(n3346) );
  ND2 U17510 ( .A(n2044), .B(n2043), .Z(n1892) );
  MUX21L U17511 ( .A(n2041), .B(n2042), .S(n5269), .Z(n2043) );
  MUX21L U17512 ( .A(n2039), .B(n2040), .S(n4908), .Z(n2044) );
  NR2 U17513 ( .A(n4908), .B(n4627), .Z(n2041) );
  ND2 U17514 ( .A(n2204), .B(n4596), .Z(n1393) );
  EO U17515 ( .A(n5230), .B(n4966), .Z(n2204) );
  ND2 U17516 ( .A(n3170), .B(n3169), .Z(n1411) );
  ND2 U17517 ( .A(n4585), .B(n4956), .Z(n3169) );
  MUX21L U17518 ( .A(n3168), .B(n4956), .S(n5233), .Z(n3170) );
  NR2 U17519 ( .A(n4956), .B(n4585), .Z(n3168) );
  AO4 U17520 ( .A(n4930), .B(n4562), .C(n5280), .D(n4562), .Z(n1911) );
  NR2 U17521 ( .A(n5253), .B(n4612), .Z(n3259) );
  NR2 U17522 ( .A(n5258), .B(n4604), .Z(n3379) );
  NR2 U17523 ( .A(n5284), .B(n4566), .Z(n2888) );
  NR2 U17524 ( .A(n5237), .B(n4583), .Z(n3140) );
  EN U17525 ( .A(n5224), .B(n4637), .Z(n2399) );
  MUX21L U17526 ( .A(n2392), .B(n5264), .S(n4636), .Z(n1901) );
  ND2 U17527 ( .A(n5264), .B(n4977), .Z(n2392) );
  ND2 U17528 ( .A(n2411), .B(n2410), .Z(n1365) );
  ND2 U17529 ( .A(n2407), .B(n5265), .Z(n2410) );
  MUX21L U17530 ( .A(n2408), .B(n2409), .S(n5265), .Z(n2411) );
  NR2 U17531 ( .A(n4976), .B(n4632), .Z(n2407) );
  AO4 U17532 ( .A(n4917), .B(n4628), .C(n5269), .D(n4628), .Z(n1355) );
  AO7 U17533 ( .A(n5237), .B(n4554), .C(n4942), .Z(n1379) );
  NR2 U17534 ( .A(n5277), .B(n4906), .Z(n2724) );
  NR2 U17535 ( .A(n5272), .B(n4602), .Z(n2095) );
  EO U17536 ( .A(n4901), .B(n4560), .Z(n1874) );
  ND2 U17537 ( .A(n3549), .B(n5248), .Z(n1889) );
  EN U17538 ( .A(n4902), .B(n4574), .Z(n3549) );
  ND2 U17539 ( .A(n2169), .B(n4598), .Z(n1861) );
  EN U17540 ( .A(n5229), .B(n4968), .Z(n2169) );
  ND2 U17541 ( .A(n4905), .B(n4559), .Z(n1373) );
  NR2 U17542 ( .A(n4918), .B(n4589), .Z(n3412) );
  NR2 U17543 ( .A(n5242), .B(n4918), .Z(n3414) );
  ND2 U17544 ( .A(n3349), .B(n4605), .Z(n1351) );
  EN U17545 ( .A(n5223), .B(n4935), .Z(n3349) );
  ND2 U17546 ( .A(n2580), .B(n2579), .Z(n1334) );
  EN U17547 ( .A(n5226), .B(n4621), .Z(n2580) );
  EO U17548 ( .A(n4903), .B(n4621), .Z(n2579) );
  ND2 U17549 ( .A(n2601), .B(n2600), .Z(n1335) );
  EN U17550 ( .A(n4903), .B(n4622), .Z(n2601) );
  EN U17551 ( .A(n5226), .B(n4622), .Z(n2600) );
  MUX21L U17552 ( .A(n3091), .B(n4940), .S(n4581), .Z(n1345) );
  ND2 U17553 ( .A(n5239), .B(n4940), .Z(n3091) );
  MUX21L U17554 ( .A(n4934), .B(n4607), .S(n5256), .Z(n1886) );
  ND2 U17555 ( .A(n2225), .B(n2224), .Z(n1826) );
  ND2 U17556 ( .A(n4965), .B(n4595), .Z(n2224) );
  EO U17557 ( .A(n5230), .B(n4595), .Z(n2225) );
  EN U17558 ( .A(n5227), .B(n4577), .Z(n1855) );
  ND2 U17559 ( .A(n4964), .B(n4594), .Z(n1327) );
  NR2 U17560 ( .A(n4910), .B(n4597), .Z(n2081) );
  ND2 U17561 ( .A(n2436), .B(n4914), .Z(n1833) );
  EN U17562 ( .A(n5224), .B(n4616), .Z(n2436) );
  ND2 U17563 ( .A(n5277), .B(n4594), .Z(n2256) );
  MUX21L U17564 ( .A(n4592), .B(n2504), .S(n5287), .Z(n1834) );
  ND2 U17565 ( .A(n4913), .B(n4592), .Z(n2504) );
  ND2 U17566 ( .A(n5256), .B(n4607), .Z(n1852) );
  NR2 U17567 ( .A(n4932), .B(n4565), .Z(n2863) );
  ND2 U17568 ( .A(n4923), .B(n3528), .Z(n1322) );
  ND2 U17569 ( .A(n5247), .B(n4572), .Z(n3528) );
  ND2 U17570 ( .A(n2841), .B(n2840), .Z(n1311) );
  ND2 U17571 ( .A(n4931), .B(n5282), .Z(n2841) );
  ND2 U17572 ( .A(n5282), .B(n4564), .Z(n2840) );
  ND2 U17573 ( .A(n2965), .B(n2964), .Z(n1810) );
  ND2 U17574 ( .A(n4946), .B(n4549), .Z(n2964) );
  EN U17575 ( .A(n5227), .B(n4549), .Z(n2965) );
  ND2 U17576 ( .A(n3074), .B(n5233), .Z(n1812) );
  EO U17577 ( .A(n4898), .B(n4579), .Z(n3074) );
  ND2 U17578 ( .A(n3118), .B(n5239), .Z(n1813) );
  EO U17579 ( .A(n4899), .B(n4582), .Z(n3118) );
  ND2 U17580 ( .A(n2227), .B(n2226), .Z(n1794) );
  ND2 U17581 ( .A(n5276), .B(n4595), .Z(n2226) );
  EO U17582 ( .A(n4902), .B(n4595), .Z(n2227) );
  EO U17583 ( .A(n5228), .B(n4603), .Z(n1792) );
  ND2 U17584 ( .A(n3161), .B(n4956), .Z(n1815) );
  EO U17585 ( .A(n5225), .B(n4585), .Z(n3161) );
  ND2 U17586 ( .A(n4910), .B(n5271), .Z(n2071) );
  ND2 U17587 ( .A(n2506), .B(n2505), .Z(n1801) );
  ND2 U17588 ( .A(n5287), .B(n4592), .Z(n2505) );
  ND2 U17589 ( .A(n4904), .B(n5287), .Z(n2506) );
  MUX21L U17590 ( .A(n4572), .B(n3527), .S(n5246), .Z(n1820) );
  ND2 U17591 ( .A(n4922), .B(n4572), .Z(n3527) );
  ND2 U17592 ( .A(n5236), .B(n4942), .Z(n1315) );
  NR2 U17593 ( .A(n5271), .B(n4602), .Z(n2085) );
  NR2 U17594 ( .A(n4959), .B(n4634), .Z(n1798) );
  ND2 U17595 ( .A(n2914), .B(n2913), .Z(n1281) );
  ND2 U17596 ( .A(n4969), .B(n4562), .Z(n2913) );
  EO U17597 ( .A(n5228), .B(n4547), .Z(n2914) );
  EN U17598 ( .A(n5229), .B(n4599), .Z(n1268) );
  ND2 U17599 ( .A(n5264), .B(n4636), .Z(n1799) );
  ND2 U17600 ( .A(n5288), .B(n4608), .Z(n2519) );
  ND2 U17601 ( .A(n5261), .B(n4961), .Z(n2317) );
  MUX21L U17602 ( .A(n4554), .B(n4942), .S(n5234), .Z(n1283) );
  ND2 U17603 ( .A(n2077), .B(n2076), .Z(n1758) );
  ND2 U17604 ( .A(n2073), .B(n5271), .Z(n2076) );
  MUX21L U17605 ( .A(n2074), .B(n2075), .S(n5271), .Z(n2077) );
  NR2 U17606 ( .A(n4910), .B(n4626), .Z(n2073) );
  NR2 U17607 ( .A(n5238), .B(n4938), .Z(n3128) );
  ND2 U17608 ( .A(n3336), .B(n4934), .Z(n1785) );
  EN U17609 ( .A(n5224), .B(n4606), .Z(n3336) );
  ND2 U17610 ( .A(n3466), .B(n3465), .Z(n1786) );
  ND2 U17611 ( .A(n5244), .B(n4568), .Z(n3465) );
  EN U17612 ( .A(n5221), .B(n4920), .Z(n3466) );
  ND2 U17613 ( .A(n3006), .B(n4944), .Z(n1777) );
  EO U17614 ( .A(n5228), .B(n4552), .Z(n3006) );
  ND2 U17615 ( .A(n4926), .B(n3598), .Z(n1788) );
  ND2 U17616 ( .A(n5249), .B(n4577), .Z(n3598) );
  ND2 U17617 ( .A(n2959), .B(n2958), .Z(n1776) );
  ND2 U17618 ( .A(n4947), .B(n5286), .Z(n2959) );
  ND2 U17619 ( .A(n5286), .B(n4548), .Z(n2958) );
  ND2 U17620 ( .A(n2568), .B(n5289), .Z(n2571) );
  NR2 U17621 ( .A(n4974), .B(n4620), .Z(n2568) );
  AO4 U17622 ( .A(n5283), .B(n4565), .C(n5283), .D(n4932), .Z(n1775) );
  NR2 U17623 ( .A(n5274), .B(n4597), .Z(n2180) );
  ND2 U17624 ( .A(n4940), .B(n5239), .Z(n3093) );
  ND2 U17625 ( .A(n3609), .B(n3608), .Z(n1264) );
  ND2 U17626 ( .A(n4577), .B(n5250), .Z(n3608) );
  MUX21L U17627 ( .A(n3607), .B(n4927), .S(n5250), .Z(n3609) );
  NR2 U17628 ( .A(n4927), .B(n4577), .Z(n3607) );
  AO4 U17629 ( .A(n4958), .B(n4584), .C(n5236), .D(n4958), .Z(n1258) );
  EO U17630 ( .A(n5222), .B(n4580), .Z(n1747) );
  EO U17631 ( .A(n5223), .B(n4959), .Z(n1733) );
  ND2 U17632 ( .A(n2806), .B(n2805), .Z(n1742) );
  ND2 U17633 ( .A(n5280), .B(n4562), .Z(n2805) );
  EN U17634 ( .A(n5222), .B(n4929), .Z(n2806) );
  ND2 U17635 ( .A(n4611), .B(n3265), .Z(n1260) );
  ND2 U17636 ( .A(n5253), .B(n4951), .Z(n3265) );
  MUX21L U17637 ( .A(n4935), .B(n4605), .S(n5257), .Z(n1262) );
  NR2 U17638 ( .A(n5231), .B(n4587), .Z(n3194) );
  NR2 U17639 ( .A(n5281), .B(n4563), .Z(n2829) );
  ND3 U17640 ( .A(n3021), .B(n3020), .C(n3019), .Z(n1745) );
  ND2 U17641 ( .A(n5240), .B(n4553), .Z(n3020) );
  ND2 U17642 ( .A(n4944), .B(n5240), .Z(n3021) );
  ND2 U17643 ( .A(n4944), .B(n4553), .Z(n3019) );
  ND3 U17644 ( .A(n4938), .B(n4583), .C(n5238), .Z(n1749) );
  ND2 U17645 ( .A(n5265), .B(n2414), .Z(n1734) );
  ND2 U17646 ( .A(n4976), .B(n4614), .Z(n2414) );
  ND2 U17647 ( .A(n2229), .B(n2228), .Z(n1212) );
  ND2 U17648 ( .A(n5276), .B(n4595), .Z(n2228) );
  EO U17649 ( .A(n4902), .B(n4595), .Z(n2229) );
  ND2 U17650 ( .A(n3624), .B(n3623), .Z(n1236) );
  EN U17651 ( .A(n5227), .B(n4578), .Z(n3624) );
  EO U17652 ( .A(n4901), .B(n4578), .Z(n3623) );
  ND2 U17653 ( .A(n2514), .B(n2513), .Z(n1219) );
  ND2 U17654 ( .A(n2510), .B(n5288), .Z(n2513) );
  MUX21L U17655 ( .A(n2511), .B(n2512), .S(n5288), .Z(n2514) );
  NR2 U17656 ( .A(n4904), .B(n4591), .Z(n2510) );
  ND2 U17657 ( .A(n4618), .B(n4916), .Z(n2476) );
  ND2 U17658 ( .A(n5264), .B(n4978), .Z(n2379) );
  MUX21L U17659 ( .A(n2475), .B(n4916), .S(n5268), .Z(n2477) );
  NR2 U17660 ( .A(n4916), .B(n4618), .Z(n2475) );
  MUX21L U17661 ( .A(n4587), .B(n3205), .S(n4954), .Z(n1231) );
  ND2 U17662 ( .A(n5230), .B(n4587), .Z(n3205) );
  ND2 U17663 ( .A(n3541), .B(n3540), .Z(n1724) );
  ND2 U17664 ( .A(n5247), .B(n4573), .Z(n3540) );
  EO U17665 ( .A(n4902), .B(n4573), .Z(n3541) );
  EN U17666 ( .A(n4903), .B(n4611), .Z(n1720) );
  ND2 U17667 ( .A(n2974), .B(n2973), .Z(n1714) );
  ND2 U17668 ( .A(n5277), .B(n4550), .Z(n2973) );
  EO U17669 ( .A(n4898), .B(n4550), .Z(n2974) );
  ND2 U17670 ( .A(n2787), .B(n4929), .Z(n1711) );
  EO U17671 ( .A(n5223), .B(n4561), .Z(n2787) );
  EO U17672 ( .A(n4900), .B(n4618), .Z(n1706) );
  EO U17673 ( .A(n5224), .B(n4977), .Z(n1704) );
  ND2 U17674 ( .A(n5242), .B(n4937), .Z(n3407) );
  ND2 U17675 ( .A(n4600), .B(n4912), .Z(n2125) );
  MUX21L U17676 ( .A(n2124), .B(n4912), .S(n5272), .Z(n2126) );
  NR2 U17677 ( .A(n4912), .B(n4600), .Z(n2124) );
  ND2 U17678 ( .A(n2324), .B(n2323), .Z(n1701) );
  ND2 U17679 ( .A(n4632), .B(n5261), .Z(n2323) );
  MUX21L U17680 ( .A(n2322), .B(n4960), .S(n5261), .Z(n2324) );
  NR2 U17681 ( .A(n4960), .B(n4632), .Z(n2322) );
  EN U17682 ( .A(n5229), .B(n4552), .Z(n1198) );
  ND2 U17683 ( .A(n4962), .B(n4630), .Z(n2301) );
  ND2 U17684 ( .A(n5233), .B(n4956), .Z(n3171) );
  ND2 U17685 ( .A(n3611), .B(n3610), .Z(n1207) );
  EN U17686 ( .A(n4902), .B(n4577), .Z(n3611) );
  EO U17687 ( .A(n5227), .B(n4577), .Z(n3610) );
  MUX21L U17688 ( .A(n2457), .B(n4915), .S(n4617), .Z(n1189) );
  ND2 U17689 ( .A(n5267), .B(n4915), .Z(n2457) );
  ND2 U17690 ( .A(n2846), .B(n2845), .Z(n1196) );
  ND2 U17691 ( .A(n2842), .B(n5282), .Z(n2845) );
  MUX21L U17692 ( .A(n2843), .B(n2844), .S(n5282), .Z(n2846) );
  NR2 U17693 ( .A(n4931), .B(n4564), .Z(n2842) );
  NR2 U17694 ( .A(n5278), .B(n4560), .Z(n2762) );
  NR2 U17695 ( .A(n4964), .B(n4594), .Z(n1185) );
  ND2 U17696 ( .A(n2164), .B(n2163), .Z(n1669) );
  ND2 U17697 ( .A(n5274), .B(n4598), .Z(n2163) );
  EO U17698 ( .A(n4902), .B(n4598), .Z(n2164) );
  EO U17699 ( .A(n5221), .B(n4963), .Z(n1672) );
  ND2 U17700 ( .A(n5286), .B(n4549), .Z(n2960) );
  MUX21L U17701 ( .A(n2090), .B(n4911), .S(n4602), .Z(n1668) );
  ND2 U17702 ( .A(n5272), .B(n4911), .Z(n2090) );
  ND2 U17703 ( .A(n4940), .B(n4581), .Z(n1200) );
  ND2 U17704 ( .A(n3067), .B(n3066), .Z(n1171) );
  ND2 U17705 ( .A(n3063), .B(n5231), .Z(n3066) );
  MUX21L U17706 ( .A(n3064), .B(n3065), .S(n5231), .Z(n3067) );
  NR2 U17707 ( .A(n4941), .B(n4556), .Z(n3063) );
  ND2 U17708 ( .A(n3326), .B(n3325), .Z(n1176) );
  ND2 U17709 ( .A(n4948), .B(n5256), .Z(n3326) );
  ND2 U17710 ( .A(n5256), .B(n4607), .Z(n3325) );
  AN2P U17711 ( .A(n4974), .B(n4621), .Z(n754) );
  EO U17712 ( .A(n5226), .B(n4624), .Z(n1646) );
  ND2 U17713 ( .A(n2933), .B(n2932), .Z(n1653) );
  MUX21L U17714 ( .A(n2930), .B(n2931), .S(n5285), .Z(n2932) );
  MUX21L U17715 ( .A(n2928), .B(n2929), .S(n4943), .Z(n2933) );
  NR2 U17716 ( .A(n4948), .B(n4549), .Z(n2930) );
  ND2 U17717 ( .A(n3626), .B(n3625), .Z(n1665) );
  EO U17718 ( .A(n5227), .B(n4578), .Z(n3626) );
  EO U17719 ( .A(n4901), .B(n4578), .Z(n3625) );
  NR2 U17720 ( .A(n5251), .B(n4953), .Z(n1660) );
  NR2 U17721 ( .A(n4946), .B(n4551), .Z(n2975) );
  NR2 U17722 ( .A(n4976), .B(n4637), .Z(n1162) );
  EN U17723 ( .A(n5228), .B(n4942), .Z(n1655) );
  EO U17724 ( .A(n5226), .B(n4586), .Z(n1151) );
  ND2 U17725 ( .A(n5285), .B(n4969), .Z(n2916) );
  ND2 U17726 ( .A(n2420), .B(n2419), .Z(n1642) );
  ND2 U17727 ( .A(n5265), .B(n4615), .Z(n2419) );
  EO U17728 ( .A(n4899), .B(n4615), .Z(n2420) );
  ND2 U17729 ( .A(n5268), .B(n4917), .Z(n2480) );
  ND2 U17730 ( .A(n4962), .B(n4631), .Z(n2305) );
  ND2 U17731 ( .A(n5260), .B(n4631), .Z(n2306) );
  ND2 U17732 ( .A(n3025), .B(n3024), .Z(n1147) );
  ND2 U17733 ( .A(n5241), .B(n4553), .Z(n3024) );
  EO U17734 ( .A(n4900), .B(n4553), .Z(n3025) );
  ND2 U17735 ( .A(n3631), .B(n3630), .Z(n1156) );
  ND2 U17736 ( .A(n4927), .B(n4579), .Z(n3630) );
  EO U17737 ( .A(n5227), .B(n4579), .Z(n3631) );
  EN U17738 ( .A(n4902), .B(n4567), .Z(n1145) );
  MUX21L U17739 ( .A(n3488), .B(n5245), .S(n4570), .Z(n1664) );
  ND2 U17740 ( .A(n5245), .B(n4920), .Z(n3488) );
  MUX21L U17741 ( .A(n2358), .B(n4959), .S(n4634), .Z(n1641) );
  ND2 U17742 ( .A(n5263), .B(n4959), .Z(n2358) );
  NR2 U17743 ( .A(n5279), .B(n4560), .Z(n2766) );
  AO4 U17744 ( .A(n4958), .B(n4634), .C(n5263), .D(n4634), .Z(n1609) );
  NR3 U17745 ( .A(n4627), .B(n5270), .C(n4909), .Z(n1604) );
  EO U17746 ( .A(n4898), .B(n4551), .Z(n1622) );
  EN U17747 ( .A(n5229), .B(n4922), .Z(n1632) );
  EO U17748 ( .A(n4900), .B(n4619), .Z(n1613) );
  EO U17749 ( .A(n4897), .B(n4593), .Z(n1612) );
  ND2 U17750 ( .A(n3042), .B(n4943), .Z(n1623) );
  EN U17751 ( .A(n5230), .B(n4554), .Z(n3042) );
  ND2 U17752 ( .A(n2422), .B(n2421), .Z(n1610) );
  ND2 U17753 ( .A(n5266), .B(n4615), .Z(n2422) );
  ND2 U17754 ( .A(n4914), .B(n4615), .Z(n2421) );
  ND2 U17755 ( .A(n4944), .B(n4553), .Z(n3026) );
  ND2 U17756 ( .A(n5241), .B(n4553), .Z(n3027) );
  OR3 U17757 ( .A(n4629), .B(n5259), .C(n4963), .Z(n755) );
  NR2 U17758 ( .A(n757), .B(n758), .Z(n756) );
  EO U17759 ( .A(n4897), .B(n4555), .Z(n757) );
  EO U17760 ( .A(n5230), .B(n4555), .Z(n758) );
  MUX21L U17761 ( .A(n3084), .B(n5237), .S(n4580), .Z(n1624) );
  ND2 U17762 ( .A(n5237), .B(n4941), .Z(n3084) );
  EN U17763 ( .A(n5224), .B(n4607), .Z(n1131) );
  EN U17764 ( .A(n5225), .B(n4951), .Z(n1130) );
  AN2P U17765 ( .A(n4969), .B(n4567), .Z(n759) );
  NR2 U17766 ( .A(n5242), .B(n4918), .Z(n3409) );
  EN U17767 ( .A(n5230), .B(n4932), .Z(n2854) );
  EO U17768 ( .A(n5224), .B(n4935), .Z(n1599) );
  ND2 U17769 ( .A(n2939), .B(n2938), .Z(n1591) );
  MUX21L U17770 ( .A(n2936), .B(n2937), .S(n5285), .Z(n2938) );
  MUX21L U17771 ( .A(n2934), .B(n2935), .S(n4948), .Z(n2939) );
  NR2 U17772 ( .A(n4948), .B(n4547), .Z(n2936) );
  ND2 U17773 ( .A(n3107), .B(n4581), .Z(n1594) );
  EO U17774 ( .A(n5223), .B(n4939), .Z(n3107) );
  ND2 U17775 ( .A(n3544), .B(n3543), .Z(n1601) );
  MUX21L U17776 ( .A(n3542), .B(n4573), .S(n4923), .Z(n3543) );
  AO2 U17777 ( .A(n5247), .B(n4573), .C(n5247), .D(n4923), .Z(n3544) );
  NR2 U17778 ( .A(n5247), .B(n4573), .Z(n3542) );
  OR2 U17779 ( .A(n4972), .B(n4622), .Z(n760) );
  NR3 U17780 ( .A(n4584), .B(n5235), .C(n4957), .Z(n1111) );
  ND2 U17781 ( .A(n5282), .B(n4565), .Z(n2853) );
  ND2 U17782 ( .A(n4577), .B(n3599), .Z(n1602) );
  ND2 U17783 ( .A(n5249), .B(n4926), .Z(n3599) );
  ND2 U17784 ( .A(n5250), .B(n4953), .Z(n3219) );
  IVP U17785 ( .A(n1578), .Z(n4186) );
  AO7 U17786 ( .A(n5273), .B(n4913), .C(n4600), .Z(n1578) );
  ND2 U17787 ( .A(n5241), .B(n4553), .Z(n3029) );
  ND2 U17788 ( .A(n4943), .B(n4554), .Z(n3028) );
  ND2 U17789 ( .A(n3023), .B(n3022), .Z(n1566) );
  ND2 U17790 ( .A(n5241), .B(n4553), .Z(n3022) );
  EN U17791 ( .A(n5229), .B(n4944), .Z(n3023) );
  NR3 U17792 ( .A(n4559), .B(n5278), .C(n4905), .Z(n1561) );
  NR2 U17793 ( .A(n5242), .B(n4589), .Z(n3422) );
  NR2 U17794 ( .A(n762), .B(n763), .Z(n761) );
  EN U17795 ( .A(n4899), .B(n4568), .Z(n762) );
  AN2P U17796 ( .A(n5244), .B(n4568), .Z(n763) );
  ND2 U17797 ( .A(n3490), .B(n3489), .Z(n1555) );
  EN U17798 ( .A(n4900), .B(n4570), .Z(n3490) );
  EN U17799 ( .A(n5230), .B(n4570), .Z(n3489) );
  OR3 U17800 ( .A(n4594), .B(n5276), .C(n4965), .Z(n764) );
  ND2 U17801 ( .A(n4927), .B(n4579), .Z(n3632) );
  EO U17802 ( .A(n5227), .B(n4579), .Z(n3633) );
  ND2 U17803 ( .A(n3628), .B(n3627), .Z(n1539) );
  ND2 U17804 ( .A(n4927), .B(n4578), .Z(n3627) );
  EO U17805 ( .A(n5227), .B(n4578), .Z(n3628) );
  ND2 U17806 ( .A(n3492), .B(n3491), .Z(n1538) );
  EN U17807 ( .A(n4900), .B(n4570), .Z(n3492) );
  EN U17808 ( .A(n5230), .B(n4570), .Z(n3491) );
  NR2 U17809 ( .A(n5243), .B(n4590), .Z(n3442) );
  ND3 U17810 ( .A(n3397), .B(n3396), .C(n3395), .Z(n1536) );
  ND2 U17811 ( .A(n4937), .B(n5259), .Z(n3397) );
  ND2 U17812 ( .A(n5259), .B(n4603), .Z(n3396) );
  ND2 U17813 ( .A(n4937), .B(n4603), .Z(n3395) );
  NR2 U17814 ( .A(n5254), .B(n4610), .Z(n3294) );
  NR2 U17815 ( .A(n4921), .B(n4570), .Z(n3494) );
  ND2 U17816 ( .A(n3274), .B(n3273), .Z(n1521) );
  EO U17817 ( .A(n5225), .B(n4611), .Z(n3274) );
  EO U17818 ( .A(n4903), .B(n4611), .Z(n3273) );
  IVP U17819 ( .A(n1093), .Z(n4196) );
  AO4 U17820 ( .A(n4922), .B(n4571), .C(n5246), .D(n4571), .Z(n1093) );
  NR2 U17821 ( .A(n4943), .B(n4554), .Z(n1518) );
  ND2 U17822 ( .A(n3330), .B(n3329), .Z(n1513) );
  ND2 U17823 ( .A(n5256), .B(n4607), .Z(n3329) );
  EO U17824 ( .A(n4897), .B(n4607), .Z(n3330) );
  EO U17825 ( .A(n4898), .B(n4589), .Z(n1515) );
  AO4 U17826 ( .A(n4947), .B(n4549), .C(n5285), .D(n4547), .Z(n1510) );
  EN U17827 ( .A(n5228), .B(n4574), .Z(n3560) );
  NR2 U17828 ( .A(n4919), .B(n4590), .Z(n3446) );
  NR2 U17829 ( .A(n5243), .B(n4590), .Z(n3447) );
  ND2 U17830 ( .A(n4950), .B(n4611), .Z(n3277) );
  ND2 U17831 ( .A(n5253), .B(n4611), .Z(n3278) );
  MUX21H U17832 ( .A(n5248), .B(n4924), .S(n4574), .Z(n765) );
  ND2 U17833 ( .A(n5244), .B(n4590), .Z(n3450) );
  NR2 U17834 ( .A(n4927), .B(n4577), .Z(n3601) );
  ND3 U17835 ( .A(n4918), .B(n4589), .C(n5242), .Z(n1497) );
  NR2 U17836 ( .A(n5262), .B(n4633), .Z(n2333) );
  NR2 U17837 ( .A(n5249), .B(n4576), .Z(n3589) );
  AO4 U17838 ( .A(n4949), .B(n4608), .C(n5255), .D(n4608), .Z(n843) );
  ND2 U17839 ( .A(n4920), .B(n4569), .Z(n3473) );
  MUX21L U17840 ( .A(n2332), .B(n2333), .S(n4960), .Z(n2334) );
  MUX21L U17841 ( .A(n2330), .B(n2331), .S(n5262), .Z(n2335) );
  AO4 U17842 ( .A(n4974), .B(n4620), .C(n5289), .D(n4620), .Z(n828) );
  NR2 U17843 ( .A(n4966), .B(n4596), .Z(n2212) );
  NR2 U17844 ( .A(n5263), .B(n4635), .Z(n2367) );
  NR2 U17845 ( .A(n4927), .B(n4578), .Z(n3613) );
  NR2 U17846 ( .A(n5250), .B(n4578), .Z(n3614) );
  NR2 U17847 ( .A(n5258), .B(n4605), .Z(n3363) );
  NR2 U17848 ( .A(n4629), .B(n4962), .Z(n2283) );
  NR2 U17849 ( .A(n4915), .B(n4617), .Z(n2460) );
  ND2 U17850 ( .A(n2353), .B(n2352), .Z(n1002) );
  EN U17851 ( .A(n5222), .B(n4633), .Z(n2353) );
  EO U17852 ( .A(n4898), .B(n4633), .Z(n2352) );
  ND2 U17853 ( .A(n4966), .B(n5275), .Z(n2219) );
  ND2 U17854 ( .A(n3211), .B(n3210), .Z(n1020) );
  ND2 U17855 ( .A(n3207), .B(n4954), .Z(n3210) );
  MUX21L U17856 ( .A(n3208), .B(n3209), .S(n5231), .Z(n3211) );
  NR2 U17857 ( .A(n5230), .B(n4588), .Z(n3207) );
  ND2 U17858 ( .A(n2911), .B(n2910), .Z(n983) );
  ND2 U17859 ( .A(n4969), .B(n4567), .Z(n2910) );
  EN U17860 ( .A(n5228), .B(n4567), .Z(n2911) );
  ND2 U17861 ( .A(n3081), .B(n3080), .Z(n986) );
  ND2 U17862 ( .A(n5236), .B(n4580), .Z(n3080) );
  EO U17863 ( .A(n4898), .B(n4580), .Z(n3081) );
  ND2 U17864 ( .A(n2385), .B(n2384), .Z(n973) );
  EN U17865 ( .A(n5223), .B(n4636), .Z(n2385) );
  EO U17866 ( .A(n4897), .B(n4636), .Z(n2384) );
  ND2 U17867 ( .A(n2522), .B(n2521), .Z(n944) );
  EO U17868 ( .A(n5225), .B(n4614), .Z(n2522) );
  EO U17869 ( .A(n4899), .B(n4614), .Z(n2521) );
  ND2 U17870 ( .A(n2967), .B(n2966), .Z(n954) );
  ND2 U17871 ( .A(n4946), .B(n4550), .Z(n2966) );
  EN U17872 ( .A(n5227), .B(n4549), .Z(n2967) );
  ND2 U17873 ( .A(n2852), .B(n2851), .Z(n952) );
  ND2 U17874 ( .A(n4564), .B(n4932), .Z(n2851) );
  MUX21L U17875 ( .A(n2850), .B(n4932), .S(n5282), .Z(n2852) );
  NR2 U17876 ( .A(n4932), .B(n4564), .Z(n2850) );
  ND2 U17877 ( .A(n3468), .B(n3467), .Z(n873) );
  EO U17878 ( .A(n5230), .B(n4568), .Z(n3468) );
  EO U17879 ( .A(n4899), .B(n4568), .Z(n3467) );
  EN U17880 ( .A(n4902), .B(n4598), .Z(n1030) );
  EN U17881 ( .A(n5222), .B(n4962), .Z(n1033) );
  ND3 U17882 ( .A(n4898), .B(n4544), .C(n5222), .Z(n766) );
  IVP U17883 ( .A(n863), .Z(n4192) );
  AO4 U17884 ( .A(n4931), .B(n4563), .C(n5282), .D(n4563), .Z(n863) );
  ND2 U17885 ( .A(n2517), .B(n2516), .Z(n1037) );
  ND2 U17886 ( .A(n4591), .B(n5288), .Z(n2516) );
  MUX21L U17887 ( .A(n2515), .B(n4904), .S(n5288), .Z(n2517) );
  NR2 U17888 ( .A(n4904), .B(n4591), .Z(n2515) );
  ND2 U17889 ( .A(n2463), .B(n2462), .Z(n975) );
  MUX21L U17890 ( .A(n2458), .B(n2459), .S(n4915), .Z(n2463) );
  MUX21L U17891 ( .A(n2460), .B(n2461), .S(n5267), .Z(n2462) );
  NR3 U17892 ( .A(n4581), .B(n5241), .C(n4939), .Z(n866) );
  NR3 U17893 ( .A(n4559), .B(n5278), .C(n4905), .Z(n1010) );
  AO7 U17894 ( .A(n5287), .B(n4917), .C(n4592), .Z(n881) );
  AO4 U17895 ( .A(n4957), .B(n4584), .C(n5235), .D(n4957), .Z(n1079) );
  AO4 U17896 ( .A(n4957), .B(n4584), .C(n5234), .D(n4584), .Z(n988) );
  AO4 U17897 ( .A(n4916), .B(n4617), .C(n5267), .D(n4617), .Z(n909) );
  NR2 U17898 ( .A(n5249), .B(n4925), .Z(n1056) );
  NR2 U17899 ( .A(n5249), .B(n4926), .Z(n995) );
  NR2 U17900 ( .A(n4929), .B(n4561), .Z(n886) );
  NR2 U17901 ( .A(n4955), .B(n4586), .Z(n869) );
  AN3 U17902 ( .A(n4898), .B(n4545), .C(n5225), .Z(n1065) );
  EN U17903 ( .A(n5229), .B(n4566), .Z(n1043) );
  EO U17904 ( .A(n5230), .B(n4594), .Z(n1000) );
  EO U17905 ( .A(n5228), .B(n4912), .Z(n966) );
  EN U17906 ( .A(n5230), .B(n4966), .Z(n968) );
  EO U17907 ( .A(n5226), .B(n4620), .Z(n977) );
  EO U17908 ( .A(n4900), .B(n4599), .Z(n935) );
  EO U17909 ( .A(n5225), .B(n4908), .Z(n948) );
  EO U17910 ( .A(n5223), .B(n4905), .Z(n950) );
  EO U17911 ( .A(n5223), .B(n4939), .Z(n923) );
  EN U17912 ( .A(n5225), .B(n4611), .Z(n927) );
  EO U17913 ( .A(n5225), .B(n4957), .Z(n925) );
  EO U17914 ( .A(n4901), .B(n4586), .Z(n894) );
  EN U17915 ( .A(n5222), .B(n4936), .Z(n897) );
  EN U17916 ( .A(n5224), .B(n4948), .Z(n896) );
  ND2 U17917 ( .A(n4920), .B(n4569), .Z(n3475) );
  ND2 U17918 ( .A(n5244), .B(n4569), .Z(n3476) );
  ND2 U17919 ( .A(n4959), .B(n5262), .Z(n2346) );
  ND2 U17920 ( .A(n3470), .B(n3469), .Z(n855) );
  ND2 U17921 ( .A(n5244), .B(n4569), .Z(n3470) );
  ND2 U17922 ( .A(n4920), .B(n4569), .Z(n3469) );
  ND2 U17923 ( .A(n4940), .B(n4581), .Z(n1017) );
  ND2 U17924 ( .A(n3272), .B(n3271), .Z(n959) );
  ND2 U17925 ( .A(n5253), .B(n4951), .Z(n3272) );
  ND2 U17926 ( .A(n4950), .B(n4611), .Z(n3271) );
  ND2 U17927 ( .A(n2524), .B(n2523), .Z(n910) );
  ND2 U17928 ( .A(n4976), .B(n4614), .Z(n2523) );
  ND2 U17929 ( .A(n5288), .B(n4614), .Z(n2524) );
  ND2 U17930 ( .A(n3280), .B(n3279), .Z(n870) );
  ND2 U17931 ( .A(n5253), .B(n4611), .Z(n3280) );
  ND2 U17932 ( .A(n4950), .B(n4610), .Z(n3279) );
  AN2P U17933 ( .A(n4934), .B(n4607), .Z(n767) );
  MUX21L U17934 ( .A(n2370), .B(n4978), .S(n4635), .Z(n941) );
  ND2 U17935 ( .A(n5263), .B(n4978), .Z(n2370) );
  MUX21L U17936 ( .A(n2835), .B(n4931), .S(n4563), .Z(n918) );
  ND2 U17937 ( .A(n5281), .B(n4931), .Z(n2835) );
  MUX21L U17938 ( .A(n4576), .B(n5249), .S(n4926), .Z(n875) );
  ND2 U17939 ( .A(n4976), .B(n4637), .Z(n908) );
  MUX21L U17940 ( .A(n4919), .B(n5243), .S(n4589), .Z(n961) );
  IVP U17941 ( .A(n4368), .Z(n4548) );
  IVP U17942 ( .A(n4370), .Z(n4562) );
  IVP U17943 ( .A(n4724), .Z(n4956) );
  IVP U17944 ( .A(n4362), .Z(n4621) );
  IVP U17945 ( .A(n4362), .Z(n4618) );
  IVP U17946 ( .A(n4722), .Z(n4971) );
  IVP U17947 ( .A(n4364), .Z(n4610) );
  IVP U17948 ( .A(n4733), .Z(n4906) );
  IVP U17949 ( .A(n4368), .Z(n4551) );
  IVP U17950 ( .A(n5069), .Z(n5228) );
  IVP U17951 ( .A(n4370), .Z(n4560) );
  IVP U17952 ( .A(n4734), .Z(n4899) );
  IVP U17953 ( .A(n4373), .Z(n4578) );
  IVP U17954 ( .A(n5067), .Z(n5240) );
  IVP U17955 ( .A(n4733), .Z(n4903) );
  IVP U17956 ( .A(n4365), .Z(n4601) );
  IVP U17957 ( .A(n4361), .Z(n4626) );
  IVP U17958 ( .A(n5069), .Z(n5229) );
  IVP U17959 ( .A(n4361), .Z(n4627) );
  IVP U17960 ( .A(n5059), .Z(n5286) );
  IVP U17961 ( .A(n4734), .Z(n4900) );
  IVP U17962 ( .A(n4368), .Z(n4550) );
  IVP U17963 ( .A(n5067), .Z(n5241) );
  IVP U17964 ( .A(n4727), .Z(n4939) );
  IVP U17965 ( .A(n4727), .Z(n4897) );
  IVP U17966 ( .A(n4361), .Z(n4628) );
  IVP U17967 ( .A(n4724), .Z(n4961) );
  IVP U17968 ( .A(n4374), .Z(n4587) );
  IVP U17969 ( .A(n4369), .Z(n4559) );
  IVP U17970 ( .A(n4723), .Z(n4967) );
  IVP U17971 ( .A(n4370), .Z(n4565) );
  IVP U17972 ( .A(n5060), .Z(n5283) );
  IVP U17973 ( .A(n4727), .Z(n4943) );
  IVP U17974 ( .A(n5061), .Z(n5278) );
  IVP U17975 ( .A(n4729), .Z(n4932) );
  NR2 U17976 ( .A(n4967), .B(n5161), .Z(n2190) );
  NR2 U17977 ( .A(n4967), .B(n4464), .Z(n2191) );
  NR2 U17978 ( .A(n4587), .B(n5085), .Z(n3185) );
  NR2 U17979 ( .A(n4587), .B(n4834), .Z(n3186) );
  ND2 U17980 ( .A(n2123), .B(n2122), .Z(n1994) );
  ND2 U17981 ( .A(n5272), .B(n4457), .Z(n2122) );
  EO U17982 ( .A(n4901), .B(n4601), .Z(n2123) );
  ND2 U17983 ( .A(n2193), .B(n2192), .Z(n1996) );
  MUX21L U17984 ( .A(n2189), .B(n4597), .S(n5275), .Z(n2192) );
  NR2 U17985 ( .A(n2191), .B(n2190), .Z(n2193) );
  NR2 U17986 ( .A(n4596), .B(n4863), .Z(n2189) );
  ND2 U17987 ( .A(n2918), .B(n2917), .Z(n2014) );
  ND2 U17988 ( .A(n4397), .B(n5185), .Z(n2917) );
  EN U17989 ( .A(n4901), .B(n4550), .Z(n2918) );
  ND2 U17990 ( .A(n2754), .B(n2753), .Z(n2010) );
  ND2 U17991 ( .A(n4904), .B(n4500), .Z(n2753) );
  EO U17992 ( .A(n5223), .B(n4559), .Z(n2754) );
  ND2 U17993 ( .A(n2472), .B(n2471), .Z(n2003) );
  ND2 U17994 ( .A(n4618), .B(n5135), .Z(n2471) );
  EO U17995 ( .A(n4898), .B(n4618), .Z(n2472) );
  ND2 U17996 ( .A(n2682), .B(n5205), .Z(n2007) );
  EO U17997 ( .A(n4897), .B(n4626), .Z(n2682) );
  ND2 U17998 ( .A(n3188), .B(n3187), .Z(n2019) );
  MUX21L U17999 ( .A(n3184), .B(n4954), .S(n5231), .Z(n3187) );
  NR2 U18000 ( .A(n3186), .B(n3185), .Z(n3188) );
  NR2 U18001 ( .A(n4954), .B(n4435), .Z(n3184) );
  ND2 U18002 ( .A(n3165), .B(n3164), .Z(n2018) );
  ND2 U18003 ( .A(n4585), .B(n5090), .Z(n3164) );
  EO U18004 ( .A(n5226), .B(n4956), .Z(n3165) );
  ND2 U18005 ( .A(n4551), .B(n5179), .Z(n2984) );
  ND2 U18006 ( .A(n2111), .B(n2110), .Z(n1961) );
  ND2 U18007 ( .A(n4852), .B(n5168), .Z(n2110) );
  MUX21L U18008 ( .A(n4852), .B(n2109), .S(n4601), .Z(n2111) );
  ND2 U18009 ( .A(n2038), .B(n2037), .Z(n1960) );
  ND2 U18010 ( .A(n4627), .B(n5174), .Z(n2037) );
  EN U18011 ( .A(n4901), .B(n4627), .Z(n2038) );
  ND2 U18012 ( .A(n2308), .B(n2307), .Z(n1966) );
  ND2 U18013 ( .A(n5260), .B(n4539), .Z(n2307) );
  EN U18014 ( .A(n5222), .B(n4961), .Z(n2308) );
  ND2 U18015 ( .A(n2592), .B(n2591), .Z(n1973) );
  ND2 U18016 ( .A(n4973), .B(n4520), .Z(n2591) );
  EN U18017 ( .A(n5226), .B(n4621), .Z(n2592) );
  ND2 U18018 ( .A(n2688), .B(n2687), .Z(n1975) );
  ND2 U18019 ( .A(n4508), .B(n4756), .Z(n2687) );
  EN U18020 ( .A(n5225), .B(n4906), .Z(n2688) );
  ND2 U18021 ( .A(n2388), .B(n2387), .Z(n1969) );
  ND2 U18022 ( .A(n4530), .B(n5142), .Z(n2387) );
  EN U18023 ( .A(n4897), .B(n4636), .Z(n2388) );
  ND2 U18024 ( .A(n3618), .B(n3617), .Z(n1990) );
  ND2 U18025 ( .A(n5250), .B(n4411), .Z(n3617) );
  EO U18026 ( .A(n4902), .B(n4578), .Z(n3618) );
  ND2 U18027 ( .A(n3190), .B(n3189), .Z(n1984) );
  ND2 U18028 ( .A(n4587), .B(n4834), .Z(n3189) );
  EO U18029 ( .A(n5226), .B(n4587), .Z(n3190) );
  MUX21L U18030 ( .A(n2856), .B(n5190), .S(n4565), .Z(n2858) );
  ND2 U18031 ( .A(n2640), .B(n2639), .Z(n1465) );
  ND2 U18032 ( .A(n4971), .B(n4624), .Z(n2639) );
  MUX21L U18033 ( .A(n2638), .B(n5209), .S(n4624), .Z(n2640) );
  NR2 U18034 ( .A(n4971), .B(n5209), .Z(n2638) );
  IVP U18035 ( .A(n5067), .Z(n5238) );
  IVP U18036 ( .A(n4365), .Z(n4603) );
  IVP U18037 ( .A(n4374), .Z(n4585) );
  IVP U18038 ( .A(n4372), .Z(n4573) );
  IVP U18039 ( .A(n4366), .Z(n4595) );
  IVP U18040 ( .A(n4732), .Z(n4910) );
  IVP U18041 ( .A(n5061), .Z(n5273) );
  IVP U18042 ( .A(n4723), .Z(n4965) );
  IVP U18043 ( .A(n4728), .Z(n4933) );
  IVP U18044 ( .A(n4369), .Z(n4557) );
  IVP U18045 ( .A(n4721), .Z(n4977) );
  IVP U18046 ( .A(n4366), .Z(n4596) );
  IVP U18047 ( .A(n4364), .Z(n4608) );
  IVP U18048 ( .A(n5066), .Z(n5245) );
  IVP U18049 ( .A(n5067), .Z(n5239) );
  IVP U18050 ( .A(n4729), .Z(n4927) );
  IVP U18051 ( .A(n4373), .Z(n4577) );
  IVP U18052 ( .A(n4723), .Z(n4963) );
  IVP U18053 ( .A(n4724), .Z(n4958) );
  IVP U18054 ( .A(n4365), .Z(n4602) );
  IVP U18055 ( .A(n4727), .Z(n4941) );
  IVP U18056 ( .A(n4369), .Z(n4554) );
  IVP U18057 ( .A(n4729), .Z(n4930) );
  IVP U18058 ( .A(n4374), .Z(n4584) );
  IVP U18059 ( .A(n4725), .Z(n4952) );
  IVP U18060 ( .A(n5069), .Z(n5227) );
  IVP U18061 ( .A(n5066), .Z(n5244) );
  IVP U18062 ( .A(n4375), .Z(n4591) );
  IVP U18063 ( .A(n4721), .Z(n4974) );
  IVP U18064 ( .A(n4371), .Z(n4569) );
  IVP U18065 ( .A(n5069), .Z(n5226) );
  IVP U18066 ( .A(n4367), .Z(n4546) );
  IVP U18067 ( .A(n5059), .Z(n5288) );
  IVP U18068 ( .A(n4733), .Z(n4904) );
  IVP U18069 ( .A(n5070), .Z(n5222) );
  IVP U18070 ( .A(n4361), .Z(n4625) );
  IVP U18071 ( .A(n4367), .Z(n4545) );
  IVP U18072 ( .A(n5070), .Z(n5225) );
  IVP U18073 ( .A(n4367), .Z(n4547) );
  IVP U18074 ( .A(n4721), .Z(n4976) );
  IVP U18075 ( .A(n4732), .Z(n4912) );
  IVP U18076 ( .A(n4733), .Z(n4905) );
  IVP U18077 ( .A(n4722), .Z(n4970) );
  IVP U18078 ( .A(n5065), .Z(n5252) );
  IVP U18079 ( .A(n4726), .Z(n4945) );
  IVP U18080 ( .A(n4727), .Z(n4940) );
  IVP U18081 ( .A(n5065), .Z(n5250) );
  IVP U18082 ( .A(n4728), .Z(n4936) );
  IVP U18083 ( .A(n4371), .Z(n4568) );
  IVP U18084 ( .A(n4734), .Z(n4898) );
  IVP U18085 ( .A(n4369), .Z(n4556) );
  IVP U18086 ( .A(n4373), .Z(n4580) );
  IVP U18087 ( .A(n4729), .Z(n4929) );
  IVP U18088 ( .A(n5062), .Z(n5267) );
  IVP U18089 ( .A(n4731), .Z(n4917) );
  IVP U18090 ( .A(n5059), .Z(n5287) );
  IVP U18091 ( .A(n4361), .Z(n4624) );
  IVP U18092 ( .A(n4725), .Z(n4951) );
  IVP U18093 ( .A(n5061), .Z(n5275) );
  IVP U18094 ( .A(n4366), .Z(n4597) );
  IVP U18095 ( .A(n4731), .Z(n4916) );
  IVP U18096 ( .A(n4730), .Z(n4923) );
  IVP U18097 ( .A(n4371), .Z(n4566) );
  IVP U18098 ( .A(n4734), .Z(n4901) );
  IVP U18099 ( .A(n4365), .Z(n4604) );
  IVP U18100 ( .A(n5064), .Z(n5258) );
  IVP U18101 ( .A(n4364), .Z(n4609) );
  IVP U18102 ( .A(n4362), .Z(n4620) );
  IVP U18103 ( .A(n4723), .Z(n4964) );
  IVP U18104 ( .A(n4373), .Z(n4579) );
  IVP U18105 ( .A(n5064), .Z(n5259) );
  IVP U18106 ( .A(n5064), .Z(n5221) );
  IVP U18107 ( .A(n4369), .Z(n4558) );
  IVP U18108 ( .A(n4366), .Z(n4600) );
  IVP U18109 ( .A(n4732), .Z(n4913) );
  IVP U18110 ( .A(n4728), .Z(n4937) );
  IVP U18111 ( .A(n4373), .Z(n4581) );
  IVP U18112 ( .A(n4732), .Z(n4914) );
  IVP U18113 ( .A(n5063), .Z(n5266) );
  IVP U18114 ( .A(n4373), .Z(n4582) );
  IVP U18115 ( .A(n4726), .Z(n4948) );
  IVP U18116 ( .A(n4731), .Z(n4920) );
  IVP U18117 ( .A(n4724), .Z(n4960) );
  IVP U18118 ( .A(n4360), .Z(n4635) );
  IVP U18119 ( .A(n4372), .Z(n4576) );
  IVP U18120 ( .A(n4360), .Z(n4634) );
  IVP U18121 ( .A(n4722), .Z(n4973) );
  IVP U18122 ( .A(n5059), .Z(n5290) );
  IVP U18123 ( .A(n5069), .Z(n5230) );
  IVP U18124 ( .A(n5064), .Z(n5260) );
  IVP U18125 ( .A(n4371), .Z(n4592) );
  IVP U18126 ( .A(n4734), .Z(n4902) );
  IVP U18127 ( .A(n4368), .Z(n4552) );
  IVP U18128 ( .A(n4366), .Z(n4599) );
  IVP U18129 ( .A(n5069), .Z(n5231) );
  IVP U18130 ( .A(n4725), .Z(n4954) );
  IVP U18131 ( .A(n4731), .Z(n4919) );
  IVP U18132 ( .A(n5062), .Z(n5272) );
  IVP U18133 ( .A(n5059), .Z(n5289) );
  IVP U18134 ( .A(n4364), .Z(n4612) );
  IVP U18135 ( .A(n5065), .Z(n5255) );
  IVP U18136 ( .A(n5061), .Z(n5277) );
  IVP U18137 ( .A(n4729), .Z(n4931) );
  IVP U18138 ( .A(n4730), .Z(n4926) );
  AO7 U18139 ( .A(n5275), .B(n4467), .C(n2223), .Z(n1422) );
  ND2 U18140 ( .A(n4965), .B(n4595), .Z(n2223) );
  AO7 U18141 ( .A(n5271), .B(n4452), .C(n2078), .Z(n1419) );
  ND2 U18142 ( .A(n4910), .B(n4626), .Z(n2078) );
  AO7 U18143 ( .A(n4908), .B(n4506), .C(n2710), .Z(n1434) );
  ND2 U18144 ( .A(n5295), .B(n4557), .Z(n2710) );
  AO7 U18145 ( .A(n4617), .B(n5137), .C(n2466), .Z(n1970) );
  ND2 U18146 ( .A(n5267), .B(n4916), .Z(n2466) );
  AO7 U18147 ( .A(n5233), .B(n4831), .C(n3166), .Z(n1983) );
  ND2 U18148 ( .A(n4956), .B(n4585), .Z(n3166) );
  AO7 U18149 ( .A(n4608), .B(n5072), .C(n3312), .Z(n1986) );
  ND2 U18150 ( .A(n5255), .B(n4948), .Z(n3312) );
  NR2 U18151 ( .A(n4620), .B(n4886), .Z(n2557) );
  NR2 U18152 ( .A(n4974), .B(n5216), .Z(n2558) );
  NR2 U18153 ( .A(n4912), .B(n4457), .Z(n2114) );
  NR2 U18154 ( .A(n5273), .B(n4767), .Z(n2142) );
  NR2 U18155 ( .A(n5273), .B(n4870), .Z(n2264) );
  ND2 U18156 ( .A(n5266), .B(n4914), .Z(n2429) );
  ND3 U18157 ( .A(n3117), .B(n3116), .C(n3115), .Z(n2016) );
  ND2 U18158 ( .A(n4582), .B(n5093), .Z(n3116) );
  ND2 U18159 ( .A(n4939), .B(n5093), .Z(n3117) );
  ND2 U18160 ( .A(n4939), .B(n4582), .Z(n3115) );
  ND3 U18161 ( .A(n2983), .B(n2982), .C(n2981), .Z(n2015) );
  ND2 U18162 ( .A(n4391), .B(n5180), .Z(n2982) );
  ND2 U18163 ( .A(n4945), .B(n5180), .Z(n2983) );
  ND2 U18164 ( .A(n4945), .B(n4391), .Z(n2981) );
  ND2 U18165 ( .A(n2561), .B(n2560), .Z(n2005) );
  NR2 U18166 ( .A(n2559), .B(n2558), .Z(n2561) );
  MUX21L U18167 ( .A(n2557), .B(n4620), .S(n5289), .Z(n2560) );
  NR2 U18168 ( .A(n4974), .B(n4524), .Z(n2559) );
  ND2 U18169 ( .A(n3387), .B(n3386), .Z(n2022) );
  ND2 U18170 ( .A(n4603), .B(n4937), .Z(n3386) );
  MUX21L U18171 ( .A(n3385), .B(n5108), .S(n4937), .Z(n3387) );
  NR2 U18172 ( .A(n4603), .B(n5108), .Z(n3385) );
  ND2 U18173 ( .A(n3479), .B(n3478), .Z(n2024) );
  ND2 U18174 ( .A(n4569), .B(n4781), .Z(n3478) );
  MUX21L U18175 ( .A(n5244), .B(n3477), .S(n4920), .Z(n3479) );
  NR2 U18176 ( .A(n5245), .B(n4569), .Z(n3477) );
  ND2 U18177 ( .A(n3088), .B(n3087), .Z(n1476) );
  MUX21L U18178 ( .A(n3085), .B(n5094), .S(n4940), .Z(n3087) );
  AO6 U18179 ( .A(n4940), .B(n4380), .C(n3086), .Z(n3088) );
  ND2 U18180 ( .A(n2757), .B(n4499), .Z(n1469) );
  EN U18181 ( .A(n5223), .B(n4903), .Z(n2757) );
  ND2 U18182 ( .A(n2802), .B(n2801), .Z(n1470) );
  ND2 U18183 ( .A(n4562), .B(n5194), .Z(n2801) );
  EO U18184 ( .A(n5222), .B(n4929), .Z(n2802) );
  ND2 U18185 ( .A(n3012), .B(n3011), .Z(n1474) );
  ND2 U18186 ( .A(n4552), .B(n4813), .Z(n3011) );
  MUX21L U18187 ( .A(n3010), .B(n5238), .S(n4552), .Z(n3012) );
  NR2 U18188 ( .A(n5239), .B(n4813), .Z(n3010) );
  ND2 U18189 ( .A(n2895), .B(n2894), .Z(n1472) );
  ND2 U18190 ( .A(n4799), .B(n5187), .Z(n2894) );
  MUX21L U18191 ( .A(n4800), .B(n2893), .S(n4566), .Z(n2895) );
  ND2 U18192 ( .A(n3299), .B(n3298), .Z(n1481) );
  ND2 U18193 ( .A(n4609), .B(n5074), .Z(n3298) );
  MUX21L U18194 ( .A(n4846), .B(n3297), .S(n5254), .Z(n3299) );
  NR2 U18195 ( .A(n4609), .B(n4846), .Z(n3297) );
  ND2 U18196 ( .A(n3384), .B(n3383), .Z(n1482) );
  ND2 U18197 ( .A(n4604), .B(n4789), .Z(n3383) );
  EO U18198 ( .A(n5223), .B(n4603), .Z(n3384) );
  ND2 U18199 ( .A(n3163), .B(n3162), .Z(n1478) );
  ND2 U18200 ( .A(n4585), .B(n4831), .Z(n3162) );
  EO U18201 ( .A(n5226), .B(n4585), .Z(n3163) );
  ND2 U18202 ( .A(n3606), .B(n3605), .Z(n1485) );
  ND2 U18203 ( .A(n4411), .B(n4768), .Z(n3605) );
  EO U18204 ( .A(n5227), .B(n4927), .Z(n3606) );
  ND2 U18205 ( .A(n2034), .B(n2033), .Z(n1453) );
  ND2 U18206 ( .A(n4444), .B(n4860), .Z(n2033) );
  EN U18207 ( .A(n5227), .B(n4628), .Z(n2034) );
  ND2 U18208 ( .A(n2144), .B(n2143), .Z(n1456) );
  ND2 U18209 ( .A(n2140), .B(n5166), .Z(n2143) );
  MUX21L U18210 ( .A(n2141), .B(n2142), .S(n4600), .Z(n2144) );
  NR2 U18211 ( .A(n4600), .B(n4913), .Z(n2140) );
  ND2 U18212 ( .A(n2092), .B(n2091), .Z(n1420) );
  ND2 U18213 ( .A(n4911), .B(n4455), .Z(n2091) );
  EN U18214 ( .A(n5228), .B(n4602), .Z(n2092) );
  ND2 U18215 ( .A(n2874), .B(n2873), .Z(n1439) );
  ND2 U18216 ( .A(n4933), .B(n4400), .Z(n2873) );
  MUX21L U18217 ( .A(n2872), .B(n4400), .S(n5284), .Z(n2874) );
  NR2 U18218 ( .A(n4933), .B(n4399), .Z(n2872) );
  ND2 U18219 ( .A(n3392), .B(n3391), .Z(n1448) );
  ND2 U18220 ( .A(n4603), .B(n5109), .Z(n3391) );
  EO U18221 ( .A(n4898), .B(n4603), .Z(n3392) );
  ND2 U18222 ( .A(n3629), .B(n5133), .Z(n1451) );
  EO U18223 ( .A(n4901), .B(n4579), .Z(n3629) );
  ND2 U18224 ( .A(n3319), .B(n3318), .Z(n1447) );
  ND2 U18225 ( .A(n4608), .B(n4825), .Z(n3318) );
  MUX21L U18226 ( .A(n3317), .B(n5255), .S(n4608), .Z(n3319) );
  NR2 U18227 ( .A(n5255), .B(n4849), .Z(n3317) );
  ND2 U18228 ( .A(n2371), .B(n5144), .Z(n1427) );
  EN U18229 ( .A(n4897), .B(n4635), .Z(n2371) );
  ND2 U18230 ( .A(n2648), .B(n2647), .Z(n1433) );
  ND3 U18231 ( .A(n4971), .B(n4515), .C(n5292), .Z(n2647) );
  MUX21L U18232 ( .A(n2645), .B(n2646), .S(n4971), .Z(n2648) );
  NR2 U18233 ( .A(n5292), .B(n4515), .Z(n2646) );
  ND2 U18234 ( .A(n3400), .B(n3399), .Z(n1988) );
  ND2 U18235 ( .A(n4937), .B(n4432), .Z(n3399) );
  MUX21L U18236 ( .A(n3398), .B(n4432), .S(n5255), .Z(n3400) );
  NR2 U18237 ( .A(n4937), .B(n4432), .Z(n3398) );
  ND2 U18238 ( .A(n3539), .B(n5125), .Z(n1989) );
  ND2 U18239 ( .A(n4923), .B(n4573), .Z(n3539) );
  ND2 U18240 ( .A(n2809), .B(n2808), .Z(n1946) );
  ND2 U18241 ( .A(n4408), .B(n4741), .Z(n2808) );
  EN U18242 ( .A(n5222), .B(n4562), .Z(n2809) );
  ND2 U18243 ( .A(n2714), .B(n5203), .Z(n1943) );
  EO U18244 ( .A(n4901), .B(n4558), .Z(n2714) );
  ND2 U18245 ( .A(n2435), .B(n2434), .Z(n1938) );
  MUX21L U18246 ( .A(n2432), .B(n2433), .S(n5266), .Z(n2434) );
  MUX21L U18247 ( .A(n2430), .B(n2431), .S(n4914), .Z(n2435) );
  NR2 U18248 ( .A(n4616), .B(n4765), .Z(n2433) );
  AN3 U18249 ( .A(n4815), .B(n5101), .C(n4554), .Z(n768) );
  MUX21L U18250 ( .A(n2262), .B(n2261), .S(n4964), .Z(n1998) );
  ND2 U18251 ( .A(n5277), .B(n4542), .Z(n2262) );
  ND2 U18252 ( .A(n4628), .B(n5153), .Z(n2261) );
  MUX21L U18253 ( .A(n4861), .B(n5269), .S(n4628), .Z(n1992) );
  MUX21L U18254 ( .A(n2156), .B(n4460), .S(n4914), .Z(n1995) );
  ND2 U18255 ( .A(n4460), .B(n5164), .Z(n2156) );
  MUX21L U18256 ( .A(n5294), .B(n4906), .S(n4556), .Z(n2008) );
  MUX21L U18257 ( .A(n5264), .B(n4881), .S(n4635), .Z(n2001) );
  MUX21L U18258 ( .A(n4889), .B(n4621), .S(n5290), .Z(n2006) );
  MUX21L U18259 ( .A(n3253), .B(n3252), .S(n5252), .Z(n2020) );
  ND2 U18260 ( .A(n4952), .B(n4481), .Z(n3253) );
  ND2 U18261 ( .A(n4952), .B(n4612), .Z(n3252) );
  MUX21L U18262 ( .A(n4907), .B(n5294), .S(n4557), .Z(n1467) );
  MUX21L U18263 ( .A(n2526), .B(n2525), .S(n4976), .Z(n1972) );
  ND2 U18264 ( .A(n5288), .B(n4618), .Z(n2526) );
  ND2 U18265 ( .A(n4618), .B(n5219), .Z(n2525) );
  MUX21L U18266 ( .A(n2503), .B(n2502), .S(n4917), .Z(n1971) );
  ND2 U18267 ( .A(n5287), .B(n4476), .Z(n2503) );
  ND2 U18268 ( .A(n5287), .B(n4592), .Z(n2502) );
  MUX21L U18269 ( .A(n5204), .B(n4509), .S(n4905), .Z(n1974) );
  MUX21L U18270 ( .A(n3375), .B(n3374), .S(n5258), .Z(n1987) );
  ND2 U18271 ( .A(n4493), .B(n4790), .Z(n3375) );
  ND2 U18272 ( .A(n4936), .B(n4604), .Z(n3374) );
  MUX21L U18273 ( .A(n3255), .B(n3254), .S(n5252), .Z(n1985) );
  ND2 U18274 ( .A(n4612), .B(n4842), .Z(n3255) );
  ND2 U18275 ( .A(n4951), .B(n4612), .Z(n3254) );
  IVP U18276 ( .A(n4364), .Z(n4607) );
  IVP U18277 ( .A(n5063), .Z(n5264) );
  IVP U18278 ( .A(n5060), .Z(n5280) );
  IVP U18279 ( .A(n4374), .Z(n4583) );
  IVP U18280 ( .A(n5064), .Z(n5256) );
  IVP U18281 ( .A(n4363), .Z(n4616) );
  IVP U18282 ( .A(n4722), .Z(n4968) );
  IVP U18283 ( .A(n4362), .Z(n4619) );
  IVP U18284 ( .A(n4732), .Z(n4911) );
  IVP U18285 ( .A(n4722), .Z(n4969) );
  IVP U18286 ( .A(n4363), .Z(n4615) );
  IVP U18287 ( .A(n5063), .Z(n5261) );
  IVP U18288 ( .A(n5068), .Z(n5233) );
  IVP U18289 ( .A(n4360), .Z(n4631) );
  IVP U18290 ( .A(n4372), .Z(n4571) );
  IVP U18291 ( .A(n4367), .Z(n4593) );
  IVP U18292 ( .A(n5065), .Z(n5251) );
  IVP U18293 ( .A(n5060), .Z(n5281) );
  IVP U18294 ( .A(n4730), .Z(n4924) );
  IVP U18295 ( .A(n4363), .Z(n4613) );
  IVP U18296 ( .A(n5063), .Z(n5263) );
  IVP U18297 ( .A(n5070), .Z(n5223) );
  IVP U18298 ( .A(n4723), .Z(n4962) );
  IVP U18299 ( .A(n5070), .Z(n5224) );
  IVP U18300 ( .A(n4728), .Z(n4934) );
  IVP U18301 ( .A(n4721), .Z(n4975) );
  IVP U18302 ( .A(n5060), .Z(n5279) );
  IVP U18303 ( .A(n4360), .Z(n4630) );
  IVP U18304 ( .A(n5061), .Z(n5274) );
  IVP U18305 ( .A(n4726), .Z(n4944) );
  IVP U18306 ( .A(n4726), .Z(n4947) );
  IVP U18307 ( .A(n5063), .Z(n5262) );
  IVP U18308 ( .A(n4731), .Z(n4915) );
  IVP U18309 ( .A(n4359), .Z(n4636) );
  IVP U18310 ( .A(n5059), .Z(n5285) );
  IVP U18311 ( .A(n4368), .Z(n4549) );
  IVP U18312 ( .A(n4370), .Z(n4561) );
  IVP U18313 ( .A(n5068), .Z(n5235) );
  IVP U18314 ( .A(n5062), .Z(n5268) );
  IVP U18315 ( .A(n5062), .Z(n5269) );
  IVP U18316 ( .A(n4728), .Z(n4938) );
  IVP U18317 ( .A(n5062), .Z(n5271) );
  IVP U18318 ( .A(n4733), .Z(n4907) );
  IVP U18319 ( .A(n5063), .Z(n5265) );
  IVP U18320 ( .A(n5060), .Z(n5284) );
  IVP U18321 ( .A(n4362), .Z(n4622) );
  IVP U18322 ( .A(n4368), .Z(n4553) );
  IVP U18323 ( .A(n5065), .Z(n5254) );
  IVP U18324 ( .A(n4363), .Z(n4617) );
  IVP U18325 ( .A(n4365), .Z(n4606) );
  IVP U18326 ( .A(n4372), .Z(n4575) );
  IVP U18327 ( .A(n4721), .Z(n4978) );
  IVP U18328 ( .A(n4362), .Z(n4623) );
  IVP U18329 ( .A(n4370), .Z(n4564) );
  IVP U18330 ( .A(n5068), .Z(n5237) );
  IVP U18331 ( .A(n4361), .Z(n4629) );
  IVP U18332 ( .A(n4374), .Z(n4588) );
  IVP U18333 ( .A(n4733), .Z(n4908) );
  AO7 U18334 ( .A(n5268), .B(n4761), .C(n4593), .Z(n2004) );
  AO7 U18335 ( .A(n5259), .B(n4870), .C(n4629), .Z(n1459) );
  AO7 U18336 ( .A(n4916), .B(n4526), .C(n2467), .Z(n1429) );
  ND2 U18337 ( .A(n5267), .B(n4617), .Z(n2467) );
  AO7 U18338 ( .A(n5264), .B(n4978), .C(n4531), .Z(n1968) );
  AO7 U18339 ( .A(n4970), .B(n4511), .C(n2667), .Z(n1942) );
  ND2 U18340 ( .A(n5293), .B(n4625), .Z(n2667) );
  AO7 U18341 ( .A(n4596), .B(n4864), .C(n2194), .Z(n1931) );
  ND2 U18342 ( .A(n5275), .B(n4967), .Z(n2194) );
  NR2 U18343 ( .A(n5285), .B(n4396), .Z(n2920) );
  NR2 U18344 ( .A(n4549), .B(n4803), .Z(n2922) );
  NR2 U18345 ( .A(n5266), .B(n4528), .Z(n2431) );
  NR2 U18346 ( .A(n4628), .B(n4860), .Z(n1927) );
  NR2 U18347 ( .A(n5293), .B(n4625), .Z(n2672) );
  ND3 U18348 ( .A(n2610), .B(n2609), .C(n2608), .Z(n1941) );
  ND2 U18349 ( .A(n5290), .B(n4892), .Z(n2609) );
  ND2 U18350 ( .A(n4623), .B(n5290), .Z(n2610) );
  ND2 U18351 ( .A(n4623), .B(n4892), .Z(n2608) );
  ND2 U18352 ( .A(n2084), .B(n4452), .Z(n1454) );
  ND2 U18353 ( .A(n5271), .B(n4910), .Z(n2084) );
  ND2 U18354 ( .A(n3503), .B(n3502), .Z(n1450) );
  ND2 U18355 ( .A(n4779), .B(n5119), .Z(n3503) );
  ND2 U18356 ( .A(n4571), .B(n5119), .Z(n3502) );
  ND2 U18357 ( .A(n4956), .B(n4436), .Z(n3173) );
  ND2 U18358 ( .A(n2391), .B(n2390), .Z(n1937) );
  ND2 U18359 ( .A(n4977), .B(n5141), .Z(n2390) );
  MUX21L U18360 ( .A(n5141), .B(n2389), .S(n4636), .Z(n2391) );
  NR2 U18361 ( .A(n4977), .B(n5141), .Z(n2389) );
  ND2 U18362 ( .A(n4592), .B(n5220), .Z(n1939) );
  ND2 U18363 ( .A(n2700), .B(n2699), .Z(n1405) );
  ND2 U18364 ( .A(n2696), .B(n5294), .Z(n2699) );
  MUX21L U18365 ( .A(n2697), .B(n2698), .S(n4557), .Z(n2700) );
  NR2 U18366 ( .A(n4907), .B(n4557), .Z(n2696) );
  ND2 U18367 ( .A(n2676), .B(n2675), .Z(n1404) );
  MUX21L U18368 ( .A(n2673), .B(n2674), .S(n5293), .Z(n2676) );
  ND2 U18369 ( .A(n2672), .B(n4969), .Z(n2675) );
  NR2 U18370 ( .A(n4969), .B(n4511), .Z(n2673) );
  ND2 U18371 ( .A(n2456), .B(n2455), .Z(n1400) );
  ND2 U18372 ( .A(n2452), .B(n5138), .Z(n2455) );
  MUX21L U18373 ( .A(n2453), .B(n2454), .S(n4915), .Z(n2456) );
  NR2 U18374 ( .A(n4616), .B(n4915), .Z(n2452) );
  ND2 U18375 ( .A(n2487), .B(n2486), .Z(n1401) );
  MUX21L U18376 ( .A(n2484), .B(n2485), .S(n5263), .Z(n2486) );
  MUX21L U18377 ( .A(n2482), .B(n2483), .S(n4917), .Z(n2487) );
  NR2 U18378 ( .A(n4593), .B(n4760), .Z(n2485) );
  ND2 U18379 ( .A(n2292), .B(n2291), .Z(n1395) );
  ND2 U18380 ( .A(n4630), .B(n5152), .Z(n2291) );
  EO U18381 ( .A(n4900), .B(n4630), .Z(n2292) );
  ND2 U18382 ( .A(n3568), .B(n3567), .Z(n1417) );
  ND2 U18383 ( .A(n5248), .B(n4773), .Z(n3567) );
  MUX21L U18384 ( .A(n4773), .B(n3566), .S(n4575), .Z(n3568) );
  NR2 U18385 ( .A(n5248), .B(n4772), .Z(n3566) );
  MUX21L U18386 ( .A(n2943), .B(n2942), .S(n4947), .Z(n1473) );
  ND2 U18387 ( .A(n4547), .B(n5183), .Z(n2942) );
  ND2 U18388 ( .A(n5285), .B(n4548), .Z(n2943) );
  MUX21L U18389 ( .A(n3241), .B(n3240), .S(n4613), .Z(n1480) );
  ND2 U18390 ( .A(n5251), .B(n4952), .Z(n3241) );
  ND2 U18391 ( .A(n4952), .B(n5079), .Z(n3240) );
  MUX21L U18392 ( .A(n3534), .B(n4419), .S(n4923), .Z(n1484) );
  ND2 U18393 ( .A(n4419), .B(n5124), .Z(n3534) );
  MUX21L U18394 ( .A(n3200), .B(n4835), .S(n5230), .Z(n1479) );
  ND2 U18395 ( .A(n4434), .B(n4836), .Z(n3200) );
  MUX21L U18396 ( .A(n2173), .B(n2172), .S(n4967), .Z(n1457) );
  ND2 U18397 ( .A(n4462), .B(n5163), .Z(n2173) );
  ND2 U18398 ( .A(n4597), .B(n5162), .Z(n2172) );
  MUX21L U18399 ( .A(n2315), .B(n2314), .S(n4631), .Z(n1425) );
  ND2 U18400 ( .A(n4961), .B(n5148), .Z(n2314) );
  ND2 U18401 ( .A(n5261), .B(n4961), .Z(n2315) );
  MUX21L U18402 ( .A(n5097), .B(n4821), .S(n4579), .Z(n1441) );
  MUX21L U18403 ( .A(n4549), .B(n2944), .S(n5285), .Z(n1440) );
  ND2 U18404 ( .A(n4548), .B(n4805), .Z(n2944) );
  MUX21L U18405 ( .A(n2533), .B(n2532), .S(n4975), .Z(n1431) );
  ND2 U18406 ( .A(n5288), .B(n4619), .Z(n2533) );
  ND2 U18407 ( .A(n4619), .B(n5217), .Z(n2532) );
  MUX21L U18408 ( .A(n4882), .B(n4637), .S(n5265), .Z(n1428) );
  MUX21L U18409 ( .A(n3333), .B(n3332), .S(n4607), .Z(n1954) );
  ND2 U18410 ( .A(n4796), .B(n5103), .Z(n3332) );
  ND2 U18411 ( .A(n5256), .B(n4934), .Z(n3333) );
  MUX21L U18412 ( .A(n5076), .B(n3283), .S(n4610), .Z(n1953) );
  ND2 U18413 ( .A(n4843), .B(n5076), .Z(n3283) );
  MUX21L U18414 ( .A(n4766), .B(n5165), .S(n4599), .Z(n1930) );
  MUX21L U18415 ( .A(n4878), .B(n4535), .S(n5262), .Z(n1934) );
  MUX21L U18416 ( .A(n4962), .B(n4540), .S(n5260), .Z(n1933) );
  MUX21L U18417 ( .A(n2896), .B(n5284), .S(n4566), .Z(n2898) );
  NR2 U18418 ( .A(n5284), .B(n4799), .Z(n2896) );
  IVP U18419 ( .A(n4360), .Z(n4632) );
  IVP U18420 ( .A(n5061), .Z(n5276) );
  IVP U18421 ( .A(n4728), .Z(n4935) );
  IVP U18422 ( .A(n5064), .Z(n5257) );
  IVP U18423 ( .A(n4731), .Z(n4918) );
  IVP U18424 ( .A(n5066), .Z(n5247) );
  IVP U18425 ( .A(n5062), .Z(n5270) );
  IVP U18426 ( .A(n4732), .Z(n4909) );
  IVP U18427 ( .A(n5065), .Z(n5253) );
  IVP U18428 ( .A(n4723), .Z(n4966) );
  IVP U18429 ( .A(n5066), .Z(n5248) );
  IVP U18430 ( .A(n4365), .Z(n4605) );
  NR2 U18431 ( .A(n5294), .B(n4907), .Z(n2698) );
  NR2 U18432 ( .A(n5267), .B(n4527), .Z(n2454) );
  NR2 U18433 ( .A(n5286), .B(n4474), .Z(n2483) );
  NR2 U18434 ( .A(n5257), .B(n4793), .Z(n3345) );
  NR2 U18435 ( .A(n4571), .B(n5120), .Z(n1416) );
  NR2 U18436 ( .A(n4918), .B(n4430), .Z(n1415) );
  ND2 U18437 ( .A(n4468), .B(n5159), .Z(n2230) );
  ND2 U18438 ( .A(n4468), .B(n4865), .Z(n2231) );
  ND2 U18439 ( .A(n4866), .B(n5159), .Z(n2232) );
  ND2 U18440 ( .A(n4593), .B(n5156), .Z(n1458) );
  ND2 U18441 ( .A(n3261), .B(n3260), .Z(n1920) );
  MUX21L U18442 ( .A(n3258), .B(n3259), .S(n4951), .Z(n3260) );
  MUX21L U18443 ( .A(n3256), .B(n3257), .S(n5252), .Z(n3261) );
  NR2 U18444 ( .A(n4612), .B(n5078), .Z(n3258) );
  ND2 U18445 ( .A(n3381), .B(n3380), .Z(n1922) );
  MUX21L U18446 ( .A(n3378), .B(n3379), .S(n4936), .Z(n3380) );
  MUX21L U18447 ( .A(n3376), .B(n3377), .S(n5258), .Z(n3381) );
  NR2 U18448 ( .A(n4604), .B(n5107), .Z(n3378) );
  ND2 U18449 ( .A(n4472), .B(n5155), .Z(n2257) );
  ND2 U18450 ( .A(n5264), .B(n4881), .Z(n1936) );
  ND2 U18451 ( .A(n2535), .B(n2534), .Z(n1402) );
  ND2 U18452 ( .A(n5288), .B(n4525), .Z(n2534) );
  EN U18453 ( .A(n5226), .B(n4975), .Z(n2535) );
  AN3 U18454 ( .A(n4480), .B(n5078), .C(n4952), .Z(n769) );
  MUX21L U18455 ( .A(n2052), .B(n2051), .S(n4909), .Z(n1390) );
  ND2 U18456 ( .A(n5270), .B(n4627), .Z(n2052) );
  ND2 U18457 ( .A(n4627), .B(n5174), .Z(n2051) );
  MUX21L U18458 ( .A(n2093), .B(n4911), .S(n4602), .Z(n1391) );
  ND2 U18459 ( .A(n4911), .B(n5169), .Z(n2093) );
  MUX21L U18460 ( .A(n2036), .B(n2035), .S(n5269), .Z(n1389) );
  ND2 U18461 ( .A(n4445), .B(n4859), .Z(n2036) );
  ND2 U18462 ( .A(n4958), .B(n4445), .Z(n2035) );
  MUX21L U18463 ( .A(n3201), .B(n5083), .S(n4954), .Z(n1412) );
  ND2 U18464 ( .A(n4587), .B(n5083), .Z(n3201) );
  IVP U18465 ( .A(n4725), .Z(n4950) );
  IVP U18466 ( .A(n4730), .Z(n4921) );
  IVP U18467 ( .A(n4369), .Z(n4555) );
  IVP U18468 ( .A(n4359), .Z(n4637) );
  IVP U18469 ( .A(n5068), .Z(n5232) );
  IVP U18470 ( .A(n4372), .Z(n4572) );
  NR2 U18471 ( .A(n4951), .B(n4482), .Z(n3256) );
  NR2 U18472 ( .A(n4936), .B(n4468), .Z(n3376) );
  NR2 U18473 ( .A(n5269), .B(n4446), .Z(n2040) );
  NR2 U18474 ( .A(n4627), .B(n4858), .Z(n2042) );
  NR2 U18475 ( .A(n4558), .B(n4754), .Z(n2720) );
  NR2 U18476 ( .A(n5245), .B(n4422), .Z(n3505) );
  NR2 U18477 ( .A(n4958), .B(n5091), .Z(n3142) );
  NR2 U18478 ( .A(n5294), .B(n4755), .Z(n2697) );
  ND2 U18479 ( .A(n4950), .B(n5076), .Z(n3284) );
  ND2 U18480 ( .A(n4950), .B(n4486), .Z(n3285) );
  ND2 U18481 ( .A(n4629), .B(n5153), .Z(n2268) );
  ND2 U18482 ( .A(n3597), .B(n3596), .Z(n1925) );
  ND2 U18483 ( .A(n4411), .B(n4769), .Z(n3596) );
  EO U18484 ( .A(n5227), .B(n4926), .Z(n3597) );
  ND2 U18485 ( .A(n2031), .B(n2030), .Z(n1891) );
  ND2 U18486 ( .A(n4968), .B(n4543), .Z(n2030) );
  MUX21L U18487 ( .A(n5175), .B(n2029), .S(n4628), .Z(n2031) );
  NR2 U18488 ( .A(n4968), .B(n5175), .Z(n2029) );
  ND2 U18489 ( .A(n2196), .B(n2195), .Z(n1895) );
  ND2 U18490 ( .A(n4596), .B(n4864), .Z(n2195) );
  EO U18491 ( .A(n5230), .B(n4967), .Z(n2196) );
  ND2 U18492 ( .A(n2786), .B(n2785), .Z(n1910) );
  ND2 U18493 ( .A(n4495), .B(n4743), .Z(n2785) );
  EO U18494 ( .A(n5223), .B(n4561), .Z(n2786) );
  ND2 U18495 ( .A(n3055), .B(n3054), .Z(n1915) );
  ND2 U18496 ( .A(n4555), .B(n4818), .Z(n3054) );
  MUX21L U18497 ( .A(n3053), .B(n5232), .S(n4555), .Z(n3055) );
  NR2 U18498 ( .A(n5231), .B(n4818), .Z(n3053) );
  ND2 U18499 ( .A(n2892), .B(n2891), .Z(n1912) );
  MUX21L U18500 ( .A(n2889), .B(n2890), .S(n5284), .Z(n2892) );
  ND2 U18501 ( .A(n2888), .B(n4933), .Z(n2891) );
  NR2 U18502 ( .A(n4933), .B(n4399), .Z(n2889) );
  ND2 U18503 ( .A(n2722), .B(n2721), .Z(n1909) );
  MUX21L U18504 ( .A(n2719), .B(n2720), .S(n5295), .Z(n2721) );
  MUX21L U18505 ( .A(n2717), .B(n2718), .S(n4907), .Z(n2722) );
  NR2 U18506 ( .A(n4907), .B(n4558), .Z(n2719) );
  ND2 U18507 ( .A(n3124), .B(n4376), .Z(n1916) );
  EO U18508 ( .A(n5224), .B(n4938), .Z(n3124) );
  ND2 U18509 ( .A(n2637), .B(n2636), .Z(n1905) );
  ND2 U18510 ( .A(n4624), .B(n4971), .Z(n2636) );
  MUX21L U18511 ( .A(n2635), .B(n5210), .S(n4971), .Z(n2637) );
  NR2 U18512 ( .A(n4624), .B(n5209), .Z(n2635) );
  ND2 U18513 ( .A(n2583), .B(n4889), .Z(n1904) );
  ND2 U18514 ( .A(n5290), .B(n4621), .Z(n2583) );
  ND2 U18515 ( .A(n4437), .B(n5088), .Z(n3174) );
  ND2 U18516 ( .A(n2375), .B(n2374), .Z(n1364) );
  ND2 U18517 ( .A(n4880), .B(n5143), .Z(n2374) );
  MUX21L U18518 ( .A(n5144), .B(n2373), .S(n4635), .Z(n2375) );
  MUX21L U18519 ( .A(n3167), .B(n4439), .S(n4956), .Z(n1918) );
  ND2 U18520 ( .A(n5233), .B(n4439), .Z(n3167) );
  MUX21L U18521 ( .A(n3401), .B(n5241), .S(n4588), .Z(n1923) );
  ND2 U18522 ( .A(n5241), .B(n4789), .Z(n3401) );
  MUX21L U18523 ( .A(n2234), .B(n2233), .S(n4595), .Z(n1896) );
  ND2 U18524 ( .A(n5276), .B(n4866), .Z(n2233) );
  ND2 U18525 ( .A(n4965), .B(n5276), .Z(n2234) );
  MUX21L U18526 ( .A(n2130), .B(n2129), .S(n4600), .Z(n1894) );
  ND2 U18527 ( .A(n4850), .B(n5167), .Z(n2129) );
  ND2 U18528 ( .A(n5273), .B(n4851), .Z(n2130) );
  MUX21L U18529 ( .A(n4388), .B(n5086), .S(n4945), .Z(n1914) );
  MUX21L U18530 ( .A(n2690), .B(n2689), .S(n4556), .Z(n1907) );
  ND2 U18531 ( .A(n5294), .B(n4756), .Z(n2689) );
  ND2 U18532 ( .A(n4906), .B(n5294), .Z(n2690) );
  MUX21L U18533 ( .A(n2678), .B(n4510), .S(n4969), .Z(n1906) );
  ND2 U18534 ( .A(n4510), .B(n5206), .Z(n2678) );
  ND2 U18535 ( .A(n3245), .B(n3244), .Z(n1383) );
  ND3 U18536 ( .A(n4952), .B(n4480), .C(n5251), .Z(n3244) );
  MUX21L U18537 ( .A(n3242), .B(n3243), .S(n4952), .Z(n3245) );
  NR2 U18538 ( .A(n5252), .B(n4480), .Z(n3243) );
  IVP U18539 ( .A(n4363), .Z(n4614) );
  IVP U18540 ( .A(n4371), .Z(n4567) );
  IVP U18541 ( .A(n4725), .Z(n4955) );
  AO7 U18542 ( .A(n4916), .B(n5135), .C(n4526), .Z(n1902) );
  NR2 U18543 ( .A(n5291), .B(n4504), .Z(n2718) );
  NR2 U18544 ( .A(n4614), .B(n4883), .Z(n2408) );
  ND3 U18545 ( .A(n4617), .B(n5136), .C(n4916), .Z(n1366) );
  ND3 U18546 ( .A(n2795), .B(n2794), .C(n2793), .Z(n1374) );
  ND2 U18547 ( .A(n5280), .B(n4494), .Z(n2794) );
  ND2 U18548 ( .A(n4929), .B(n5279), .Z(n2795) );
  ND2 U18549 ( .A(n4929), .B(n4495), .Z(n2793) );
  ND2 U18550 ( .A(n4425), .B(n4781), .Z(n1483) );
  ND2 U18551 ( .A(n5232), .B(n4393), .Z(n1913) );
  ND2 U18552 ( .A(n4635), .B(n5145), .Z(n1900) );
  MUX21L U18553 ( .A(n2564), .B(n2563), .S(n5289), .Z(n1869) );
  ND2 U18554 ( .A(n4524), .B(n4887), .Z(n2564) );
  ND2 U18555 ( .A(n4974), .B(n4620), .Z(n2563) );
  ND2 U18556 ( .A(n4532), .B(n4880), .Z(n2372) );
  ND2 U18557 ( .A(n2206), .B(n2205), .Z(n1359) );
  ND2 U18558 ( .A(n4596), .B(n4865), .Z(n2205) );
  EO U18559 ( .A(n5230), .B(n4596), .Z(n2206) );
  ND2 U18560 ( .A(n2119), .B(n2118), .Z(n1357) );
  ND2 U18561 ( .A(n4457), .B(n4851), .Z(n2118) );
  EO U18562 ( .A(n5229), .B(n4601), .Z(n2119) );
  ND2 U18563 ( .A(n2279), .B(n2278), .Z(n1361) );
  ND2 U18564 ( .A(n4629), .B(n4871), .Z(n2278) );
  MUX21L U18565 ( .A(n5259), .B(n2277), .S(n4963), .Z(n2279) );
  NR2 U18566 ( .A(n5259), .B(n4629), .Z(n2277) );
  ND2 U18567 ( .A(n2054), .B(n2053), .Z(n1356) );
  ND2 U18568 ( .A(n5270), .B(n4448), .Z(n2054) );
  ND2 U18569 ( .A(n5270), .B(n4857), .Z(n2053) );
  ND2 U18570 ( .A(n2912), .B(n5185), .Z(n1376) );
  EO U18571 ( .A(n4901), .B(n4567), .Z(n2912) );
  ND2 U18572 ( .A(n2828), .B(n2827), .Z(n1375) );
  ND2 U18573 ( .A(n4405), .B(n4738), .Z(n2828) );
  ND2 U18574 ( .A(n5281), .B(n4404), .Z(n2827) );
  MUX21L U18575 ( .A(n5212), .B(n2599), .S(n4973), .Z(n1369) );
  ND2 U18576 ( .A(n4622), .B(n5213), .Z(n2599) );
  MUX21L U18577 ( .A(n4754), .B(n5203), .S(n4557), .Z(n1371) );
  MUX21L U18578 ( .A(n2946), .B(n2945), .S(n5286), .Z(n1377) );
  ND2 U18579 ( .A(n4947), .B(n4395), .Z(n2946) );
  ND2 U18580 ( .A(n4548), .B(n4806), .Z(n2945) );
  MUX21L U18581 ( .A(n3090), .B(n3089), .S(n4580), .Z(n1380) );
  ND2 U18582 ( .A(n5238), .B(n4823), .Z(n3089) );
  ND2 U18583 ( .A(n4940), .B(n5238), .Z(n3090) );
  IVP U18584 ( .A(n4372), .Z(n4574) );
  IVP U18585 ( .A(n4727), .Z(n4942) );
  AO7 U18586 ( .A(n4591), .B(n5219), .C(n4758), .Z(n1903) );
  ND2 U18587 ( .A(n2726), .B(n2725), .Z(n1873) );
  MUX21L U18588 ( .A(n2723), .B(n5202), .S(n4558), .Z(n2725) );
  AO6 U18589 ( .A(n4558), .B(n4753), .C(n2724), .Z(n2726) );
  AO7 U18590 ( .A(n4920), .B(n5116), .C(n4426), .Z(n1386) );
  ND2 U18591 ( .A(n2692), .B(n2691), .Z(n1871) );
  ND2 U18592 ( .A(n4906), .B(n4508), .Z(n2691) );
  EN U18593 ( .A(n5225), .B(n4556), .Z(n2692) );
  ND2 U18594 ( .A(n3481), .B(n3480), .Z(n1888) );
  ND2 U18595 ( .A(n4424), .B(n5117), .Z(n3480) );
  EN U18596 ( .A(n4900), .B(n4569), .Z(n3481) );
  ND2 U18597 ( .A(n3263), .B(n3262), .Z(n1884) );
  ND2 U18598 ( .A(n4612), .B(n4842), .Z(n3262) );
  EO U18599 ( .A(n5225), .B(n4612), .Z(n3263) );
  ND2 U18600 ( .A(n3314), .B(n3313), .Z(n1885) );
  ND2 U18601 ( .A(n4608), .B(n4848), .Z(n3313) );
  EO U18602 ( .A(n5224), .B(n4948), .Z(n3314) );
  ND2 U18603 ( .A(n2290), .B(n4872), .Z(n1863) );
  EN U18604 ( .A(n5222), .B(n4630), .Z(n2290) );
  ND3 U18605 ( .A(n4796), .B(n5102), .C(n4490), .Z(n1413) );
  MUX21L U18606 ( .A(n4554), .B(n3036), .S(n4943), .Z(n1879) );
  ND2 U18607 ( .A(n4554), .B(n5101), .Z(n3036) );
  MUX21L U18608 ( .A(n2811), .B(n2810), .S(n4562), .Z(n1875) );
  ND2 U18609 ( .A(n4740), .B(n5193), .Z(n2810) );
  ND2 U18610 ( .A(n4930), .B(n5193), .Z(n2811) );
  MUX21L U18611 ( .A(n2987), .B(n2986), .S(n4551), .Z(n1878) );
  ND2 U18612 ( .A(n4809), .B(n5179), .Z(n2986) );
  ND2 U18613 ( .A(n5233), .B(n4809), .Z(n2987) );
  MUX21L U18614 ( .A(n3126), .B(n3125), .S(n4582), .Z(n1882) );
  ND2 U18615 ( .A(n4938), .B(n5238), .Z(n3126) );
  ND2 U18616 ( .A(n5238), .B(n4826), .Z(n3125) );
  MUX21L U18617 ( .A(n4968), .B(n2032), .S(n5269), .Z(n1857) );
  ND2 U18618 ( .A(n4968), .B(n4518), .Z(n2032) );
  ND2 U18619 ( .A(n2236), .B(n2235), .Z(n1862) );
  ND2 U18620 ( .A(n4469), .B(n5158), .Z(n2236) );
  ND2 U18621 ( .A(n4965), .B(n5158), .Z(n2235) );
  ND2 U18622 ( .A(n4553), .B(n4815), .Z(n1378) );
  ND2 U18623 ( .A(n2069), .B(n2068), .Z(n1858) );
  ND2 U18624 ( .A(n4910), .B(n5271), .Z(n2068) );
  MUX21L U18625 ( .A(n2067), .B(n4451), .S(n5271), .Z(n2069) );
  NR2 U18626 ( .A(n4910), .B(n4451), .Z(n2067) );
  ND2 U18627 ( .A(n2097), .B(n2096), .Z(n1325) );
  MUX21L U18628 ( .A(n2094), .B(n5169), .S(n4911), .Z(n2096) );
  AO6 U18629 ( .A(n4911), .B(n4455), .C(n2095), .Z(n2097) );
  IVP U18630 ( .A(n4366), .Z(n4598) );
  AO7 U18631 ( .A(n4913), .B(n5167), .C(n4458), .Z(n1859) );
  NR2 U18632 ( .A(n4631), .B(n4873), .Z(n1864) );
  ND3 U18633 ( .A(n4588), .B(n4837), .C(n5250), .Z(n1883) );
  ND2 U18634 ( .A(n4968), .B(n5184), .Z(n2925) );
  ND2 U18635 ( .A(n4968), .B(n4396), .Z(n2926) );
  ND2 U18636 ( .A(n4920), .B(n4427), .Z(n1887) );
  ND2 U18637 ( .A(n2132), .B(n2131), .Z(n1860) );
  ND2 U18638 ( .A(n4459), .B(n4850), .Z(n2132) );
  ND2 U18639 ( .A(n5273), .B(n4459), .Z(n2131) );
  ND2 U18640 ( .A(n3416), .B(n3415), .Z(n1352) );
  MUX21L U18641 ( .A(n3413), .B(n3414), .S(n4589), .Z(n3416) );
  ND2 U18642 ( .A(n3412), .B(n5242), .Z(n3415) );
  NR2 U18643 ( .A(n5242), .B(n4788), .Z(n3413) );
  MUX21L U18644 ( .A(n3301), .B(n3300), .S(n4949), .Z(n1350) );
  ND2 U18645 ( .A(n5255), .B(n4488), .Z(n3301) );
  ND2 U18646 ( .A(n4609), .B(n5074), .Z(n3300) );
  MUX21L U18647 ( .A(n2649), .B(n5292), .S(n4624), .Z(n1336) );
  ND2 U18648 ( .A(n5292), .B(n4971), .Z(n2649) );
  AO7 U18649 ( .A(n4552), .B(n4814), .C(n3015), .Z(n1343) );
  ND2 U18650 ( .A(n5239), .B(n4944), .Z(n3015) );
  MUX21L U18651 ( .A(n2839), .B(n2838), .S(n5282), .Z(n1341) );
  ND2 U18652 ( .A(n4931), .B(n4404), .Z(n2839) );
  ND2 U18653 ( .A(n4931), .B(n4564), .Z(n2838) );
  ND2 U18654 ( .A(n4632), .B(n4875), .Z(n2316) );
  AN3 U18655 ( .A(n4571), .B(n5120), .C(n4921), .Z(n770) );
  ND2 U18656 ( .A(n3204), .B(n3203), .Z(n1348) );
  ND2 U18657 ( .A(n4836), .B(n5082), .Z(n3203) );
  MUX21L U18658 ( .A(n5083), .B(n3202), .S(n4587), .Z(n3204) );
  ND2 U18659 ( .A(n2470), .B(n2469), .Z(n1332) );
  ND2 U18660 ( .A(n4761), .B(n5136), .Z(n2469) );
  MUX21L U18661 ( .A(n5136), .B(n2468), .S(n4618), .Z(n2470) );
  ND2 U18662 ( .A(n2704), .B(n2703), .Z(n1337) );
  ND3 U18663 ( .A(n4907), .B(n4508), .C(n5295), .Z(n2703) );
  MUX21L U18664 ( .A(n2701), .B(n2702), .S(n4907), .Z(n2704) );
  NR2 U18665 ( .A(n5295), .B(n4507), .Z(n2702) );
  IVP U18666 ( .A(n5060), .Z(n5282) );
  IVP U18667 ( .A(n4375), .Z(n4589) );
  IVP U18668 ( .A(n5067), .Z(n5242) );
  IVP U18669 ( .A(n4367), .Z(n4594) );
  IVP U18670 ( .A(n4726), .Z(n4949) );
  IVP U18671 ( .A(n5068), .Z(n5236) );
  AO6 U18672 ( .A(n4967), .B(n4463), .C(n2176), .Z(n2178) );
  NR2 U18673 ( .A(n5274), .B(n4597), .Z(n2176) );
  AO7 U18674 ( .A(n4561), .B(n4742), .C(n5194), .Z(n1340) );
  NR2 U18675 ( .A(n5284), .B(n4735), .Z(n1342) );
  ND2 U18676 ( .A(n3038), .B(n3037), .Z(n1845) );
  ND2 U18677 ( .A(n4385), .B(n5101), .Z(n3037) );
  EN U18678 ( .A(n4897), .B(n4554), .Z(n3038) );
  ND2 U18679 ( .A(n3103), .B(n3102), .Z(n1846) );
  ND2 U18680 ( .A(n4939), .B(n4377), .Z(n3102) );
  EO U18681 ( .A(n5223), .B(n4581), .Z(n3103) );
  ND2 U18682 ( .A(n2584), .B(n4889), .Z(n1835) );
  EO U18683 ( .A(n5226), .B(n4621), .Z(n2584) );
  ND2 U18684 ( .A(n2273), .B(n2272), .Z(n1828) );
  ND2 U18685 ( .A(n2269), .B(n5153), .Z(n2272) );
  MUX21L U18686 ( .A(n2270), .B(n2271), .S(n4963), .Z(n2273) );
  NR2 U18687 ( .A(n4629), .B(n4963), .Z(n2269) );
  ND2 U18688 ( .A(n2615), .B(n2614), .Z(n1836) );
  ND2 U18689 ( .A(n2611), .B(n5291), .Z(n2614) );
  MUX21L U18690 ( .A(n2612), .B(n2613), .S(n5291), .Z(n2615) );
  NR2 U18691 ( .A(n4972), .B(n4623), .Z(n2611) );
  ND2 U18692 ( .A(n3484), .B(n3483), .Z(n1854) );
  ND2 U18693 ( .A(n4920), .B(n5117), .Z(n3483) );
  MUX21L U18694 ( .A(n5117), .B(n3482), .S(n4569), .Z(n3484) );
  NR2 U18695 ( .A(n4920), .B(n5118), .Z(n3482) );
  MUX21L U18696 ( .A(n2175), .B(n5161), .S(n4967), .Z(n2177) );
  MUX21L U18697 ( .A(n3076), .B(n4381), .S(n4941), .Z(n1344) );
  ND2 U18698 ( .A(n4382), .B(n5097), .Z(n3076) );
  ND2 U18699 ( .A(n2567), .B(n2566), .Z(n1304) );
  ND2 U18700 ( .A(n4887), .B(n5215), .Z(n2566) );
  MUX21L U18701 ( .A(n4887), .B(n2565), .S(n4620), .Z(n2567) );
  IVP U18702 ( .A(n4724), .Z(n4957) );
  IVP U18703 ( .A(n4360), .Z(n4633) );
  IVP U18704 ( .A(n5068), .Z(n5234) );
  IVP U18705 ( .A(n4722), .Z(n4972) );
  AO7 U18706 ( .A(n4587), .B(n4835), .C(n5085), .Z(n1849) );
  NR2 U18707 ( .A(n5259), .B(n4542), .Z(n2271) );
  NR2 U18708 ( .A(n4972), .B(n4518), .Z(n2612) );
  NR2 U18709 ( .A(n4960), .B(n5147), .Z(n2326) );
  NR2 U18710 ( .A(n4960), .B(n4537), .Z(n2327) );
  MUX21L U18711 ( .A(n2325), .B(n4632), .S(n5261), .Z(n2328) );
  NR2 U18712 ( .A(n4633), .B(n4876), .Z(n2325) );
  ND3 U18713 ( .A(n2311), .B(n2310), .C(n2309), .Z(n1829) );
  ND2 U18714 ( .A(n4538), .B(n5149), .Z(n2310) );
  ND2 U18715 ( .A(n4961), .B(n5149), .Z(n2311) );
  ND2 U18716 ( .A(n4961), .B(n4538), .Z(n2309) );
  ND3 U18717 ( .A(n2814), .B(n2813), .C(n2812), .Z(n1841) );
  ND2 U18718 ( .A(n4407), .B(n4740), .Z(n2813) );
  ND2 U18719 ( .A(n5280), .B(n4740), .Z(n2814) );
  ND2 U18720 ( .A(n5280), .B(n4407), .Z(n2812) );
  ND2 U18721 ( .A(n4565), .B(n5189), .Z(n2860) );
  ND2 U18722 ( .A(n5283), .B(n4402), .Z(n2861) );
  MUX21L U18723 ( .A(n2800), .B(n4409), .S(n4929), .Z(n1840) );
  ND2 U18724 ( .A(n5280), .B(n4493), .Z(n2800) );
  AO7 U18725 ( .A(n4976), .B(n4530), .C(n2406), .Z(n1832) );
  ND2 U18726 ( .A(n5265), .B(n4637), .Z(n2406) );
  MUX21L U18727 ( .A(n4610), .B(n3286), .S(n5254), .Z(n1851) );
  ND2 U18728 ( .A(n4610), .B(n4843), .Z(n3286) );
  MUX21L U18729 ( .A(n4838), .B(n3220), .S(n4614), .Z(n1850) );
  ND2 U18730 ( .A(n5251), .B(n4838), .Z(n3220) );
  MUX21L U18731 ( .A(n3403), .B(n3402), .S(n4937), .Z(n1853) );
  ND2 U18732 ( .A(n4431), .B(n5110), .Z(n3402) );
  ND2 U18733 ( .A(n5242), .B(n4431), .Z(n3403) );
  ND2 U18734 ( .A(n4380), .B(n5095), .Z(n3082) );
  AO7 U18735 ( .A(n4905), .B(n4505), .C(n2711), .Z(n1307) );
  ND2 U18736 ( .A(n5295), .B(n4557), .Z(n2711) );
  AN3 U18737 ( .A(n4444), .B(n5174), .C(n4968), .Z(n771) );
  MUX21L U18738 ( .A(n4856), .B(n5171), .S(n4626), .Z(n1823) );
  ND2 U18739 ( .A(n2729), .B(n2728), .Z(n1839) );
  ND2 U18740 ( .A(n4558), .B(n5202), .Z(n2728) );
  MUX21L U18741 ( .A(n4753), .B(n2727), .S(n5277), .Z(n2729) );
  NR2 U18742 ( .A(n4558), .B(n4753), .Z(n2727) );
  MUX21L U18743 ( .A(n5203), .B(n4505), .S(n4907), .Z(n1837) );
  MUX21L U18744 ( .A(n5264), .B(n4882), .S(n4635), .Z(n1831) );
  MUX21L U18745 ( .A(n4957), .B(n4440), .S(n5234), .Z(n1848) );
  ND2 U18746 ( .A(n3147), .B(n3146), .Z(n1318) );
  ND2 U18747 ( .A(n5236), .B(n4829), .Z(n3146) );
  MUX21L U18748 ( .A(n4829), .B(n3145), .S(n4584), .Z(n3147) );
  NR2 U18749 ( .A(n5236), .B(n4828), .Z(n3145) );
  IVP U18750 ( .A(n4364), .Z(n4611) );
  ND2 U18751 ( .A(n2865), .B(n2864), .Z(n1809) );
  MUX21L U18752 ( .A(n5283), .B(n2862), .S(n4932), .Z(n2864) );
  AO6 U18753 ( .A(n5283), .B(n4401), .C(n2863), .Z(n2865) );
  NR2 U18754 ( .A(n5283), .B(n4401), .Z(n2862) );
  ND3 U18755 ( .A(n2745), .B(n2744), .C(n2743), .Z(n1339) );
  ND2 U18756 ( .A(n4750), .B(n5199), .Z(n2745) );
  ND2 U18757 ( .A(n4503), .B(n4750), .Z(n2744) );
  ND2 U18758 ( .A(n4503), .B(n5200), .Z(n2743) );
  ND3 U18759 ( .A(n2949), .B(n2948), .C(n2947), .Z(n1313) );
  ND2 U18760 ( .A(n4806), .B(n5183), .Z(n2948) );
  ND2 U18761 ( .A(n4547), .B(n4806), .Z(n2947) );
  ND2 U18762 ( .A(n4548), .B(n5183), .Z(n2949) );
  ND2 U18763 ( .A(n4533), .B(n5146), .Z(n2359) );
  MUX21L U18764 ( .A(n2630), .B(n2629), .S(n5291), .Z(n1305) );
  ND2 U18765 ( .A(n4517), .B(n4893), .Z(n2630) );
  ND2 U18766 ( .A(n4971), .B(n4623), .Z(n2629) );
  ND2 U18767 ( .A(n4611), .B(n5077), .Z(n3264) );
  ND2 U18768 ( .A(n5242), .B(n4788), .Z(n3417) );
  ND2 U18769 ( .A(n5242), .B(n4429), .Z(n3418) );
  MUX21L U18770 ( .A(n2876), .B(n2875), .S(n4565), .Z(n1312) );
  ND2 U18771 ( .A(n5284), .B(n4785), .Z(n2875) );
  ND2 U18772 ( .A(n4933), .B(n5284), .Z(n2876) );
  ND2 U18773 ( .A(n2771), .B(n2770), .Z(n1310) );
  ND2 U18774 ( .A(n4747), .B(n5195), .Z(n2771) );
  ND2 U18775 ( .A(n4560), .B(n4747), .Z(n2770) );
  ND2 U18776 ( .A(n2747), .B(n2746), .Z(n1309) );
  ND2 U18777 ( .A(n4502), .B(n5199), .Z(n2747) );
  ND2 U18778 ( .A(n4905), .B(n4502), .Z(n2746) );
  ND2 U18779 ( .A(n3030), .B(n4387), .Z(n1314) );
  ND2 U18780 ( .A(n5240), .B(n4943), .Z(n3030) );
  IVP U18781 ( .A(n5066), .Z(n5246) );
  IVP U18782 ( .A(n4724), .Z(n4959) );
  IVP U18783 ( .A(n4726), .Z(n4946) );
  IVP U18784 ( .A(n4730), .Z(n4922) );
  NR2 U18785 ( .A(n5288), .B(n4884), .Z(n2538) );
  ND2 U18786 ( .A(n2350), .B(n2349), .Z(n1796) );
  ND2 U18787 ( .A(n4633), .B(n5146), .Z(n2349) );
  EO U18788 ( .A(n5222), .B(n4959), .Z(n2350) );
  ND2 U18789 ( .A(n2474), .B(n2473), .Z(n1800) );
  ND2 U18790 ( .A(n4618), .B(n5135), .Z(n2473) );
  EO U18791 ( .A(n4898), .B(n4618), .Z(n2474) );
  ND2 U18792 ( .A(n3551), .B(n3550), .Z(n1821) );
  ND2 U18793 ( .A(n4416), .B(n5125), .Z(n3550) );
  EN U18794 ( .A(n4902), .B(n4574), .Z(n3551) );
  ND2 U18795 ( .A(n3218), .B(n4837), .Z(n1816) );
  EO U18796 ( .A(n5229), .B(n4588), .Z(n3218) );
  ND2 U18797 ( .A(n4804), .B(n5184), .Z(n2927) );
  MUX21L U18798 ( .A(n2989), .B(n2988), .S(n4551), .Z(n1811) );
  ND2 U18799 ( .A(n4809), .B(n5178), .Z(n2988) );
  ND2 U18800 ( .A(n5234), .B(n4810), .Z(n2989) );
  MUX21L U18801 ( .A(n2709), .B(n2708), .S(n5295), .Z(n1805) );
  ND2 U18802 ( .A(n4557), .B(n4755), .Z(n2709) );
  ND2 U18803 ( .A(n4908), .B(n4557), .Z(n2708) );
  MUX21L U18804 ( .A(n3335), .B(n3334), .S(n4607), .Z(n1818) );
  ND2 U18805 ( .A(n4796), .B(n5103), .Z(n3334) );
  ND2 U18806 ( .A(n5256), .B(n4934), .Z(n3335) );
  MUX21L U18807 ( .A(n2070), .B(n4452), .S(n5271), .Z(n2072) );
  NR2 U18808 ( .A(n4910), .B(n4451), .Z(n2070) );
  ND2 U18809 ( .A(n2135), .B(n2134), .Z(n1793) );
  ND2 U18810 ( .A(n5273), .B(n4849), .Z(n2134) );
  MUX21L U18811 ( .A(n4850), .B(n2133), .S(n4600), .Z(n2135) );
  NR2 U18812 ( .A(n5273), .B(n4849), .Z(n2133) );
  ND2 U18813 ( .A(n2670), .B(n2669), .Z(n1804) );
  ND2 U18814 ( .A(n4625), .B(n4803), .Z(n2669) );
  MUX21L U18815 ( .A(n2668), .B(n5293), .S(n4625), .Z(n2670) );
  NR2 U18816 ( .A(n5293), .B(n4802), .Z(n2668) );
  ND2 U18817 ( .A(n3436), .B(n3435), .Z(n1819) );
  ND2 U18818 ( .A(n4428), .B(n5113), .Z(n3435) );
  MUX21L U18819 ( .A(n4785), .B(n3434), .S(n4590), .Z(n3436) );
  ND2 U18820 ( .A(n2774), .B(n2773), .Z(n1279) );
  ND2 U18821 ( .A(n5279), .B(n4746), .Z(n2773) );
  MUX21L U18822 ( .A(n2772), .B(n4497), .S(n5279), .Z(n2774) );
  ND2 U18823 ( .A(n2540), .B(n2539), .Z(n1275) );
  ND2 U18824 ( .A(n2536), .B(n5217), .Z(n2539) );
  MUX21L U18825 ( .A(n2537), .B(n2538), .S(n4619), .Z(n2540) );
  NR2 U18826 ( .A(n4619), .B(n4975), .Z(n2536) );
  IVP U18827 ( .A(n4374), .Z(n4586) );
  IVP U18828 ( .A(n4375), .Z(n4590) );
  IVP U18829 ( .A(n4730), .Z(n4925) );
  NR2 U18830 ( .A(n4626), .B(n4856), .Z(n2074) );
  NR2 U18831 ( .A(n4966), .B(n5160), .Z(n2208) );
  NR2 U18832 ( .A(n4966), .B(n4466), .Z(n2209) );
  ND2 U18833 ( .A(n2211), .B(n2210), .Z(n1269) );
  MUX21L U18834 ( .A(n2207), .B(n4596), .S(n5275), .Z(n2210) );
  NR2 U18835 ( .A(n2209), .B(n2208), .Z(n2211) );
  NR2 U18836 ( .A(n4596), .B(n4865), .Z(n2207) );
  ND2 U18837 ( .A(n2121), .B(n2120), .Z(n1267) );
  ND2 U18838 ( .A(n4601), .B(n4851), .Z(n2120) );
  EO U18839 ( .A(n5229), .B(n4601), .Z(n2121) );
  ND2 U18840 ( .A(n3351), .B(n3350), .Z(n1290) );
  ND2 U18841 ( .A(n4491), .B(n5105), .Z(n3350) );
  EN U18842 ( .A(n4897), .B(n4605), .Z(n3351) );
  ND3 U18843 ( .A(n4568), .B(n4782), .C(n5244), .Z(n1291) );
  ND2 U18844 ( .A(n2528), .B(n2527), .Z(n1802) );
  ND2 U18845 ( .A(n4975), .B(n4525), .Z(n2528) );
  ND2 U18846 ( .A(n4975), .B(n5219), .Z(n2527) );
  ND2 U18847 ( .A(n4909), .B(n5173), .Z(n2055) );
  ND2 U18848 ( .A(n4964), .B(n5157), .Z(n2246) );
  ND2 U18849 ( .A(n4964), .B(n4471), .Z(n2247) );
  MUX21L U18850 ( .A(n4586), .B(n3175), .S(n5232), .Z(n1287) );
  ND2 U18851 ( .A(n4586), .B(n4833), .Z(n3175) );
  AO7 U18852 ( .A(n5247), .B(n4418), .C(n3535), .Z(n1292) );
  ND2 U18853 ( .A(n4923), .B(n4573), .Z(n3535) );
  MUX21L U18854 ( .A(n3270), .B(n4484), .S(n4951), .Z(n1288) );
  ND2 U18855 ( .A(n5253), .B(n4484), .Z(n3270) );
  MUX21L U18856 ( .A(n3570), .B(n3569), .S(n4925), .Z(n1293) );
  ND2 U18857 ( .A(n4414), .B(n5128), .Z(n3570) );
  ND2 U18858 ( .A(n4575), .B(n5128), .Z(n3569) );
  AN3 U18859 ( .A(n4548), .B(n5182), .C(n4947), .Z(n772) );
  MUX21L U18860 ( .A(n4838), .B(n5251), .S(n4614), .Z(n1817) );
  ND2 U18861 ( .A(n2295), .B(n2294), .Z(n1271) );
  ND2 U18862 ( .A(n4630), .B(n4962), .Z(n2294) );
  MUX21L U18863 ( .A(n2293), .B(n5152), .S(n4962), .Z(n2295) );
  NR2 U18864 ( .A(n4630), .B(n5151), .Z(n2293) );
  ND2 U18865 ( .A(n3322), .B(n3321), .Z(n1289) );
  ND2 U18866 ( .A(n4608), .B(n4768), .Z(n3321) );
  MUX21L U18867 ( .A(n3320), .B(n5255), .S(n4608), .Z(n3322) );
  NR2 U18868 ( .A(n5256), .B(n4896), .Z(n3320) );
  IVP U18869 ( .A(n4729), .Z(n4928) );
  ND2 U18870 ( .A(n3130), .B(n3129), .Z(n1781) );
  MUX21L U18871 ( .A(n3127), .B(n5092), .S(n4583), .Z(n3129) );
  AO6 U18872 ( .A(n4583), .B(n4826), .C(n3128), .Z(n3130) );
  AO7 U18873 ( .A(n4584), .B(n5090), .C(n4958), .Z(n1286) );
  NR2 U18874 ( .A(n5274), .B(n4765), .Z(n2159) );
  NR2 U18875 ( .A(n5274), .B(n4461), .Z(n2160) );
  NR2 U18876 ( .A(n4906), .B(n5201), .Z(n2732) );
  ND2 U18877 ( .A(n3328), .B(n5071), .Z(n1784) );
  EO U18878 ( .A(n4897), .B(n4607), .Z(n3328) );
  ND2 U18879 ( .A(n2836), .B(n5191), .Z(n1774) );
  EN U18880 ( .A(n4900), .B(n4564), .Z(n2836) );
  ND2 U18881 ( .A(n2577), .B(n2576), .Z(n1767) );
  ND2 U18882 ( .A(n4621), .B(n5215), .Z(n2576) );
  EO U18883 ( .A(n5226), .B(n4974), .Z(n2577) );
  ND3 U18884 ( .A(n3041), .B(n3040), .C(n3039), .Z(n1778) );
  ND2 U18885 ( .A(n4384), .B(n4816), .Z(n3040) );
  ND2 U18886 ( .A(n5239), .B(n4816), .Z(n3041) );
  ND2 U18887 ( .A(n5239), .B(n4385), .Z(n3039) );
  ND3 U18888 ( .A(n4826), .B(n5092), .C(n4376), .Z(n1316) );
  ND2 U18889 ( .A(n2642), .B(n2641), .Z(n1769) );
  ND2 U18890 ( .A(n5292), .B(n4896), .Z(n2642) );
  ND2 U18891 ( .A(n4624), .B(n4895), .Z(n2641) );
  ND2 U18892 ( .A(n5291), .B(n4516), .Z(n1803) );
  ND2 U18893 ( .A(n4564), .B(n4737), .Z(n1280) );
  MUX21L U18894 ( .A(n2158), .B(n4598), .S(n4914), .Z(n2161) );
  NR2 U18895 ( .A(n4598), .B(n5163), .Z(n2158) );
  ND2 U18896 ( .A(n2760), .B(n2759), .Z(n1773) );
  ND2 U18897 ( .A(n4928), .B(n4498), .Z(n2759) );
  MUX21L U18898 ( .A(n5197), .B(n2758), .S(n4560), .Z(n2760) );
  NR2 U18899 ( .A(n4928), .B(n5197), .Z(n2758) );
  ND2 U18900 ( .A(n2734), .B(n2733), .Z(n1772) );
  ND2 U18901 ( .A(n2730), .B(n4752), .Z(n2733) );
  MUX21L U18902 ( .A(n2731), .B(n2732), .S(n4558), .Z(n2734) );
  NR2 U18903 ( .A(n5277), .B(n4558), .Z(n2730) );
  ND2 U18904 ( .A(n2439), .B(n2438), .Z(n1765) );
  ND2 U18905 ( .A(n4616), .B(n4764), .Z(n2438) );
  MUX21L U18906 ( .A(n5266), .B(n2437), .S(n4915), .Z(n2439) );
  NR2 U18907 ( .A(n5266), .B(n4616), .Z(n2437) );
  MUX21L U18908 ( .A(n2569), .B(n2570), .S(n5289), .Z(n2572) );
  NR2 U18909 ( .A(n4974), .B(n4523), .Z(n2569) );
  ND2 U18910 ( .A(n2881), .B(n2880), .Z(n1253) );
  ND2 U18911 ( .A(n2877), .B(n5189), .Z(n2880) );
  MUX21L U18912 ( .A(n2878), .B(n2879), .S(n4566), .Z(n2881) );
  NR2 U18913 ( .A(n4566), .B(n4933), .Z(n2877) );
  ND2 U18914 ( .A(n2378), .B(n2377), .Z(n1246) );
  ND2 U18915 ( .A(n4880), .B(n5143), .Z(n2377) );
  MUX21L U18916 ( .A(n5143), .B(n2376), .S(n4635), .Z(n2378) );
  IVP U18917 ( .A(n4725), .Z(n4953) );
  IVP U18918 ( .A(n5066), .Z(n5249) );
  AO7 U18919 ( .A(n5238), .B(n4825), .C(n4378), .Z(n1779) );
  ND2 U18920 ( .A(n2182), .B(n2181), .Z(n1241) );
  MUX21L U18921 ( .A(n2179), .B(n5161), .S(n4967), .Z(n2181) );
  AO6 U18922 ( .A(n4967), .B(n4463), .C(n2180), .Z(n2182) );
  NR2 U18923 ( .A(n5284), .B(n4801), .Z(n2879) );
  ND2 U18924 ( .A(n4614), .B(n5081), .Z(n3221) );
  ND2 U18925 ( .A(n2594), .B(n2593), .Z(n1768) );
  ND2 U18926 ( .A(n4519), .B(n5214), .Z(n2594) );
  ND2 U18927 ( .A(n4973), .B(n4519), .Z(n2593) );
  ND2 U18928 ( .A(n4625), .B(n5208), .Z(n2653) );
  ND2 U18929 ( .A(n2509), .B(n2508), .Z(n1248) );
  ND2 U18930 ( .A(n4591), .B(n4758), .Z(n2508) );
  MUX21L U18931 ( .A(n2507), .B(n5287), .S(n4592), .Z(n2509) );
  NR2 U18932 ( .A(n5287), .B(n4758), .Z(n2507) );
  ND2 U18933 ( .A(n2100), .B(n2099), .Z(n1239) );
  ND2 U18934 ( .A(n4911), .B(n5169), .Z(n2099) );
  MUX21L U18935 ( .A(n2098), .B(n4455), .S(n4911), .Z(n2100) );
  ND2 U18936 ( .A(n2152), .B(n2151), .Z(n1240) );
  ND2 U18937 ( .A(n4766), .B(n5165), .Z(n2151) );
  MUX21L U18938 ( .A(n4766), .B(n2150), .S(n4599), .Z(n2152) );
  ND2 U18939 ( .A(n2289), .B(n2288), .Z(n1243) );
  ND2 U18940 ( .A(n4962), .B(n4540), .Z(n2288) );
  EO U18941 ( .A(n5222), .B(n4630), .Z(n2289) );
  MUX21L U18942 ( .A(n3177), .B(n3176), .S(n4955), .Z(n1259) );
  ND2 U18943 ( .A(n4436), .B(n5087), .Z(n3177) );
  ND2 U18944 ( .A(n4586), .B(n5087), .Z(n3176) );
  AN3 U18945 ( .A(n4429), .B(n5111), .C(n4918), .Z(n773) );
  MUX21L U18946 ( .A(n2395), .B(n2394), .S(n4977), .Z(n1764) );
  ND2 U18947 ( .A(n4636), .B(n5140), .Z(n2394) );
  ND2 U18948 ( .A(n5265), .B(n4636), .Z(n2395) );
  MUX21L U18949 ( .A(n2318), .B(n4538), .S(n5261), .Z(n2320) );
  ND2 U18950 ( .A(n2089), .B(n2088), .Z(n1728) );
  ND2 U18951 ( .A(n4454), .B(n4853), .Z(n2088) );
  EN U18952 ( .A(n5228), .B(n4602), .Z(n2089) );
  AO7 U18953 ( .A(n5295), .B(n4754), .C(n4505), .Z(n1770) );
  NR2 U18954 ( .A(n4595), .B(n5160), .Z(n2220) );
  ND2 U18955 ( .A(n4591), .B(n4757), .Z(n1766) );
  ND2 U18956 ( .A(n4600), .B(n4751), .Z(n2136) );
  ND2 U18957 ( .A(n5270), .B(n4447), .Z(n2045) );
  ND2 U18958 ( .A(n2972), .B(n5180), .Z(n1744) );
  EO U18959 ( .A(n4899), .B(n4550), .Z(n2972) );
  ND2 U18960 ( .A(n2816), .B(n2815), .Z(n1743) );
  ND2 U18961 ( .A(n5280), .B(n4407), .Z(n2815) );
  EN U18962 ( .A(n5222), .B(n4930), .Z(n2816) );
  ND2 U18963 ( .A(n5261), .B(n4875), .Z(n2319) );
  ND2 U18964 ( .A(n4594), .B(n4867), .Z(n2248) );
  ND2 U18965 ( .A(n3509), .B(n3508), .Z(n1263) );
  ND2 U18966 ( .A(n4422), .B(n5120), .Z(n3509) );
  ND2 U18967 ( .A(n4921), .B(n4422), .Z(n3508) );
  ND2 U18968 ( .A(n2239), .B(n2238), .Z(n1731) );
  ND2 U18969 ( .A(n4965), .B(n4469), .Z(n2238) );
  MUX21L U18970 ( .A(n2237), .B(n4470), .S(n5276), .Z(n2239) );
  NR2 U18971 ( .A(n4965), .B(n4469), .Z(n2237) );
  ND2 U18972 ( .A(n3196), .B(n3195), .Z(n1750) );
  MUX21L U18973 ( .A(n3193), .B(n3194), .S(n4954), .Z(n3195) );
  MUX21L U18974 ( .A(n3191), .B(n3192), .S(n5231), .Z(n3196) );
  NR2 U18975 ( .A(n4587), .B(n5085), .Z(n3193) );
  ND2 U18976 ( .A(n3406), .B(n3405), .Z(n1754) );
  ND2 U18977 ( .A(n4937), .B(n5110), .Z(n3405) );
  MUX21L U18978 ( .A(n3404), .B(n4431), .S(n4937), .Z(n3406) );
  ND2 U18979 ( .A(n2797), .B(n2796), .Z(n1224) );
  ND2 U18980 ( .A(n4929), .B(n4494), .Z(n2796) );
  EO U18981 ( .A(n5222), .B(n4561), .Z(n2797) );
  IVP U18982 ( .A(n4370), .Z(n4563) );
  AO7 U18983 ( .A(n4572), .B(n4776), .C(n5122), .Z(n1755) );
  AO7 U18984 ( .A(n5289), .B(n4888), .C(n2578), .Z(n1736) );
  ND2 U18985 ( .A(n4974), .B(n4621), .Z(n2578) );
  AO7 U18986 ( .A(n4625), .B(n5206), .C(n4803), .Z(n1738) );
  NR2 U18987 ( .A(n4954), .B(n4434), .Z(n3191) );
  ND2 U18988 ( .A(n4478), .B(n5081), .Z(n3222) );
  ND2 U18989 ( .A(n4566), .B(n4801), .Z(n2882) );
  ND2 U18990 ( .A(n4566), .B(n5188), .Z(n2884) );
  ND2 U18991 ( .A(n3553), .B(n3552), .Z(n1756) );
  ND2 U18992 ( .A(n4775), .B(n5126), .Z(n3553) );
  ND2 U18993 ( .A(n4574), .B(n4775), .Z(n3552) );
  ND2 U18994 ( .A(n2618), .B(n2617), .Z(n1737) );
  ND2 U18995 ( .A(n4623), .B(n5291), .Z(n2617) );
  MUX21L U18996 ( .A(n2616), .B(n4972), .S(n5291), .Z(n2618) );
  NR2 U18997 ( .A(n4972), .B(n4623), .Z(n2616) );
  ND2 U18998 ( .A(n2441), .B(n2440), .Z(n1735) );
  ND2 U18999 ( .A(n4528), .B(n4764), .Z(n2440) );
  EN U19000 ( .A(n5224), .B(n4616), .Z(n2441) );
  ND2 U19001 ( .A(n4942), .B(n4384), .Z(n3046) );
  ND2 U19002 ( .A(n2545), .B(n2544), .Z(n1220) );
  ND2 U19003 ( .A(n2541), .B(n5217), .Z(n2544) );
  MUX21L U19004 ( .A(n2542), .B(n2543), .S(n4619), .Z(n2545) );
  NR2 U19005 ( .A(n4619), .B(n4975), .Z(n2541) );
  ND2 U19006 ( .A(n2604), .B(n2603), .Z(n1221) );
  ND2 U19007 ( .A(n4972), .B(n4519), .Z(n2603) );
  MUX21L U19008 ( .A(n5212), .B(n2602), .S(n4622), .Z(n2604) );
  NR2 U19009 ( .A(n4972), .B(n5212), .Z(n2602) );
  ND2 U19010 ( .A(n2282), .B(n2281), .Z(n1214) );
  ND2 U19011 ( .A(n5260), .B(n4871), .Z(n2281) );
  MUX21L U19012 ( .A(n4872), .B(n2280), .S(n4629), .Z(n2282) );
  NR2 U19013 ( .A(n5260), .B(n4871), .Z(n2280) );
  ND2 U19014 ( .A(n3453), .B(n3452), .Z(n1234) );
  ND2 U19015 ( .A(n4783), .B(n5114), .Z(n3452) );
  MUX21L U19016 ( .A(n5114), .B(n3451), .S(n4591), .Z(n3453) );
  ND2 U19017 ( .A(n3530), .B(n3529), .Z(n1235) );
  ND2 U19018 ( .A(n4419), .B(n5123), .Z(n3529) );
  EO U19019 ( .A(n5229), .B(n4923), .Z(n3530) );
  MUX21L U19020 ( .A(n5080), .B(n3223), .S(n4613), .Z(n1751) );
  ND2 U19021 ( .A(n4953), .B(n5081), .Z(n3223) );
  MUX21L U19022 ( .A(n4604), .B(n4790), .S(n5258), .Z(n1753) );
  MUX21L U19023 ( .A(n4486), .B(n4950), .S(n5254), .Z(n1752) );
  MUX21L U19024 ( .A(n2693), .B(n5294), .S(n4556), .Z(n1739) );
  ND2 U19025 ( .A(n5294), .B(n4906), .Z(n2693) );
  MUX21L U19026 ( .A(n5100), .B(n3045), .S(n4555), .Z(n3047) );
  NR2 U19027 ( .A(n4942), .B(n5100), .Z(n3045) );
  ND2 U19028 ( .A(n3355), .B(n3354), .Z(n1233) );
  ND3 U19029 ( .A(n4935), .B(n4491), .C(n5257), .Z(n3354) );
  MUX21L U19030 ( .A(n3352), .B(n3353), .S(n4935), .Z(n3355) );
  NR2 U19031 ( .A(n5257), .B(n4491), .Z(n3353) );
  NR2 U19032 ( .A(n5288), .B(n4885), .Z(n2543) );
  NR2 U19033 ( .A(n4904), .B(n4477), .Z(n2511) );
  ND2 U19034 ( .A(n4448), .B(n5173), .Z(n2056) );
  ND2 U19035 ( .A(n4960), .B(n4537), .Z(n2321) );
  ND2 U19036 ( .A(n4599), .B(n5166), .Z(n2145) );
  ND2 U19037 ( .A(n4599), .B(n4767), .Z(n2146) );
  ND2 U19038 ( .A(n2059), .B(n2058), .Z(n1209) );
  ND2 U19039 ( .A(n4909), .B(n4449), .Z(n2058) );
  MUX21L U19040 ( .A(n2057), .B(n4449), .S(n5270), .Z(n2059) );
  NR2 U19041 ( .A(n4909), .B(n4449), .Z(n2057) );
  AN3 U19042 ( .A(n4481), .B(n5078), .C(n4952), .Z(n774) );
  ND2 U19043 ( .A(n3557), .B(n3556), .Z(n1725) );
  AO6 U19044 ( .A(n4574), .B(n4774), .C(n3555), .Z(n3557) );
  MUX21L U19045 ( .A(n3554), .B(n5126), .S(n4574), .Z(n3556) );
  NR2 U19046 ( .A(n5248), .B(n4924), .Z(n3555) );
  MUX21L U19047 ( .A(n4853), .B(n2101), .S(n4602), .Z(n1210) );
  ND2 U19048 ( .A(n4853), .B(n5168), .Z(n2101) );
  MUX21L U19049 ( .A(n3149), .B(n3148), .S(n5236), .Z(n1230) );
  ND2 U19050 ( .A(n4443), .B(n4829), .Z(n3149) );
  ND2 U19051 ( .A(n4958), .B(n4442), .Z(n3148) );
  MUX21L U19052 ( .A(n5073), .B(n3302), .S(n4609), .Z(n1232) );
  ND2 U19053 ( .A(n4949), .B(n5073), .Z(n3302) );
  AO7 U19054 ( .A(n4970), .B(n4625), .C(n5207), .Z(n1708) );
  ND2 U19055 ( .A(n2200), .B(n2199), .Z(n1699) );
  ND2 U19056 ( .A(n4966), .B(n4465), .Z(n2199) );
  EO U19057 ( .A(n5230), .B(n4596), .Z(n2200) );
  ND2 U19058 ( .A(n4610), .B(n5075), .Z(n3287) );
  ND2 U19059 ( .A(n4965), .B(n5158), .Z(n2240) );
  ND2 U19060 ( .A(n3390), .B(n3389), .Z(n1722) );
  ND2 U19061 ( .A(n4603), .B(n4937), .Z(n3389) );
  MUX21L U19062 ( .A(n3388), .B(n5109), .S(n4937), .Z(n3390) );
  NR2 U19063 ( .A(n4603), .B(n5109), .Z(n3388) );
  MUX21L U19064 ( .A(n4890), .B(n2595), .S(n5290), .Z(n1707) );
  ND2 U19065 ( .A(n4622), .B(n4890), .Z(n2595) );
  ND2 U19066 ( .A(n4490), .B(n4797), .Z(n1261) );
  ND2 U19067 ( .A(n5292), .B(n4873), .Z(n2655) );
  ND2 U19068 ( .A(n5292), .B(n4514), .Z(n2656) );
  AN3 U19069 ( .A(n4504), .B(n5201), .C(n4906), .Z(n775) );
  ND2 U19070 ( .A(n2139), .B(n2138), .Z(n1698) );
  ND2 U19071 ( .A(n4913), .B(n4459), .Z(n2138) );
  MUX21L U19072 ( .A(n5167), .B(n2137), .S(n4600), .Z(n2139) );
  NR2 U19073 ( .A(n4913), .B(n5166), .Z(n2137) );
  MUX21L U19074 ( .A(n3083), .B(n5237), .S(n4580), .Z(n1717) );
  ND2 U19075 ( .A(n5237), .B(n4822), .Z(n3083) );
  MUX21L U19076 ( .A(n4736), .B(n4403), .S(n5282), .Z(n1712) );
  MUX21L U19077 ( .A(n4555), .B(n4819), .S(n5231), .Z(n1716) );
  ND2 U19078 ( .A(n2357), .B(n2356), .Z(n1703) );
  ND2 U19079 ( .A(n5262), .B(n4534), .Z(n2356) );
  MUX21L U19080 ( .A(n4879), .B(n2355), .S(n4634), .Z(n2357) );
  NR2 U19081 ( .A(n5263), .B(n4878), .Z(n2355) );
  MUX21L U19082 ( .A(n2695), .B(n2694), .S(n4907), .Z(n1709) );
  ND2 U19083 ( .A(n5294), .B(n4556), .Z(n2695) );
  ND2 U19084 ( .A(n4556), .B(n5204), .Z(n2694) );
  ND2 U19085 ( .A(n2444), .B(n2443), .Z(n1705) );
  ND2 U19086 ( .A(n5266), .B(n4763), .Z(n2443) );
  MUX21L U19087 ( .A(n4764), .B(n2442), .S(n4616), .Z(n2444) );
  NR2 U19088 ( .A(n5266), .B(n4763), .Z(n2442) );
  NR2 U19089 ( .A(n4941), .B(n4383), .Z(n3060) );
  NR2 U19090 ( .A(n4942), .B(n5098), .Z(n3059) );
  NR2 U19091 ( .A(n4931), .B(n4403), .Z(n2843) );
  ND2 U19092 ( .A(n3062), .B(n3061), .Z(n1199) );
  MUX21L U19093 ( .A(n3058), .B(n4556), .S(n5231), .Z(n3061) );
  NR2 U19094 ( .A(n3060), .B(n3059), .Z(n3062) );
  NR2 U19095 ( .A(n4556), .B(n4819), .Z(n3058) );
  ND2 U19096 ( .A(n2362), .B(n2361), .Z(n1187) );
  ND2 U19097 ( .A(n4634), .B(n5145), .Z(n2361) );
  EN U19098 ( .A(n4897), .B(n4634), .Z(n2362) );
  ND3 U19099 ( .A(n2909), .B(n2908), .C(n2907), .Z(n1197) );
  ND2 U19100 ( .A(n4934), .B(n5186), .Z(n2909) );
  ND2 U19101 ( .A(n4567), .B(n5186), .Z(n2908) );
  ND2 U19102 ( .A(n4934), .B(n4567), .Z(n2907) );
  ND2 U19103 ( .A(n4944), .B(n5177), .Z(n1715) );
  ND2 U19104 ( .A(n4867), .B(n5157), .Z(n2249) );
  ND2 U19105 ( .A(n4593), .B(n4760), .Z(n2491) );
  ND2 U19106 ( .A(n4593), .B(n5134), .Z(n2493) );
  ND2 U19107 ( .A(n3357), .B(n3356), .Z(n1204) );
  ND2 U19108 ( .A(n5257), .B(n4492), .Z(n3356) );
  EN U19109 ( .A(n4897), .B(n4605), .Z(n3357) );
  MUX21L U19110 ( .A(n3324), .B(n3323), .S(n5256), .Z(n1203) );
  ND2 U19111 ( .A(n4948), .B(n4489), .Z(n3324) );
  ND2 U19112 ( .A(n4948), .B(n4608), .Z(n3323) );
  ND2 U19113 ( .A(n2582), .B(n2581), .Z(n1191) );
  ND2 U19114 ( .A(n4522), .B(n5214), .Z(n2581) );
  EO U19115 ( .A(n4903), .B(n4621), .Z(n2582) );
  ND2 U19116 ( .A(n2684), .B(n2683), .Z(n1193) );
  ND2 U19117 ( .A(n5293), .B(n4620), .Z(n2683) );
  EN U19118 ( .A(n5225), .B(n4905), .Z(n2684) );
  MUX21L U19119 ( .A(n4746), .B(n2776), .S(n5279), .Z(n1195) );
  ND2 U19120 ( .A(n4560), .B(n4746), .Z(n2776) );
  ND2 U19121 ( .A(n5262), .B(n4959), .Z(n2354) );
  AN3 U19122 ( .A(n4481), .B(n4839), .C(n5252), .Z(n776) );
  ND2 U19123 ( .A(n3281), .B(n4485), .Z(n1691) );
  EN U19124 ( .A(n5225), .B(n4950), .Z(n3281) );
  IVP U19125 ( .A(n4371), .Z(n4570) );
  NR2 U19126 ( .A(n4915), .B(n5138), .Z(n2447) );
  NR2 U19127 ( .A(n4972), .B(n5211), .Z(n2620) );
  NR2 U19128 ( .A(n4972), .B(n4518), .Z(n2621) );
  ND2 U19129 ( .A(n4416), .B(n5126), .Z(n3559) );
  ND2 U19130 ( .A(n4924), .B(n5127), .Z(n3558) );
  ND2 U19131 ( .A(n4570), .B(n4781), .Z(n3485) );
  ND2 U19132 ( .A(n4570), .B(n5118), .Z(n3487) );
  ND2 U19133 ( .A(n2764), .B(n2763), .Z(n1683) );
  MUX21L U19134 ( .A(n2761), .B(n5196), .S(n4928), .Z(n2763) );
  AO6 U19135 ( .A(n4928), .B(n4497), .C(n2762), .Z(n2764) );
  ND2 U19136 ( .A(n2915), .B(n4397), .Z(n1685) );
  EO U19137 ( .A(n5228), .B(n4969), .Z(n2915) );
  MUX21L U19138 ( .A(n2818), .B(n2817), .S(n4563), .Z(n1684) );
  ND2 U19139 ( .A(n5280), .B(n4930), .Z(n2818) );
  ND2 U19140 ( .A(n4930), .B(n5192), .Z(n2817) );
  MUX21L U19141 ( .A(n4873), .B(n2312), .S(n5260), .Z(n1673) );
  ND2 U19142 ( .A(n4631), .B(n4874), .Z(n2312) );
  ND2 U19143 ( .A(n2531), .B(n2530), .Z(n1678) );
  ND2 U19144 ( .A(n4618), .B(n5218), .Z(n2530) );
  MUX21L U19145 ( .A(n2529), .B(n5218), .S(n4975), .Z(n2531) );
  NR2 U19146 ( .A(n4619), .B(n5218), .Z(n2529) );
  ND2 U19147 ( .A(n2623), .B(n2622), .Z(n1679) );
  MUX21L U19148 ( .A(n2619), .B(n4623), .S(n5291), .Z(n2622) );
  NR2 U19149 ( .A(n2621), .B(n2620), .Z(n2623) );
  NR2 U19150 ( .A(n4623), .B(n4892), .Z(n2619) );
  AN3 U19151 ( .A(n4580), .B(n5095), .C(n4941), .Z(n777) );
  MUX21L U19152 ( .A(n4430), .B(n5242), .S(n4933), .Z(n1694) );
  ND2 U19153 ( .A(n3009), .B(n3008), .Z(n1687) );
  ND2 U19154 ( .A(n4812), .B(n5102), .Z(n3008) );
  MUX21L U19155 ( .A(n4813), .B(n3007), .S(n4552), .Z(n3009) );
  ND2 U19156 ( .A(n2260), .B(n2259), .Z(n1671) );
  ND2 U19157 ( .A(n4593), .B(n4964), .Z(n2259) );
  MUX21L U19158 ( .A(n2258), .B(n5155), .S(n4964), .Z(n2260) );
  NR2 U19159 ( .A(n4593), .B(n5154), .Z(n2258) );
  ND2 U19160 ( .A(n2203), .B(n2202), .Z(n1670) );
  ND2 U19161 ( .A(n5275), .B(n4966), .Z(n2202) );
  MUX21L U19162 ( .A(n2201), .B(n4465), .S(n4966), .Z(n2203) );
  NR2 U19163 ( .A(n5275), .B(n4465), .Z(n2201) );
  ND2 U19164 ( .A(n2050), .B(n2049), .Z(n1667) );
  ND2 U19165 ( .A(n4909), .B(n4447), .Z(n2049) );
  MUX21L U19166 ( .A(n2048), .B(n4448), .S(n5270), .Z(n2050) );
  NR2 U19167 ( .A(n4909), .B(n4447), .Z(n2048) );
  ND2 U19168 ( .A(n2449), .B(n2448), .Z(n1677) );
  ND2 U19169 ( .A(n2445), .B(n4763), .Z(n2448) );
  MUX21L U19170 ( .A(n2446), .B(n2447), .S(n4616), .Z(n2449) );
  NR2 U19171 ( .A(n5266), .B(n4616), .Z(n2445) );
  NR2 U19172 ( .A(n4941), .B(n4383), .Z(n3064) );
  ND2 U19173 ( .A(n2381), .B(n2380), .Z(n1675) );
  ND2 U19174 ( .A(n4635), .B(n5142), .Z(n2380) );
  EO U19175 ( .A(n5223), .B(n4978), .Z(n2381) );
  ND3 U19176 ( .A(n4907), .B(n4557), .C(n5294), .Z(n1680) );
  ND2 U19177 ( .A(n4563), .B(n4738), .Z(n2832) );
  ND2 U19178 ( .A(n4563), .B(n5192), .Z(n2834) );
  ND2 U19179 ( .A(n3000), .B(n2999), .Z(n1170) );
  ND2 U19180 ( .A(n4945), .B(n5178), .Z(n2999) );
  MUX21L U19181 ( .A(n2998), .B(n4389), .S(n4945), .Z(n3000) );
  ND2 U19182 ( .A(n3113), .B(n3112), .Z(n1172) );
  ND2 U19183 ( .A(n4825), .B(n5093), .Z(n3112) );
  MUX21L U19184 ( .A(n5094), .B(n3111), .S(n4582), .Z(n3113) );
  ND2 U19185 ( .A(n3511), .B(n3510), .Z(n1179) );
  ND2 U19186 ( .A(n5246), .B(n4779), .Z(n3511) );
  ND2 U19187 ( .A(n4571), .B(n4778), .Z(n3510) );
  ND2 U19188 ( .A(n2659), .B(n2658), .Z(n1165) );
  ND2 U19189 ( .A(n4970), .B(n4513), .Z(n2658) );
  MUX21L U19190 ( .A(n2657), .B(n4514), .S(n5292), .Z(n2659) );
  NR2 U19191 ( .A(n4970), .B(n4513), .Z(n2657) );
  ND2 U19192 ( .A(n2398), .B(n2397), .Z(n1676) );
  ND2 U19193 ( .A(n4977), .B(n4530), .Z(n2397) );
  MUX21L U19194 ( .A(n5140), .B(n2396), .S(n4636), .Z(n2398) );
  NR2 U19195 ( .A(n4977), .B(n5140), .Z(n2396) );
  MUX21L U19196 ( .A(n3420), .B(n3419), .S(n4589), .Z(n1178) );
  ND2 U19197 ( .A(n4787), .B(n5112), .Z(n3419) );
  ND2 U19198 ( .A(n4918), .B(n5111), .Z(n3420) );
  MUX21L U19199 ( .A(n3150), .B(n5236), .S(n4584), .Z(n1174) );
  ND2 U19200 ( .A(n5236), .B(n4830), .Z(n3150) );
  ND2 U19201 ( .A(n2171), .B(n2170), .Z(n1638) );
  ND2 U19202 ( .A(n4598), .B(n5163), .Z(n2170) );
  EN U19203 ( .A(n4903), .B(n4598), .Z(n2171) );
  NR2 U19204 ( .A(n4548), .B(n4804), .Z(n2931) );
  NR2 U19205 ( .A(n4929), .B(n5194), .Z(n2789) );
  NR2 U19206 ( .A(n4929), .B(n4495), .Z(n2790) );
  ND2 U19207 ( .A(n2242), .B(n2241), .Z(n1639) );
  ND2 U19208 ( .A(n5276), .B(n4470), .Z(n2241) );
  EN U19209 ( .A(n4902), .B(n4595), .Z(n2242) );
  ND2 U19210 ( .A(n4398), .B(n5185), .Z(n1713) );
  ND2 U19211 ( .A(n2792), .B(n2791), .Z(n1650) );
  MUX21L U19212 ( .A(n2788), .B(n4561), .S(n5279), .Z(n2791) );
  NR2 U19213 ( .A(n2790), .B(n2789), .Z(n2792) );
  NR2 U19214 ( .A(n4561), .B(n4743), .Z(n2788) );
  ND2 U19215 ( .A(n3106), .B(n3105), .Z(n1656) );
  ND2 U19216 ( .A(n4581), .B(n4824), .Z(n3105) );
  MUX21L U19217 ( .A(n3104), .B(n5241), .S(n4581), .Z(n3106) );
  NR2 U19218 ( .A(n5240), .B(n4824), .Z(n3104) );
  ND2 U19219 ( .A(n2737), .B(n2736), .Z(n1649) );
  ND2 U19220 ( .A(n4559), .B(n5200), .Z(n2736) );
  MUX21L U19221 ( .A(n2735), .B(n5201), .S(n4906), .Z(n2737) );
  NR2 U19222 ( .A(n4559), .B(n5200), .Z(n2735) );
  ND2 U19223 ( .A(n3460), .B(n3459), .Z(n1663) );
  ND2 U19224 ( .A(n4568), .B(n5115), .Z(n3459) );
  EO U19225 ( .A(n4899), .B(n4568), .Z(n3460) );
  ND2 U19226 ( .A(n2628), .B(n2627), .Z(n1645) );
  ND2 U19227 ( .A(n2624), .B(n5291), .Z(n2627) );
  MUX21L U19228 ( .A(n2625), .B(n2626), .S(n5291), .Z(n2628) );
  NR2 U19229 ( .A(n4972), .B(n4623), .Z(n2624) );
  ND2 U19230 ( .A(n4891), .B(n5211), .Z(n2605) );
  ND2 U19231 ( .A(n4759), .B(n5134), .Z(n2492) );
  ND2 U19232 ( .A(n2479), .B(n4473), .Z(n1163) );
  ND2 U19233 ( .A(n5268), .B(n4916), .Z(n2479) );
  MUX21L U19234 ( .A(n2274), .B(n4541), .S(n5259), .Z(n2276) );
  NR2 U19235 ( .A(n4963), .B(n4541), .Z(n2274) );
  AO7 U19236 ( .A(n5233), .B(n4832), .C(n4585), .Z(n1659) );
  AO7 U19237 ( .A(n4935), .B(n4490), .C(n5256), .Z(n1662) );
  AO7 U19238 ( .A(n5289), .B(n4621), .C(n4888), .Z(n1644) );
  NR2 U19239 ( .A(n5285), .B(n4396), .Z(n2929) );
  NR2 U19240 ( .A(n4972), .B(n4517), .Z(n2625) );
  NR2 U19241 ( .A(n4938), .B(n5092), .Z(n1658) );
  ND2 U19242 ( .A(n5232), .B(n4382), .Z(n3069) );
  ND2 U19243 ( .A(n4941), .B(n5232), .Z(n3070) );
  ND2 U19244 ( .A(n4941), .B(n4382), .Z(n3068) );
  ND2 U19245 ( .A(n4563), .B(n5192), .Z(n2819) );
  ND2 U19246 ( .A(n4563), .B(n4739), .Z(n2820) );
  ND2 U19247 ( .A(n5233), .B(n4810), .Z(n2990) );
  ND2 U19248 ( .A(n5295), .B(n2712), .Z(n1647) );
  ND2 U19249 ( .A(n4908), .B(n4557), .Z(n2712) );
  ND2 U19250 ( .A(n3153), .B(n3152), .Z(n1150) );
  ND2 U19251 ( .A(n4584), .B(n4830), .Z(n3152) );
  MUX21L U19252 ( .A(n5235), .B(n3151), .S(n4957), .Z(n3153) );
  NR2 U19253 ( .A(n5235), .B(n4584), .Z(n3151) );
  MUX21L U19254 ( .A(n4487), .B(n5254), .S(n4950), .Z(n1661) );
  MUX21L U19255 ( .A(n2451), .B(n2450), .S(n4616), .Z(n1643) );
  ND2 U19256 ( .A(n4762), .B(n5138), .Z(n2450) );
  ND2 U19257 ( .A(n5267), .B(n4915), .Z(n2451) );
  ND2 U19258 ( .A(n2768), .B(n2767), .Z(n1618) );
  MUX21L U19259 ( .A(n2765), .B(n5196), .S(n4928), .Z(n2767) );
  AO6 U19260 ( .A(n4928), .B(n4497), .C(n2766), .Z(n2768) );
  ND2 U19261 ( .A(n3228), .B(n3227), .Z(n1628) );
  ND2 U19262 ( .A(n3224), .B(n4839), .Z(n3227) );
  MUX21L U19263 ( .A(n3225), .B(n3226), .S(n4613), .Z(n3228) );
  NR2 U19264 ( .A(n5251), .B(n4613), .Z(n3224) );
  ND2 U19265 ( .A(n4737), .B(n5191), .Z(n2833) );
  ND2 U19266 ( .A(n4745), .B(n5195), .Z(n2777) );
  ND2 U19267 ( .A(n4607), .B(n4797), .Z(n1152) );
  NR2 U19268 ( .A(n4953), .B(n5080), .Z(n3226) );
  ND3 U19269 ( .A(n2963), .B(n2962), .C(n2961), .Z(n1621) );
  ND2 U19270 ( .A(n5282), .B(n4808), .Z(n2962) );
  ND2 U19271 ( .A(n4548), .B(n5286), .Z(n2963) );
  ND2 U19272 ( .A(n4550), .B(n4808), .Z(n2961) );
  ND3 U19273 ( .A(n2598), .B(n2597), .C(n2596), .Z(n1614) );
  ND2 U19274 ( .A(n4890), .B(n5213), .Z(n2597) );
  ND2 U19275 ( .A(n4622), .B(n5213), .Z(n2598) );
  ND2 U19276 ( .A(n4622), .B(n4891), .Z(n2596) );
  ND2 U19277 ( .A(n4391), .B(n4810), .Z(n2991) );
  ND2 U19278 ( .A(n5281), .B(n4739), .Z(n2821) );
  ND2 U19279 ( .A(n5281), .B(n4406), .Z(n2822) );
  ND2 U19280 ( .A(n5283), .B(n4735), .Z(n2866) );
  ND2 U19281 ( .A(n4559), .B(n4752), .Z(n2738) );
  ND2 U19282 ( .A(n5278), .B(n4752), .Z(n2739) );
  ND2 U19283 ( .A(n3339), .B(n3338), .Z(n1630) );
  ND2 U19284 ( .A(n4606), .B(n5103), .Z(n3338) );
  MUX21L U19285 ( .A(n4795), .B(n3337), .S(n5257), .Z(n3339) );
  NR2 U19286 ( .A(n4606), .B(n4795), .Z(n3337) );
  ND2 U19287 ( .A(n2681), .B(n2680), .Z(n1615) );
  ND2 U19288 ( .A(n4626), .B(n4904), .Z(n2680) );
  MUX21L U19289 ( .A(n2679), .B(n5206), .S(n4904), .Z(n2681) );
  NR2 U19290 ( .A(n4626), .B(n5205), .Z(n2679) );
  ND2 U19291 ( .A(n2478), .B(n4473), .Z(n1611) );
  ND2 U19292 ( .A(n5268), .B(n4916), .Z(n2478) );
  ND2 U19293 ( .A(n4531), .B(n4882), .Z(n1161) );
  ND2 U19294 ( .A(n4516), .B(n4894), .Z(n1164) );
  MUX21L U19295 ( .A(n3132), .B(n3131), .S(n4583), .Z(n1626) );
  ND2 U19296 ( .A(n4827), .B(n5091), .Z(n3131) );
  ND2 U19297 ( .A(n4938), .B(n5091), .Z(n3132) );
  MUX21L U19298 ( .A(n3290), .B(n5254), .S(n4610), .Z(n1629) );
  ND2 U19299 ( .A(n5254), .B(n4844), .Z(n3290) );
  ND2 U19300 ( .A(n4575), .B(n5129), .Z(n3571) );
  ND2 U19301 ( .A(n4957), .B(n4442), .Z(n3154) );
  ND2 U19302 ( .A(n5235), .B(n4442), .Z(n3155) );
  ND2 U19303 ( .A(n3513), .B(n3512), .Z(n1134) );
  ND2 U19304 ( .A(n5246), .B(n4421), .Z(n3512) );
  EN U19305 ( .A(n4900), .B(n4571), .Z(n3513) );
  ND2 U19306 ( .A(n3180), .B(n3179), .Z(n1129) );
  ND2 U19307 ( .A(n4586), .B(n4833), .Z(n3179) );
  MUX21L U19308 ( .A(n4834), .B(n3178), .S(n5232), .Z(n3180) );
  NR2 U19309 ( .A(n4586), .B(n4833), .Z(n3178) );
  ND2 U19310 ( .A(n3360), .B(n3359), .Z(n1132) );
  ND2 U19311 ( .A(n4605), .B(n5105), .Z(n3359) );
  MUX21L U19312 ( .A(n4792), .B(n3358), .S(n5258), .Z(n3360) );
  NR2 U19313 ( .A(n4605), .B(n4792), .Z(n3358) );
  ND2 U19314 ( .A(n2644), .B(n2643), .Z(n1585) );
  ND2 U19315 ( .A(n5292), .B(n4515), .Z(n2643) );
  EN U19316 ( .A(n4903), .B(n4624), .Z(n2644) );
  NR2 U19317 ( .A(n4548), .B(n4805), .Z(n2937) );
  ND2 U19318 ( .A(n4905), .B(n4503), .Z(n2740) );
  ND2 U19319 ( .A(n3057), .B(n3056), .Z(n1593) );
  ND2 U19320 ( .A(n4942), .B(n4383), .Z(n3056) );
  EO U19321 ( .A(n5221), .B(n4556), .Z(n3057) );
  ND2 U19322 ( .A(n2994), .B(n2993), .Z(n1592) );
  ND2 U19323 ( .A(n5234), .B(n4811), .Z(n2993) );
  MUX21L U19324 ( .A(n2992), .B(n4390), .S(n5234), .Z(n2994) );
  ND2 U19325 ( .A(n2869), .B(n2868), .Z(n1590) );
  ND2 U19326 ( .A(n4565), .B(n4735), .Z(n2868) );
  MUX21L U19327 ( .A(n5283), .B(n2867), .S(n4933), .Z(n2869) );
  NR2 U19328 ( .A(n5283), .B(n4565), .Z(n2867) );
  ND2 U19329 ( .A(n3411), .B(n3410), .Z(n1600) );
  MUX21L U19330 ( .A(n3408), .B(n5111), .S(n4588), .Z(n3410) );
  AO6 U19331 ( .A(n4589), .B(n4788), .C(n3409), .Z(n3411) );
  ND2 U19332 ( .A(n3230), .B(n3229), .Z(n1598) );
  ND2 U19333 ( .A(n4478), .B(n5080), .Z(n3230) );
  ND2 U19334 ( .A(n4953), .B(n5079), .Z(n3229) );
  ND2 U19335 ( .A(n4516), .B(n4895), .Z(n1142) );
  ND2 U19336 ( .A(n3575), .B(n3574), .Z(n1118) );
  ND2 U19337 ( .A(n4925), .B(n4413), .Z(n3574) );
  MUX21L U19338 ( .A(n5129), .B(n3573), .S(n4575), .Z(n3575) );
  NR2 U19339 ( .A(n4925), .B(n5129), .Z(n3573) );
  ND2 U19340 ( .A(n3305), .B(n3304), .Z(n1114) );
  ND2 U19341 ( .A(n5255), .B(n4847), .Z(n3304) );
  MUX21L U19342 ( .A(n4847), .B(n3303), .S(n4609), .Z(n3305) );
  NR2 U19343 ( .A(n5255), .B(n4846), .Z(n3303) );
  ND2 U19344 ( .A(n3455), .B(n3454), .Z(n1116) );
  ND2 U19345 ( .A(n4427), .B(n4783), .Z(n3454) );
  EO U19346 ( .A(n5221), .B(n4591), .Z(n3455) );
  ND2 U19347 ( .A(n3248), .B(n3247), .Z(n1113) );
  ND2 U19348 ( .A(n4613), .B(n4840), .Z(n3247) );
  MUX21L U19349 ( .A(n4613), .B(n3246), .S(n5252), .Z(n3248) );
  NR2 U19350 ( .A(n4613), .B(n4840), .Z(n3246) );
  AO7 U19351 ( .A(n4956), .B(n5090), .C(n4439), .Z(n1596) );
  NR2 U19352 ( .A(n5285), .B(n4395), .Z(n2935) );
  ND2 U19353 ( .A(n5278), .B(n4504), .Z(n2741) );
  AN3 U19354 ( .A(n4487), .B(n4845), .C(n5254), .Z(n778) );
  MUX21L U19355 ( .A(n4954), .B(n4434), .S(n5231), .Z(n1597) );
  MUX21L U19356 ( .A(n3361), .B(n4935), .S(n4605), .Z(n1115) );
  ND2 U19357 ( .A(n4935), .B(n5105), .Z(n3361) );
  ND2 U19358 ( .A(n3235), .B(n3234), .Z(n1572) );
  ND2 U19359 ( .A(n3231), .B(n4839), .Z(n3234) );
  MUX21L U19360 ( .A(n3232), .B(n3233), .S(n4613), .Z(n3235) );
  NR2 U19361 ( .A(n5251), .B(n4613), .Z(n3231) );
  ND2 U19362 ( .A(n3134), .B(n3133), .Z(n1570) );
  ND2 U19363 ( .A(n4375), .B(n4827), .Z(n3133) );
  EN U19364 ( .A(n5224), .B(n4583), .Z(n3134) );
  ND2 U19365 ( .A(n3109), .B(n3108), .Z(n1568) );
  ND2 U19366 ( .A(n4581), .B(n4824), .Z(n3108) );
  EO U19367 ( .A(n5223), .B(n4581), .Z(n3109) );
  ND2 U19368 ( .A(n4414), .B(n5128), .Z(n3572) );
  NR2 U19369 ( .A(n4953), .B(n5079), .Z(n3233) );
  ND2 U19370 ( .A(n4748), .B(n5196), .Z(n2769) );
  ND2 U19371 ( .A(n3438), .B(n3437), .Z(n1574) );
  ND2 U19372 ( .A(n4590), .B(n4784), .Z(n3437) );
  EO U19373 ( .A(n5221), .B(n4590), .Z(n3438) );
  ND2 U19374 ( .A(n3547), .B(n4417), .Z(n1575) );
  ND2 U19375 ( .A(n5247), .B(n4924), .Z(n3547) );
  ND2 U19376 ( .A(n2825), .B(n2824), .Z(n1563) );
  ND2 U19377 ( .A(n4930), .B(n4406), .Z(n2824) );
  MUX21L U19378 ( .A(n2823), .B(n4406), .S(n5281), .Z(n2825) );
  NR2 U19379 ( .A(n4930), .B(n4405), .Z(n2823) );
  ND2 U19380 ( .A(n2871), .B(n2870), .Z(n1564) );
  ND2 U19381 ( .A(n5284), .B(n4401), .Z(n2871) );
  ND2 U19382 ( .A(n4933), .B(n4400), .Z(n2870) );
  AN3 U19383 ( .A(n4610), .B(n4845), .C(n5254), .Z(n779) );
  MUX21L U19384 ( .A(n4816), .B(n3043), .S(n5237), .Z(n1567) );
  ND2 U19385 ( .A(n4554), .B(n4817), .Z(n3043) );
  MUX21L U19386 ( .A(n2941), .B(n2940), .S(n4548), .Z(n1565) );
  ND2 U19387 ( .A(n4805), .B(n5184), .Z(n2940) );
  ND2 U19388 ( .A(n5285), .B(n4948), .Z(n2941) );
  ND2 U19389 ( .A(n3282), .B(n4485), .Z(n1104) );
  ND2 U19390 ( .A(n5254), .B(n4950), .Z(n3282) );
  ND2 U19391 ( .A(n3137), .B(n3136), .Z(n1549) );
  ND2 U19392 ( .A(n4583), .B(n4827), .Z(n3136) );
  MUX21L U19393 ( .A(n5238), .B(n3135), .S(n4938), .Z(n3137) );
  NR2 U19394 ( .A(n5237), .B(n4583), .Z(n3135) );
  ND2 U19395 ( .A(n3620), .B(n3619), .Z(n1556) );
  ND2 U19396 ( .A(n4578), .B(n5132), .Z(n3619) );
  EO U19397 ( .A(n5227), .B(n4927), .Z(n3620) );
  ND2 U19398 ( .A(n3199), .B(n3198), .Z(n1550) );
  ND2 U19399 ( .A(n4835), .B(n5084), .Z(n3198) );
  MUX21L U19400 ( .A(n5084), .B(n3197), .S(n4587), .Z(n3199) );
  ND2 U19401 ( .A(n3424), .B(n3423), .Z(n1107) );
  MUX21L U19402 ( .A(n3421), .B(n5112), .S(n4918), .Z(n3423) );
  AO6 U19403 ( .A(n4918), .B(n4428), .C(n3422), .Z(n3424) );
  ND2 U19404 ( .A(n2978), .B(n4393), .Z(n1546) );
  ND2 U19405 ( .A(n5232), .B(n4946), .Z(n2978) );
  ND2 U19406 ( .A(n2997), .B(n2996), .Z(n1547) );
  ND2 U19407 ( .A(n4945), .B(n4390), .Z(n2996) );
  MUX21L U19408 ( .A(n2995), .B(n4390), .S(n5234), .Z(n2997) );
  NR2 U19409 ( .A(n4945), .B(n4389), .Z(n2995) );
  ND2 U19410 ( .A(n4795), .B(n5104), .Z(n3340) );
  ND2 U19411 ( .A(n5246), .B(n4421), .Z(n3515) );
  MUX21L U19412 ( .A(n3292), .B(n3291), .S(n4610), .Z(n1552) );
  ND2 U19413 ( .A(n4845), .B(n5075), .Z(n3291) );
  ND2 U19414 ( .A(n4949), .B(n5075), .Z(n3292) );
  MUX21L U19415 ( .A(n4430), .B(n5242), .S(n4918), .Z(n1554) );
  MUX21L U19416 ( .A(n4606), .B(n3341), .S(n5257), .Z(n1553) );
  ND2 U19417 ( .A(n4606), .B(n4794), .Z(n3341) );
  NR2 U19418 ( .A(n5251), .B(n4479), .Z(n3236) );
  ND2 U19419 ( .A(n3316), .B(n3315), .Z(n1535) );
  ND2 U19420 ( .A(n4488), .B(n4848), .Z(n3315) );
  EO U19421 ( .A(n5224), .B(n4608), .Z(n3316) );
  ND2 U19422 ( .A(n3239), .B(n3238), .Z(n1534) );
  AO6 U19423 ( .A(n5251), .B(n4479), .C(n3237), .Z(n3239) );
  MUX21L U19424 ( .A(n5251), .B(n3236), .S(n4953), .Z(n3238) );
  NR2 U19425 ( .A(n4953), .B(n4613), .Z(n3237) );
  ND2 U19426 ( .A(n4408), .B(n4741), .Z(n1562) );
  IVP U19427 ( .A(n5067), .Z(n5243) );
  NR2 U19428 ( .A(n4919), .B(n4428), .Z(n3439) );
  ND2 U19429 ( .A(n3444), .B(n3443), .Z(n1537) );
  MUX21L U19430 ( .A(n3441), .B(n3442), .S(n4919), .Z(n3443) );
  MUX21L U19431 ( .A(n3439), .B(n3440), .S(n5243), .Z(n3444) );
  NR2 U19432 ( .A(n4590), .B(n5113), .Z(n3441) );
  ND2 U19433 ( .A(n3139), .B(n3138), .Z(n1532) );
  ND2 U19434 ( .A(n5237), .B(n4426), .Z(n3139) );
  ND2 U19435 ( .A(n4938), .B(n4443), .Z(n3138) );
  MUX21L U19436 ( .A(n5130), .B(n3576), .S(n4575), .Z(n3578) );
  NR2 U19437 ( .A(n4925), .B(n5130), .Z(n3576) );
  ND2 U19438 ( .A(n3296), .B(n3295), .Z(n1522) );
  MUX21L U19439 ( .A(n3293), .B(n5074), .S(n4949), .Z(n3295) );
  AO6 U19440 ( .A(n4949), .B(n4487), .C(n3294), .Z(n3296) );
  ND2 U19441 ( .A(n3496), .B(n3495), .Z(n1525) );
  MUX21L U19442 ( .A(n5245), .B(n3493), .S(n4921), .Z(n3495) );
  AO6 U19443 ( .A(n5245), .B(n4424), .C(n3494), .Z(n3496) );
  NR2 U19444 ( .A(n5245), .B(n4424), .Z(n3493) );
  ND2 U19445 ( .A(n4925), .B(n5130), .Z(n3577) );
  MUX21L U19446 ( .A(n4771), .B(n3579), .S(n5249), .Z(n3581) );
  NR2 U19447 ( .A(n4576), .B(n4771), .Z(n3579) );
  ND3 U19448 ( .A(n4577), .B(n5132), .C(n4927), .Z(n1526) );
  ND2 U19449 ( .A(n4423), .B(n4780), .Z(n3498) );
  ND2 U19450 ( .A(n4921), .B(n4423), .Z(n3497) );
  ND2 U19451 ( .A(n3533), .B(n3532), .Z(n1508) );
  ND2 U19452 ( .A(n4572), .B(n4923), .Z(n3532) );
  MUX21L U19453 ( .A(n3531), .B(n5123), .S(n4923), .Z(n3533) );
  NR2 U19454 ( .A(n4573), .B(n5124), .Z(n3531) );
  ND2 U19455 ( .A(n3449), .B(n3448), .Z(n1507) );
  MUX21L U19456 ( .A(n4784), .B(n3445), .S(n5243), .Z(n3448) );
  NR2 U19457 ( .A(n3447), .B(n3446), .Z(n3449) );
  ND2 U19458 ( .A(n4793), .B(n5104), .Z(n3343) );
  ND2 U19459 ( .A(n3501), .B(n3500), .Z(n1503) );
  ND2 U19460 ( .A(n4570), .B(n4780), .Z(n3500) );
  MUX21L U19461 ( .A(n4570), .B(n3499), .S(n5245), .Z(n3501) );
  NR2 U19462 ( .A(n4570), .B(n4779), .Z(n3499) );
  ND2 U19463 ( .A(n4925), .B(n4413), .Z(n3582) );
  ND2 U19464 ( .A(n4415), .B(n4774), .Z(n3562) );
  ND2 U19465 ( .A(n4574), .B(n4774), .Z(n3561) );
  ND2 U19466 ( .A(n3604), .B(n3603), .Z(n1499) );
  NR2 U19467 ( .A(n3602), .B(n3601), .Z(n3604) );
  MUX21L U19468 ( .A(n4769), .B(n3600), .S(n5250), .Z(n3603) );
  NR2 U19469 ( .A(n5250), .B(n4577), .Z(n3602) );
  NR2 U19470 ( .A(n4960), .B(n4536), .Z(n2330) );
  NR2 U19471 ( .A(n4633), .B(n5147), .Z(n2332) );
  NR2 U19472 ( .A(n4926), .B(n5132), .Z(n3591) );
  OR3 U19473 ( .A(n4557), .B(n5295), .C(n4908), .Z(n780) );
  ND2 U19474 ( .A(n3589), .B(n4769), .Z(n3592) );
  MUX21L U19475 ( .A(n3590), .B(n3591), .S(n4576), .Z(n3593) );
  AO6 U19476 ( .A(n4601), .B(n4852), .C(n2103), .Z(n2105) );
  NR2 U19477 ( .A(n5272), .B(n4911), .Z(n2103) );
  ND2 U19478 ( .A(n3365), .B(n3364), .Z(n1083) );
  MUX21L U19479 ( .A(n3362), .B(n5106), .S(n4936), .Z(n3364) );
  AO6 U19480 ( .A(n4936), .B(n4492), .C(n3363), .Z(n3365) );
  NR2 U19481 ( .A(n4966), .B(n4466), .Z(n2213) );
  NR2 U19482 ( .A(n5241), .B(n4379), .Z(n3095) );
  NR2 U19483 ( .A(n4954), .B(n4433), .Z(n3208) );
  NR2 U19484 ( .A(n4633), .B(n4877), .Z(n2339) );
  NR2 U19485 ( .A(n4959), .B(n5147), .Z(n2340) );
  NR2 U19486 ( .A(n5267), .B(n4527), .Z(n2459) );
  NR2 U19487 ( .A(n5287), .B(n4476), .Z(n2498) );
  NR2 U19488 ( .A(n5265), .B(n4883), .Z(n2403) );
  NR2 U19489 ( .A(n4567), .B(n4798), .Z(n2902) );
  NR2 U19490 ( .A(n4934), .B(n5186), .Z(n2903) );
  NR2 U19491 ( .A(n4588), .B(n5082), .Z(n3213) );
  NR2 U19492 ( .A(n5250), .B(n4837), .Z(n3214) );
  NR2 U19493 ( .A(n4919), .B(n5112), .Z(n3431) );
  ND2 U19494 ( .A(n5262), .B(n4876), .Z(n2337) );
  ND2 U19495 ( .A(n4633), .B(n5262), .Z(n2338) );
  ND2 U19496 ( .A(n4633), .B(n4876), .Z(n2336) );
  ND2 U19497 ( .A(n3522), .B(n3521), .Z(n1025) );
  ND2 U19498 ( .A(n4572), .B(n4777), .Z(n3521) );
  EN U19499 ( .A(n5229), .B(n4922), .Z(n3522) );
  ND2 U19500 ( .A(n2300), .B(n2299), .Z(n938) );
  ND2 U19501 ( .A(n4540), .B(n5150), .Z(n2299) );
  EO U19502 ( .A(n4900), .B(n4630), .Z(n2300) );
  ND2 U19503 ( .A(n2686), .B(n2685), .Z(n947) );
  ND2 U19504 ( .A(n5293), .B(n4614), .Z(n2685) );
  EN U19505 ( .A(n5225), .B(n4906), .Z(n2686) );
  ND2 U19506 ( .A(n3634), .B(n4410), .Z(n931) );
  EO U19507 ( .A(n5227), .B(n4923), .Z(n3634) );
  ND2 U19508 ( .A(n4592), .B(n4759), .Z(n2496) );
  ND2 U19509 ( .A(n2549), .B(n5216), .Z(n2552) );
  NR2 U19510 ( .A(n4619), .B(n4975), .Z(n2549) );
  ND2 U19511 ( .A(n5275), .B(n4466), .Z(n2218) );
  ND2 U19512 ( .A(n4966), .B(n4467), .Z(n2217) );
  ND2 U19513 ( .A(n5289), .B(n4523), .Z(n2574) );
  ND2 U19514 ( .A(n2495), .B(n2494), .Z(n1066) );
  ND2 U19515 ( .A(n4592), .B(n5134), .Z(n2494) );
  EN U19516 ( .A(n4897), .B(n4592), .Z(n2495) );
  ND2 U19517 ( .A(n2548), .B(n2547), .Z(n1067) );
  ND2 U19518 ( .A(n4975), .B(n5216), .Z(n2547) );
  MUX21L U19519 ( .A(n2546), .B(n4524), .S(n4975), .Z(n2548) );
  ND2 U19520 ( .A(n2416), .B(n2415), .Z(n1064) );
  ND2 U19521 ( .A(n4529), .B(n5139), .Z(n2415) );
  EO U19522 ( .A(n4900), .B(n4614), .Z(n2416) );
  ND2 U19523 ( .A(n3097), .B(n3096), .Z(n1077) );
  ND3 U19524 ( .A(n4940), .B(n4379), .C(n5235), .Z(n3096) );
  MUX21L U19525 ( .A(n3094), .B(n3095), .S(n4940), .Z(n3097) );
  ND2 U19526 ( .A(n3031), .B(n4387), .Z(n1076) );
  EO U19527 ( .A(n5230), .B(n4943), .Z(n3031) );
  ND2 U19528 ( .A(n3616), .B(n3615), .Z(n1086) );
  MUX21L U19529 ( .A(n4768), .B(n3612), .S(n5250), .Z(n3615) );
  NR2 U19530 ( .A(n3614), .B(n3613), .Z(n3616) );
  ND2 U19531 ( .A(n3394), .B(n3393), .Z(n1053) );
  ND2 U19532 ( .A(n4494), .B(n5110), .Z(n3393) );
  EO U19533 ( .A(n4898), .B(n4603), .Z(n3394) );
  ND2 U19534 ( .A(n3206), .B(n5082), .Z(n1050) );
  EN U19535 ( .A(n4901), .B(n4588), .Z(n3206) );
  ND2 U19536 ( .A(n2849), .B(n2848), .Z(n1042) );
  ND2 U19537 ( .A(n4564), .B(n4737), .Z(n2848) );
  EO U19538 ( .A(n5229), .B(n4564), .Z(n2849) );
  ND2 U19539 ( .A(n2155), .B(n2154), .Z(n998) );
  ND2 U19540 ( .A(n4765), .B(n5164), .Z(n2154) );
  MUX21L U19541 ( .A(n5164), .B(n2153), .S(n4599), .Z(n2155) );
  ND2 U19542 ( .A(n3308), .B(n3307), .Z(n1022) );
  ND2 U19543 ( .A(n4949), .B(n5072), .Z(n3307) );
  MUX21L U19544 ( .A(n3306), .B(n4488), .S(n4949), .Z(n3308) );
  ND2 U19545 ( .A(n2901), .B(n2900), .Z(n1013) );
  ND2 U19546 ( .A(n4798), .B(n5187), .Z(n2900) );
  MUX21L U19547 ( .A(n4798), .B(n2899), .S(n4567), .Z(n2901) );
  ND2 U19548 ( .A(n3073), .B(n3072), .Z(n1016) );
  ND2 U19549 ( .A(n4820), .B(n5097), .Z(n3072) );
  MUX21L U19550 ( .A(n4820), .B(n3071), .S(n4556), .Z(n3073) );
  ND2 U19551 ( .A(n2953), .B(n2952), .Z(n1014) );
  ND2 U19552 ( .A(n5286), .B(n4807), .Z(n2952) );
  MUX21L U19553 ( .A(n2951), .B(n4395), .S(n5286), .Z(n2953) );
  ND2 U19554 ( .A(n2799), .B(n2798), .Z(n981) );
  ND2 U19555 ( .A(n4929), .B(n4392), .Z(n2798) );
  EO U19556 ( .A(n5222), .B(n4561), .Z(n2799) );
  ND2 U19557 ( .A(n3018), .B(n3017), .Z(n985) );
  ND2 U19558 ( .A(n5240), .B(n4944), .Z(n3017) );
  MUX21L U19559 ( .A(n3016), .B(n4388), .S(n4944), .Z(n3018) );
  NR2 U19560 ( .A(n5240), .B(n4388), .Z(n3016) );
  ND2 U19561 ( .A(n2287), .B(n2286), .Z(n970) );
  MUX21L U19562 ( .A(n2284), .B(n2285), .S(n4629), .Z(n2287) );
  ND2 U19563 ( .A(n2283), .B(n5152), .Z(n2286) );
  NR2 U19564 ( .A(n5260), .B(n4872), .Z(n2285) );
  ND2 U19565 ( .A(n2501), .B(n2500), .Z(n976) );
  AO6 U19566 ( .A(n5287), .B(n4476), .C(n2499), .Z(n2501) );
  MUX21L U19567 ( .A(n5287), .B(n2498), .S(n4917), .Z(n2500) );
  NR2 U19568 ( .A(n4917), .B(n4592), .Z(n2499) );
  ND2 U19569 ( .A(n2633), .B(n2632), .Z(n978) );
  ND2 U19570 ( .A(n4893), .B(n5210), .Z(n2632) );
  MUX21L U19571 ( .A(n5210), .B(n2631), .S(n4624), .Z(n2633) );
  ND2 U19572 ( .A(n2418), .B(n2417), .Z(n942) );
  ND2 U19573 ( .A(n4529), .B(n5139), .Z(n2417) );
  EO U19574 ( .A(n4899), .B(n4615), .Z(n2418) );
  ND2 U19575 ( .A(n3217), .B(n3216), .Z(n958) );
  NR2 U19576 ( .A(n3215), .B(n3214), .Z(n3217) );
  MUX21L U19577 ( .A(n3213), .B(n4588), .S(n4953), .Z(n3216) );
  NR2 U19578 ( .A(n5250), .B(n4433), .Z(n3215) );
  ND2 U19579 ( .A(n3005), .B(n3004), .Z(n921) );
  ND2 U19580 ( .A(n4552), .B(n4812), .Z(n3004) );
  MUX21L U19581 ( .A(n4812), .B(n3003), .S(n5236), .Z(n3005) );
  NR2 U19582 ( .A(n4552), .B(n4811), .Z(n3003) );
  ND2 U19583 ( .A(n3538), .B(n3537), .Z(n930) );
  ND2 U19584 ( .A(n5247), .B(n4418), .Z(n3537) );
  EO U19585 ( .A(n4901), .B(n4573), .Z(n3538) );
  ND2 U19586 ( .A(n2607), .B(n2606), .Z(n912) );
  ND2 U19587 ( .A(n4623), .B(n5211), .Z(n2606) );
  EN U19588 ( .A(n4901), .B(n4623), .Z(n2607) );
  ND2 U19589 ( .A(n2666), .B(n2665), .Z(n913) );
  ND2 U19590 ( .A(n4970), .B(n4512), .Z(n2665) );
  MUX21L U19591 ( .A(n2664), .B(n4512), .S(n5293), .Z(n2666) );
  NR2 U19592 ( .A(n4970), .B(n4512), .Z(n2664) );
  ND2 U19593 ( .A(n2707), .B(n2706), .Z(n914) );
  ND2 U19594 ( .A(n4908), .B(n4506), .Z(n2706) );
  MUX21L U19595 ( .A(n2705), .B(n4507), .S(n5295), .Z(n2707) );
  NR2 U19596 ( .A(n4908), .B(n4506), .Z(n2705) );
  ND2 U19597 ( .A(n3251), .B(n3250), .Z(n895) );
  ND2 U19598 ( .A(n5252), .B(n4841), .Z(n3250) );
  MUX21L U19599 ( .A(n4841), .B(n3249), .S(n4612), .Z(n3251) );
  NR2 U19600 ( .A(n5252), .B(n4841), .Z(n3249) );
  ND2 U19601 ( .A(n3433), .B(n3432), .Z(n898) );
  ND2 U19602 ( .A(n3429), .B(n4785), .Z(n3432) );
  MUX21L U19603 ( .A(n3430), .B(n3431), .S(n4589), .Z(n3433) );
  NR2 U19604 ( .A(n5243), .B(n4590), .Z(n3429) );
  ND2 U19605 ( .A(n3052), .B(n3051), .Z(n890) );
  ND2 U19606 ( .A(n5232), .B(n4384), .Z(n3051) );
  EN U19607 ( .A(n4897), .B(n4555), .Z(n3052) );
  ND2 U19608 ( .A(n4535), .B(n4877), .Z(n2348) );
  ND2 U19609 ( .A(n4959), .B(n4633), .Z(n2347) );
  MUX21L U19610 ( .A(n2102), .B(n5168), .S(n4602), .Z(n2104) );
  MUX21L U19611 ( .A(n2550), .B(n2551), .S(n4619), .Z(n2553) );
  NR2 U19612 ( .A(n5289), .B(n4885), .Z(n2551) );
  ND2 U19613 ( .A(n2780), .B(n2779), .Z(n1072) );
  ND2 U19614 ( .A(n5279), .B(n4745), .Z(n2779) );
  MUX21L U19615 ( .A(n2778), .B(n4496), .S(n5279), .Z(n2780) );
  ND2 U19616 ( .A(n2062), .B(n2061), .Z(n997) );
  ND2 U19617 ( .A(n4627), .B(n5172), .Z(n2061) );
  MUX21L U19618 ( .A(n2060), .B(n5172), .S(n4909), .Z(n2062) );
  NR2 U19619 ( .A(n4627), .B(n5171), .Z(n2060) );
  ND2 U19620 ( .A(n2298), .B(n2297), .Z(n1001) );
  ND2 U19621 ( .A(n4962), .B(n4630), .Z(n2297) );
  MUX21L U19622 ( .A(n2296), .B(n5151), .S(n4630), .Z(n2298) );
  NR2 U19623 ( .A(n4962), .B(n5151), .Z(n2296) );
  ND2 U19624 ( .A(n2343), .B(n2342), .Z(n971) );
  NR2 U19625 ( .A(n2341), .B(n2340), .Z(n2343) );
  MUX21L U19626 ( .A(n2339), .B(n4633), .S(n5262), .Z(n2342) );
  NR2 U19627 ( .A(n4959), .B(n4536), .Z(n2341) );
  ND2 U19628 ( .A(n2255), .B(n2254), .Z(n969) );
  ND2 U19629 ( .A(n4594), .B(n4869), .Z(n2254) );
  MUX21L U19630 ( .A(n5277), .B(n2253), .S(n4964), .Z(n2255) );
  NR2 U19631 ( .A(n5277), .B(n4594), .Z(n2253) );
  ND2 U19632 ( .A(n2663), .B(n2662), .Z(n979) );
  ND2 U19633 ( .A(n5293), .B(n4802), .Z(n2662) );
  MUX21L U19634 ( .A(n2661), .B(n4513), .S(n5293), .Z(n2663) );
  ND2 U19635 ( .A(n2405), .B(n2404), .Z(n974) );
  ND2 U19636 ( .A(n2401), .B(n5139), .Z(n2404) );
  MUX21L U19637 ( .A(n2402), .B(n2403), .S(n4637), .Z(n2405) );
  NR2 U19638 ( .A(n4637), .B(n4976), .Z(n2401) );
  ND2 U19639 ( .A(n2188), .B(n2187), .Z(n936) );
  ND2 U19640 ( .A(n4597), .B(n4863), .Z(n2187) );
  MUX21L U19641 ( .A(n4597), .B(n2186), .S(n5275), .Z(n2188) );
  NR2 U19642 ( .A(n4597), .B(n4863), .Z(n2186) );
  ND2 U19643 ( .A(n2108), .B(n2107), .Z(n934) );
  ND2 U19644 ( .A(n4912), .B(n4456), .Z(n2107) );
  MUX21L U19645 ( .A(n2106), .B(n4456), .S(n5272), .Z(n2108) );
  NR2 U19646 ( .A(n4912), .B(n4456), .Z(n2106) );
  ND2 U19647 ( .A(n2556), .B(n2555), .Z(n945) );
  ND2 U19648 ( .A(n4620), .B(n4886), .Z(n2555) );
  MUX21L U19649 ( .A(n4886), .B(n2554), .S(n5289), .Z(n2556) );
  NR2 U19650 ( .A(n4620), .B(n4885), .Z(n2554) );
  ND2 U19651 ( .A(n2906), .B(n2905), .Z(n953) );
  NR2 U19652 ( .A(n2904), .B(n2903), .Z(n2906) );
  MUX21L U19653 ( .A(n2902), .B(n4567), .S(n5285), .Z(n2905) );
  NR2 U19654 ( .A(n4934), .B(n4398), .Z(n2904) );
  ND2 U19655 ( .A(n3050), .B(n3049), .Z(n956) );
  ND2 U19656 ( .A(n4555), .B(n5099), .Z(n3049) );
  MUX21L U19657 ( .A(n3048), .B(n5099), .S(n4942), .Z(n3050) );
  NR2 U19658 ( .A(n4555), .B(n5098), .Z(n3048) );
  ND2 U19659 ( .A(n2970), .B(n2969), .Z(n920) );
  ND2 U19660 ( .A(n4550), .B(n4946), .Z(n2969) );
  MUX21L U19661 ( .A(n2968), .B(n5181), .S(n4946), .Z(n2970) );
  NR2 U19662 ( .A(n4549), .B(n5181), .Z(n2968) );
  ND2 U19663 ( .A(n2752), .B(n2751), .Z(n916) );
  ND2 U19664 ( .A(n4904), .B(n4500), .Z(n2751) );
  MUX21L U19665 ( .A(n2750), .B(n4501), .S(n5278), .Z(n2752) );
  NR2 U19666 ( .A(n4905), .B(n4500), .Z(n2750) );
  ND2 U19667 ( .A(n3428), .B(n3427), .Z(n929) );
  ND2 U19668 ( .A(n5243), .B(n4786), .Z(n3427) );
  MUX21L U19669 ( .A(n4786), .B(n3426), .S(n4589), .Z(n3428) );
  NR2 U19670 ( .A(n5243), .B(n4786), .Z(n3426) );
  ND2 U19671 ( .A(n3525), .B(n3524), .Z(n899) );
  ND2 U19672 ( .A(n4922), .B(n5122), .Z(n3524) );
  MUX21L U19673 ( .A(n3523), .B(n4420), .S(n4922), .Z(n3525) );
  ND2 U19674 ( .A(n3160), .B(n3159), .Z(n893) );
  ND2 U19675 ( .A(n4957), .B(n4440), .Z(n3159) );
  MUX21L U19676 ( .A(n3158), .B(n4441), .S(n5234), .Z(n3160) );
  NR2 U19677 ( .A(n4957), .B(n4440), .Z(n3158) );
  ND2 U19678 ( .A(n3100), .B(n3099), .Z(n891) );
  ND2 U19679 ( .A(n4939), .B(n4378), .Z(n3099) );
  MUX21L U19680 ( .A(n3098), .B(n4378), .S(n5241), .Z(n3100) );
  NR2 U19681 ( .A(n4939), .B(n4377), .Z(n3098) );
  ND2 U19682 ( .A(n3373), .B(n3372), .Z(n872) );
  ND2 U19683 ( .A(n4604), .B(n4791), .Z(n3372) );
  MUX21L U19684 ( .A(n4604), .B(n3371), .S(n5258), .Z(n3373) );
  NR2 U19685 ( .A(n4604), .B(n4790), .Z(n3371) );
  ND2 U19686 ( .A(n3311), .B(n3310), .Z(n871) );
  ND2 U19687 ( .A(n4609), .B(n4848), .Z(n3310) );
  MUX21L U19688 ( .A(n4609), .B(n3309), .S(n5255), .Z(n3311) );
  NR2 U19689 ( .A(n4609), .B(n4847), .Z(n3309) );
  ND2 U19690 ( .A(n2365), .B(n2364), .Z(n1035) );
  ND2 U19691 ( .A(n5263), .B(n4533), .Z(n2364) );
  MUX21L U19692 ( .A(n4879), .B(n2363), .S(n4634), .Z(n2365) );
  NR2 U19693 ( .A(n5263), .B(n4879), .Z(n2363) );
  ND2 U19694 ( .A(n2369), .B(n2368), .Z(n1004) );
  MUX21L U19695 ( .A(n2366), .B(n5145), .S(n4978), .Z(n2368) );
  AO6 U19696 ( .A(n4978), .B(n4533), .C(n2367), .Z(n2369) );
  AO7 U19697 ( .A(n4939), .B(n4376), .C(n3114), .Z(n1047) );
  ND2 U19698 ( .A(n5239), .B(n4582), .Z(n3114) );
  AO7 U19699 ( .A(n4591), .B(n5114), .C(n3456), .Z(n1024) );
  ND2 U19700 ( .A(n5241), .B(n4919), .Z(n3456) );
  AO7 U19701 ( .A(n4576), .B(n4770), .C(n5249), .Z(n1026) );
  AO7 U19702 ( .A(n5281), .B(n4404), .C(n4931), .Z(n1012) );
  AO7 U19703 ( .A(n4948), .B(n4489), .C(n3327), .Z(n991) );
  ND2 U19704 ( .A(n5256), .B(n4607), .Z(n3327) );
  AO7 U19705 ( .A(n4624), .B(n4893), .C(n2634), .Z(n946) );
  ND2 U19706 ( .A(n5291), .B(n4971), .Z(n2634) );
  AO7 U19707 ( .A(n5247), .B(n4418), .C(n3536), .Z(n962) );
  ND2 U19708 ( .A(n4923), .B(n4573), .Z(n3536) );
  AO7 U19709 ( .A(n4580), .B(n5096), .C(n4821), .Z(n922) );
  AO7 U19710 ( .A(n4936), .B(n4603), .C(n5108), .Z(n928) );
  NR2 U19711 ( .A(n4617), .B(n4762), .Z(n2461) );
  NR2 U19712 ( .A(n4955), .B(n5087), .Z(n1080) );
  ND2 U19713 ( .A(n2383), .B(n2382), .Z(n1063) );
  ND2 U19714 ( .A(n4636), .B(n5142), .Z(n2382) );
  EO U19715 ( .A(n5223), .B(n4978), .Z(n2383) );
  ND3 U19716 ( .A(n3464), .B(n3463), .C(n3462), .Z(n1054) );
  ND2 U19717 ( .A(n4919), .B(n5115), .Z(n3464) );
  ND2 U19718 ( .A(n4568), .B(n5115), .Z(n3463) );
  ND2 U19719 ( .A(n4919), .B(n4568), .Z(n3462) );
  ND3 U19720 ( .A(n4425), .B(n5116), .C(n4920), .Z(n993) );
  ND3 U19721 ( .A(n2887), .B(n2886), .C(n2885), .Z(n919) );
  ND2 U19722 ( .A(n4800), .B(n5187), .Z(n2886) );
  ND2 U19723 ( .A(n4566), .B(n5188), .Z(n2887) );
  ND2 U19724 ( .A(n4566), .B(n4800), .Z(n2885) );
  ND2 U19725 ( .A(n2413), .B(n2412), .Z(n1005) );
  ND2 U19726 ( .A(n4529), .B(n4884), .Z(n2412) );
  EO U19727 ( .A(n5224), .B(n4976), .Z(n2413) );
  ND2 U19728 ( .A(n4947), .B(n5182), .Z(n2954) );
  ND2 U19729 ( .A(n4947), .B(n4394), .Z(n2955) );
  ND2 U19730 ( .A(n4959), .B(n4536), .Z(n2344) );
  ND2 U19731 ( .A(n5262), .B(n4535), .Z(n2345) );
  ND2 U19732 ( .A(n4909), .B(n4450), .Z(n2065) );
  ND2 U19733 ( .A(n5270), .B(n4450), .Z(n2066) );
  ND2 U19734 ( .A(n2716), .B(n2715), .Z(n1069) );
  ND2 U19735 ( .A(n5295), .B(n4558), .Z(n2716) );
  ND2 U19736 ( .A(n4907), .B(n4558), .Z(n2715) );
  ND2 U19737 ( .A(n4969), .B(n4398), .Z(n1074) );
  ND2 U19738 ( .A(n3032), .B(n4386), .Z(n1045) );
  ND2 U19739 ( .A(n5240), .B(n4943), .Z(n3032) );
  ND3 U19740 ( .A(n2185), .B(n2184), .C(n2183), .Z(n999) );
  ND2 U19741 ( .A(n4464), .B(n4862), .Z(n2184) );
  ND2 U19742 ( .A(n5274), .B(n4862), .Z(n2185) );
  ND2 U19743 ( .A(n5274), .B(n4464), .Z(n2183) );
  ND3 U19744 ( .A(n3268), .B(n3267), .C(n3266), .Z(n1021) );
  ND2 U19745 ( .A(n5253), .B(n4482), .Z(n3267) );
  ND2 U19746 ( .A(n4951), .B(n5253), .Z(n3268) );
  ND2 U19747 ( .A(n4951), .B(n4483), .Z(n3266) );
  ND2 U19748 ( .A(n3172), .B(n4438), .Z(n1019) );
  ND2 U19749 ( .A(n5232), .B(n4956), .Z(n3172) );
  ND2 U19750 ( .A(n2807), .B(n4409), .Z(n1011) );
  ND2 U19751 ( .A(n5280), .B(n4930), .Z(n2807) );
  ND2 U19752 ( .A(n2064), .B(n2063), .Z(n965) );
  ND2 U19753 ( .A(n5270), .B(n4857), .Z(n2064) );
  ND2 U19754 ( .A(n4627), .B(n4856), .Z(n2063) );
  ND2 U19755 ( .A(n2148), .B(n2147), .Z(n967) );
  ND2 U19756 ( .A(n4913), .B(n4460), .Z(n2148) );
  ND2 U19757 ( .A(n4913), .B(n5165), .Z(n2147) );
  ND3 U19758 ( .A(n3586), .B(n3585), .C(n3584), .Z(n963) );
  ND2 U19759 ( .A(n4412), .B(n5131), .Z(n3585) );
  ND2 U19760 ( .A(n4926), .B(n5131), .Z(n3586) );
  ND2 U19761 ( .A(n4926), .B(n4412), .Z(n3584) );
  ND3 U19762 ( .A(n3183), .B(n3182), .C(n3181), .Z(n926) );
  ND2 U19763 ( .A(n4435), .B(n5086), .Z(n3182) );
  ND2 U19764 ( .A(n4955), .B(n5086), .Z(n3183) );
  ND2 U19765 ( .A(n4955), .B(n4435), .Z(n3181) );
  ND2 U19766 ( .A(n2386), .B(n4531), .Z(n907) );
  ND2 U19767 ( .A(n5264), .B(n4977), .Z(n2386) );
  ND2 U19768 ( .A(n2585), .B(n4522), .Z(n911) );
  ND2 U19769 ( .A(n5290), .B(n4973), .Z(n2585) );
  ND2 U19770 ( .A(n3588), .B(n3587), .Z(n900) );
  ND2 U19771 ( .A(n4412), .B(n4770), .Z(n3588) );
  ND2 U19772 ( .A(n5249), .B(n4770), .Z(n3587) );
  ND2 U19773 ( .A(n3033), .B(n4386), .Z(n889) );
  ND2 U19774 ( .A(n5240), .B(n4943), .Z(n3033) );
  ND2 U19775 ( .A(n2855), .B(n4403), .Z(n887) );
  ND2 U19776 ( .A(n5282), .B(n4932), .Z(n2855) );
  AN3 U19777 ( .A(n4818), .B(n5099), .C(n4555), .Z(n781) );
  MUX21L U19778 ( .A(n2250), .B(n5277), .S(n4594), .Z(n1061) );
  ND2 U19779 ( .A(n5276), .B(n4868), .Z(n2250) );
  MUX21L U19780 ( .A(n2677), .B(n4510), .S(n5293), .Z(n1068) );
  ND2 U19781 ( .A(n4969), .B(n4511), .Z(n2677) );
  MUX21L U19782 ( .A(n4807), .B(n2950), .S(n5286), .Z(n1075) );
  ND2 U19783 ( .A(n4549), .B(n4807), .Z(n2950) );
  MUX21L U19784 ( .A(n2749), .B(n2748), .S(n4905), .Z(n1071) );
  ND2 U19785 ( .A(n4501), .B(n5198), .Z(n2748) );
  ND2 U19786 ( .A(n5278), .B(n4501), .Z(n2749) );
  MUX21L U19787 ( .A(n2847), .B(n5190), .S(n4931), .Z(n1073) );
  ND2 U19788 ( .A(n4564), .B(n5191), .Z(n2847) );
  MUX21L U19789 ( .A(n5073), .B(n4949), .S(n4609), .Z(n1082) );
  MUX21L U19790 ( .A(n3520), .B(n3519), .S(n4571), .Z(n1085) );
  ND2 U19791 ( .A(n4777), .B(n5121), .Z(n3519) );
  ND2 U19792 ( .A(n4922), .B(n5121), .Z(n3520) );
  MUX21L U19793 ( .A(n4787), .B(n3425), .S(n4589), .Z(n1084) );
  ND2 U19794 ( .A(n5243), .B(n4787), .Z(n3425) );
  MUX21L U19795 ( .A(n5122), .B(n4572), .S(n4922), .Z(n1055) );
  MUX21L U19796 ( .A(n3157), .B(n3156), .S(n5235), .Z(n1049) );
  ND2 U19797 ( .A(n4441), .B(n4830), .Z(n3157) );
  ND2 U19798 ( .A(n4957), .B(n4441), .Z(n3156) );
  MUX21L U19799 ( .A(n4840), .B(n4612), .S(n5252), .Z(n1051) );
  MUX21L U19800 ( .A(n5096), .B(n4821), .S(n4579), .Z(n1046) );
  MUX21L U19801 ( .A(n4394), .B(n5182), .S(n4947), .Z(n1044) );
  MUX21L U19802 ( .A(n4928), .B(n2781), .S(n5279), .Z(n1041) );
  ND2 U19803 ( .A(n4928), .B(n4496), .Z(n2781) );
  MUX21L U19804 ( .A(n3367), .B(n3366), .S(n4605), .Z(n1023) );
  ND2 U19805 ( .A(n5258), .B(n4791), .Z(n3366) );
  ND2 U19806 ( .A(n4936), .B(n5258), .Z(n3367) );
  MUX21L U19807 ( .A(n3001), .B(n5236), .S(n4551), .Z(n1015) );
  ND2 U19808 ( .A(n5236), .B(n4811), .Z(n3001) );
  MUX21L U19809 ( .A(n5106), .B(n3368), .S(n4604), .Z(n992) );
  ND2 U19810 ( .A(n4791), .B(n5106), .Z(n3368) );
  MUX21L U19811 ( .A(n5124), .B(n4775), .S(n4573), .Z(n994) );
  MUX21L U19812 ( .A(n3269), .B(n4483), .S(n5253), .Z(n990) );
  ND2 U19813 ( .A(n4951), .B(n4483), .Z(n3269) );
  MUX21L U19814 ( .A(n4588), .B(n4836), .S(n5232), .Z(n989) );
  MUX21L U19815 ( .A(n2465), .B(n2464), .S(n4617), .Z(n943) );
  ND2 U19816 ( .A(n4762), .B(n5137), .Z(n2464) );
  ND2 U19817 ( .A(n5267), .B(n4916), .Z(n2465) );
  MUX21L U19818 ( .A(n5177), .B(n3002), .S(n4551), .Z(n955) );
  ND2 U19819 ( .A(n4945), .B(n5178), .Z(n3002) );
  MUX21L U19820 ( .A(n4744), .B(n2782), .S(n5279), .Z(n951) );
  ND2 U19821 ( .A(n4561), .B(n4744), .Z(n2782) );
  MUX21L U19822 ( .A(n3370), .B(n3369), .S(n4936), .Z(n960) );
  ND2 U19823 ( .A(n4492), .B(n5107), .Z(n3369) );
  ND2 U19824 ( .A(n5258), .B(n4493), .Z(n3370) );
  MUX21L U19825 ( .A(n4743), .B(n2783), .S(n4561), .Z(n917) );
  ND2 U19826 ( .A(n4744), .B(n5195), .Z(n2783) );
  MUX21L U19827 ( .A(n2971), .B(n4393), .S(n4946), .Z(n888) );
  ND2 U19828 ( .A(n4394), .B(n5181), .Z(n2971) );
  MUX21L U19829 ( .A(n4572), .B(n3526), .S(n5246), .Z(n874) );
  ND2 U19830 ( .A(n4572), .B(n4777), .Z(n3526) );
  ND2 U19831 ( .A(n2252), .B(n2251), .Z(n1032) );
  ND2 U19832 ( .A(n4868), .B(n5156), .Z(n2252) );
  ND2 U19833 ( .A(n4594), .B(n4868), .Z(n2251) );
  ND2 U19834 ( .A(n4948), .B(n5071), .Z(n1052) );
  ND3 U19835 ( .A(n4832), .B(n5089), .C(n4437), .Z(n842) );
  ND3 U19836 ( .A(n4749), .B(n5198), .C(n4499), .Z(n1040) );
  ND3 U19837 ( .A(n4748), .B(n5198), .C(n4498), .Z(n885) );
  ND3 U19838 ( .A(n4831), .B(n5089), .C(n4438), .Z(n868) );
  ND2 U19839 ( .A(n4843), .B(n5077), .Z(n1081) );
  MUX41 U19840 ( .D0(n1991), .D1(n1976), .D2(n1982), .D3(n1967), .A(n4208), 
        .B(n4221), .Z(N133) );
  ND4 U19841 ( .A(n4162), .B(n4161), .C(n4160), .D(n4159), .Z(n1982) );
  MUX21L U19842 ( .A(n4156), .B(n4155), .S(n4258), .Z(n4161) );
  AO2 U19843 ( .A(n4152), .B(n4295), .C(n4151), .D(n4295), .Z(n4160) );
  MUX21L U19844 ( .A(n4153), .B(n4154), .S(n4258), .Z(n4162) );
  MUX21L U19845 ( .A(n4158), .B(n4157), .S(n4260), .Z(n4159) );
  AN3 U19846 ( .A(n4333), .B(n1979), .C(n4290), .Z(n4158) );
  ND2 U19847 ( .A(n2756), .B(n2755), .Z(n1977) );
  NR3 U19848 ( .A(n4334), .B(n4194), .C(n4295), .Z(n4153) );
  IVP U19849 ( .A(n1981), .Z(n4194) );
  AO7 U19850 ( .A(n4581), .B(n5094), .C(n3101), .Z(n1981) );
  ND2 U19851 ( .A(n5241), .B(n4939), .Z(n3101) );
  MUX41 U19852 ( .D0(n1486), .D1(n1468), .D2(n1477), .D3(n1461), .A(n4209), 
        .B(n4220), .Z(N186) );
  NR2 U19853 ( .A(n4335), .B(n362), .Z(n4152) );
  ND2 U19854 ( .A(n4808), .B(n5179), .Z(n2985) );
  MUX41 U19855 ( .D0(n2026), .D1(n2009), .D2(n2017), .D3(n2000), .A(n4208), 
        .B(n4221), .Z(N134) );
  NR2 U19856 ( .A(n4335), .B(n363), .Z(n4154) );
  AO6 U19857 ( .A(n4565), .B(n4736), .C(n2857), .Z(n2859) );
  ND4 U19858 ( .A(n4102), .B(n4101), .C(n4100), .D(n4099), .Z(n1468) );
  AO2 U19859 ( .A(n4092), .B(n4260), .C(n4091), .D(n1467), .Z(n4100) );
  MUX21L U19860 ( .A(n4098), .B(n4097), .S(n4258), .Z(n4099) );
  MUX21L U19861 ( .A(n4096), .B(n4095), .S(n4258), .Z(n4101) );
  ND3 U19862 ( .A(n2232), .B(n2231), .C(n2230), .Z(n1997) );
  AO7 U19863 ( .A(n4960), .B(n4537), .C(n5148), .Z(n1999) );
  AO7 U19864 ( .A(n4910), .B(n4450), .C(n5171), .Z(n1993) );
  ND2 U19865 ( .A(n5280), .B(n4742), .Z(n2011) );
  AO7 U19866 ( .A(n4932), .B(n4565), .C(n5283), .Z(n2013) );
  AO7 U19867 ( .A(n4930), .B(n4562), .C(n5280), .Z(n2012) );
  MUX21L U19868 ( .A(n2257), .B(n4471), .S(n4964), .Z(n1964) );
  MUX21L U19869 ( .A(n5159), .B(n4467), .S(n4965), .Z(n1963) );
  AO7 U19870 ( .A(n5274), .B(n4461), .C(n2157), .Z(n1962) );
  MUX41 U19871 ( .D0(n1958), .D1(n1944), .D2(n1949), .D3(n1935), .A(n4208), 
        .B(n4221), .Z(N132) );
  MUX41 U19872 ( .D0(n1452), .D1(n1435), .D2(n1443), .D3(n1426), .A(n4209), 
        .B(n4220), .Z(N185) );
  NR2 U19873 ( .A(n4294), .B(n4190), .Z(n4095) );
  IVP U19874 ( .A(n1463), .Z(n4190) );
  AO7 U19875 ( .A(n4916), .B(n4526), .C(n5137), .Z(n1463) );
  ND3 U19876 ( .A(n4539), .B(n5150), .C(n4961), .Z(n1424) );
  MUX21L U19877 ( .A(n4472), .B(n4869), .S(n5277), .Z(n1423) );
  MUX21L U19878 ( .A(n4599), .B(n2149), .S(n5274), .Z(n1421) );
  NR2 U19879 ( .A(n4559), .B(n4751), .Z(n1436) );
  NR2 U19880 ( .A(n5281), .B(n4739), .Z(n1438) );
  MUX21L U19881 ( .A(n4828), .B(n4583), .S(n5237), .Z(n1444) );
  ND2 U19882 ( .A(n5250), .B(n3212), .Z(n1445) );
  MUX21L U19883 ( .A(n4479), .B(n5251), .S(n4952), .Z(n1446) );
  ND2 U19884 ( .A(n4943), .B(n4554), .Z(n1948) );
  AO7 U19885 ( .A(n5253), .B(n4484), .C(n4842), .Z(n1952) );
  AO7 U19886 ( .A(n5247), .B(n4924), .C(n4417), .Z(n1956) );
  ND2 U19887 ( .A(n3174), .B(n3173), .Z(n1951) );
  AN3 U19888 ( .A(n4333), .B(n4289), .C(n1462), .Z(n4097) );
  MUX21L U19889 ( .A(n4958), .B(n5263), .S(n4634), .Z(n1462) );
  IVP U19890 ( .A(n5058), .Z(n5294) );
  IVP U19891 ( .A(n5058), .Z(n5292) );
  IVP U19892 ( .A(n5058), .Z(n5293) );
  NR3 U19893 ( .A(n364), .B(n4336), .C(n4291), .Z(n3886) );
  ND2 U19894 ( .A(n5238), .B(n4582), .Z(n3122) );
  NR3 U19895 ( .A(n366), .B(n4336), .C(n4291), .Z(n3885) );
  ND2 U19896 ( .A(n4566), .B(n4799), .Z(n2897) );
  NR3 U19897 ( .A(n367), .B(n4335), .C(n4264), .Z(n3882) );
  ND2 U19898 ( .A(n4552), .B(n4814), .Z(n3014) );
  MUX41 U19899 ( .D0(n1418), .D1(n1406), .D2(n1410), .D3(n1397), .A(n4209), 
        .B(n4220), .Z(N184) );
  AO7 U19900 ( .A(n5291), .B(n4517), .C(n4894), .Z(n1403) );
  ND2 U19901 ( .A(n2399), .B(n4977), .Z(n1399) );
  MUX21L U19902 ( .A(n2372), .B(n4532), .S(n5263), .Z(n1398) );
  ND2 U19903 ( .A(n4461), .B(n4861), .Z(n1392) );
  ND2 U19904 ( .A(n4593), .B(n5156), .Z(n1394) );
  AO7 U19905 ( .A(n4961), .B(n5148), .C(n4632), .Z(n1396) );
  AN3 U19906 ( .A(n1408), .B(n4251), .C(n4331), .Z(n3884) );
  MUX21L U19907 ( .A(n2826), .B(n5281), .S(n4930), .Z(n1408) );
  ND2 U19908 ( .A(n5281), .B(n4405), .Z(n2826) );
  AN3 U19909 ( .A(n1407), .B(n4251), .C(n4331), .Z(n3883) );
  MUX21L U19910 ( .A(n4750), .B(n2742), .S(n5278), .Z(n1407) );
  ND2 U19911 ( .A(n4559), .B(n4751), .Z(n2742) );
  ND3 U19912 ( .A(n3889), .B(n3888), .C(n3887), .Z(n1410) );
  MUX21L U19913 ( .A(n3881), .B(n3882), .S(n4292), .Z(n3889) );
  MUX21L U19914 ( .A(n3884), .B(n3883), .S(n4291), .Z(n3887) );
  MUX21L U19915 ( .A(n3886), .B(n3885), .S(n4264), .Z(n3888) );
  MUX41 U19916 ( .D0(n1926), .D1(n1908), .D2(n1917), .D3(n1899), .A(n4210), 
        .B(n4221), .Z(N131) );
  IVP U19917 ( .A(n5058), .Z(n5295) );
  NR2 U19918 ( .A(n4339), .B(n4292), .Z(n4091) );
  NR2 U19919 ( .A(n4339), .B(n4294), .Z(n4092) );
  AO4 U19920 ( .A(n4955), .B(n4585), .C(n5233), .D(n4956), .Z(n1919) );
  ND2 U19921 ( .A(n3285), .B(n3284), .Z(n1921) );
  MUX21L U19922 ( .A(n5247), .B(n4776), .S(n4572), .Z(n1924) );
  ND3 U19923 ( .A(n4912), .B(n4458), .C(n5273), .Z(n1893) );
  MUX21L U19924 ( .A(n5150), .B(n4631), .S(n4961), .Z(n1898) );
  MUX21L U19925 ( .A(n4629), .B(n2268), .S(n4963), .Z(n1897) );
  AN3 U19926 ( .A(n4289), .B(n1464), .C(n4333), .Z(n4098) );
  ND2 U19927 ( .A(n4522), .B(n5214), .Z(n1464) );
  IVP U19928 ( .A(n5058), .Z(n5291) );
  MUX41 U19929 ( .D0(n1388), .D1(n1372), .D2(n1381), .D3(n1363), .A(n4209), 
        .B(n4219), .Z(N183) );
  NR2 U19930 ( .A(n4917), .B(n4475), .Z(n1367) );
  AO7 U19931 ( .A(n4621), .B(n5215), .C(n4888), .Z(n1368) );
  ND3 U19932 ( .A(n4906), .B(n4509), .C(n5294), .Z(n1370) );
  AN3 U19933 ( .A(n1382), .B(n4332), .C(n4251), .Z(n3986) );
  ND2 U19934 ( .A(n3144), .B(n3143), .Z(n1382) );
  ND2 U19935 ( .A(n3140), .B(n4828), .Z(n3143) );
  MUX21L U19936 ( .A(n3141), .B(n3142), .S(n4583), .Z(n3144) );
  EO U19937 ( .A(n5227), .B(n4927), .Z(n782) );
  MUX41 U19938 ( .D0(n1890), .D1(n1872), .D2(n1881), .D3(n1865), .A(n4210), 
        .B(n4221), .Z(N130) );
  ND4 U19939 ( .A(n4114), .B(n4113), .C(n4112), .D(n4111), .Z(n1872) );
  MUX21L U19940 ( .A(n4105), .B(n4106), .S(n4258), .Z(n4114) );
  AO2 U19941 ( .A(n4104), .B(n4338), .C(n4103), .D(n1871), .Z(n4112) );
  MUX21L U19942 ( .A(n4107), .B(n4108), .S(n4294), .Z(n4113) );
  NR2 U19943 ( .A(n4965), .B(n4470), .Z(n1360) );
  NR2 U19944 ( .A(n4913), .B(n4599), .Z(n1358) );
  AO7 U19945 ( .A(n5261), .B(n4875), .C(n4632), .Z(n1362) );
  MUX21L U19946 ( .A(n4110), .B(n4109), .S(n4260), .Z(n4111) );
  AN3 U19947 ( .A(n1866), .B(n4289), .C(n4333), .Z(n4109) );
  MUX21L U19948 ( .A(n4532), .B(n5144), .S(n4978), .Z(n1866) );
  MUX41 U19949 ( .D0(n1354), .D1(n1338), .D2(n1346), .D3(n1329), .A(n4209), 
        .B(n4219), .Z(N182) );
  ND2 U19950 ( .A(n4567), .B(n4797), .Z(n1876) );
  ND2 U19951 ( .A(n2926), .B(n2925), .Z(n1877) );
  MUX21L U19952 ( .A(n5095), .B(n3082), .S(n4941), .Z(n1880) );
  AN3 U19953 ( .A(n1324), .B(n4253), .C(n4288), .Z(n3666) );
  ND2 U19954 ( .A(n2080), .B(n2079), .Z(n1324) );
  ND2 U19955 ( .A(n5271), .B(n4626), .Z(n2079) );
  EN U19956 ( .A(n5228), .B(n4910), .Z(n2080) );
  NR3 U19957 ( .A(n4294), .B(n4337), .C(n368), .Z(n4106) );
  ND2 U19958 ( .A(n5288), .B(n4477), .Z(n2518) );
  ND2 U19959 ( .A(n4618), .B(n4761), .Z(n1868) );
  NR2 U19960 ( .A(n4294), .B(n4260), .Z(n4103) );
  NR2 U19961 ( .A(n4294), .B(n4258), .Z(n4104) );
  ND2 U19962 ( .A(n4950), .B(n4485), .Z(n1349) );
  AO7 U19963 ( .A(n5236), .B(n4958), .C(n4583), .Z(n1347) );
  ND3 U19964 ( .A(n4802), .B(n5133), .C(n4579), .Z(n1353) );
  NR3 U19965 ( .A(n4637), .B(n5265), .C(n4976), .Z(n1331) );
  ND3 U19966 ( .A(n4592), .B(n5220), .C(n4903), .Z(n1333) );
  MUX21L U19967 ( .A(n5146), .B(n2359), .S(n4958), .Z(n1330) );
  NR3 U19968 ( .A(n4187), .B(n4297), .C(n4268), .Z(n3665) );
  IVP U19969 ( .A(n1328), .Z(n4187) );
  AO7 U19970 ( .A(n5260), .B(n4961), .C(n4539), .Z(n1328) );
  MUX41 U19971 ( .D0(n1856), .D1(n1838), .D2(n1847), .D3(n1830), .A(n4210), 
        .B(n4221), .Z(N129) );
  MUX41 U19972 ( .D0(n1323), .D1(n1308), .D2(n1317), .D3(n1300), .A(n4209), 
        .B(n4219), .Z(N181) );
  ND4 U19973 ( .A(n4047), .B(n4046), .C(n4045), .D(n4044), .Z(n1300) );
  MUX21L U19974 ( .A(n4042), .B(n4043), .S(n4259), .Z(n4044) );
  MUX21L U19975 ( .A(n4038), .B(n4039), .S(n4260), .Z(n4046) );
  MUX21L U19976 ( .A(n4036), .B(n4037), .S(n4341), .Z(n4047) );
  AO7 U19977 ( .A(n5273), .B(n4913), .C(n4458), .Z(n1824) );
  MUX21L U19978 ( .A(n4593), .B(n2256), .S(n4964), .Z(n1827) );
  MUX21L U19979 ( .A(n4913), .B(n5273), .S(n4600), .Z(n1825) );
  MUX21L U19980 ( .A(n5102), .B(n4814), .S(n4553), .Z(n1844) );
  MUX21L U19981 ( .A(n4804), .B(n2927), .S(n4549), .Z(n1843) );
  MUX21L U19982 ( .A(n2861), .B(n2860), .S(n4932), .Z(n1842) );
  NR3 U19983 ( .A(n370), .B(n4294), .C(n4259), .Z(n4036) );
  NR2 U19984 ( .A(n2327), .B(n2326), .Z(n2329) );
  ND2 U19985 ( .A(n3418), .B(n3417), .Z(n1321) );
  MUX21L U19986 ( .A(n5255), .B(n4949), .S(n4609), .Z(n1320) );
  MUX21L U19987 ( .A(n3264), .B(n5077), .S(n4951), .Z(n1319) );
  AN3 U19988 ( .A(n1301), .B(n4331), .C(n4252), .Z(n3770) );
  MUX21L U19989 ( .A(n2360), .B(n4958), .S(n4634), .Z(n1301) );
  ND2 U19990 ( .A(n5263), .B(n4958), .Z(n2360) );
  ND2 U19991 ( .A(n2083), .B(n2082), .Z(n1295) );
  ND2 U19992 ( .A(n4910), .B(n4626), .Z(n2082) );
  MUX21L U19993 ( .A(n2081), .B(n4626), .S(n5271), .Z(n2083) );
  ND2 U19994 ( .A(n2128), .B(n2127), .Z(n1296) );
  ND2 U19995 ( .A(n5273), .B(n4600), .Z(n2127) );
  EO U19996 ( .A(n4900), .B(n4600), .Z(n2128) );
  MUX41 U19997 ( .D0(n1822), .D1(n1806), .D2(n1814), .D3(n1797), .A(n4209), 
        .B(n4220), .Z(N128) );
  NR2 U19998 ( .A(n4558), .B(n5202), .Z(n1807) );
  AO7 U19999 ( .A(n5280), .B(n4562), .C(n4742), .Z(n1808) );
  MUX41 U20000 ( .D0(n1294), .D1(n1277), .D2(n1285), .D3(n1273), .A(n4209), 
        .B(n4219), .Z(N180) );
  ND4 U20001 ( .A(n4090), .B(n4089), .C(n4088), .D(n4087), .Z(n1277) );
  AO2 U20002 ( .A(n4080), .B(n4294), .C(n4079), .D(n4294), .Z(n4088) );
  MUX21L U20003 ( .A(n4081), .B(n4082), .S(n4258), .Z(n4090) );
  MUX21L U20004 ( .A(n4084), .B(n4083), .S(n4258), .Z(n4089) );
  NR2 U20005 ( .A(n4963), .B(n4628), .Z(n1790) );
  AN3 U20006 ( .A(n4900), .B(n4546), .C(n5222), .Z(n1795) );
  ND2 U20007 ( .A(n2072), .B(n2071), .Z(n1791) );
  NR2 U20008 ( .A(n5235), .B(n4389), .Z(n1282) );
  NR2 U20009 ( .A(n5239), .B(n4823), .Z(n1284) );
  NR2 U20010 ( .A(n4905), .B(n4559), .Z(n1278) );
  MUX21L U20011 ( .A(n4086), .B(n4085), .S(n4258), .Z(n4087) );
  AN3 U20012 ( .A(n4333), .B(n1275), .C(n4289), .Z(n4086) );
  ND2 U20013 ( .A(n4973), .B(n4634), .Z(n1274) );
  MUX41 U20014 ( .D0(n1789), .D1(n1771), .D2(n1780), .D3(n1763), .A(n4210), 
        .B(n4220), .Z(N127) );
  NR2 U20015 ( .A(n4340), .B(n372), .Z(n4082) );
  EN U20016 ( .A(n5225), .B(n4976), .Z(n2520) );
  ND4 U20017 ( .A(n4035), .B(n4034), .C(n4033), .D(n4032), .Z(n1763) );
  MUX21L U20018 ( .A(n4024), .B(n4025), .S(n4293), .Z(n4035) );
  MUX21L U20019 ( .A(n4027), .B(n4026), .S(n4260), .Z(n4034) );
  MUX21L U20020 ( .A(n4030), .B(n4031), .S(n4262), .Z(n4032) );
  ND2 U20021 ( .A(n2247), .B(n2246), .Z(n1270) );
  MUX21L U20022 ( .A(n2317), .B(n4960), .S(n4632), .Z(n1272) );
  MUX21L U20023 ( .A(n5173), .B(n2055), .S(n4627), .Z(n1266) );
  NR3 U20024 ( .A(n4340), .B(n2713), .C(n4294), .Z(n4081) );
  ND2 U20025 ( .A(n4907), .B(n4557), .Z(n2713) );
  ND2 U20026 ( .A(n2198), .B(n2197), .Z(n1760) );
  ND2 U20027 ( .A(n4596), .B(n4864), .Z(n2197) );
  EO U20028 ( .A(n5230), .B(n4596), .Z(n2198) );
  ND2 U20029 ( .A(n2087), .B(n2086), .Z(n1759) );
  ND2 U20030 ( .A(n4602), .B(n4854), .Z(n2086) );
  MUX21L U20031 ( .A(n5271), .B(n2085), .S(n4910), .Z(n2087) );
  NR2 U20032 ( .A(n4340), .B(n5295), .Z(n4080) );
  MUX41 U20033 ( .D0(n1265), .D1(n1250), .D2(n1257), .D3(n1245), .A(n4209), 
        .B(n4219), .Z(N179) );
  NR3 U20034 ( .A(n4293), .B(n4340), .C(n371), .Z(n4026) );
  NR2 U20035 ( .A(n2160), .B(n2159), .Z(n2162) );
  ND4 U20036 ( .A(n4150), .B(n4149), .C(n4148), .D(n4147), .Z(n1257) );
  MUX21L U20037 ( .A(n4139), .B(n4140), .S(n4336), .Z(n4150) );
  MUX21L U20038 ( .A(n4141), .B(n4142), .S(n4259), .Z(n4149) );
  MUX21L U20039 ( .A(n4145), .B(n4146), .S(n4258), .Z(n4147) );
  MUX21L U20040 ( .A(n3222), .B(n3221), .S(n4953), .Z(n1783) );
  MUX21L U20041 ( .A(n5123), .B(n4776), .S(n4572), .Z(n1787) );
  MUX21L U20042 ( .A(n5088), .B(n4955), .S(n4585), .Z(n1782) );
  NR2 U20043 ( .A(n4293), .B(n4189), .Z(n4027) );
  IVP U20044 ( .A(n1762), .Z(n4189) );
  AO7 U20045 ( .A(n5262), .B(n4877), .C(n2351), .Z(n1762) );
  ND2 U20046 ( .A(n4959), .B(n4633), .Z(n2351) );
  EN U20047 ( .A(n5230), .B(n4564), .Z(n1252) );
  MUX21L U20048 ( .A(n4122), .B(n4121), .S(n4259), .Z(n4123) );
  AN3 U20049 ( .A(n4290), .B(n1249), .C(n4334), .Z(n4122) );
  AN3 U20050 ( .A(n4334), .B(n4290), .C(n1246), .Z(n4121) );
  ND2 U20051 ( .A(n2572), .B(n2571), .Z(n1249) );
  MUX41 U20052 ( .D0(n1757), .D1(n1740), .D2(n1748), .D3(n1732), .A(n4208), 
        .B(n4220), .Z(N126) );
  EN U20053 ( .A(n5227), .B(n4973), .Z(n783) );
  NR2 U20054 ( .A(n4294), .B(n373), .Z(n4120) );
  ND2 U20055 ( .A(n4624), .B(n4896), .Z(n2654) );
  MUX21L U20056 ( .A(n4594), .B(n2248), .S(n5276), .Z(n1242) );
  MUX21L U20057 ( .A(n5172), .B(n2056), .S(n4909), .Z(n1238) );
  ND2 U20058 ( .A(n2320), .B(n2319), .Z(n1244) );
  MUX21L U20059 ( .A(n4928), .B(n2775), .S(n5279), .Z(n1251) );
  ND2 U20060 ( .A(n4928), .B(n4496), .Z(n2775) );
  NR3 U20061 ( .A(n374), .B(n4295), .C(n4259), .Z(n4139) );
  ND2 U20062 ( .A(n5240), .B(n4823), .Z(n3092) );
  EN U20063 ( .A(n4899), .B(n4631), .Z(n784) );
  NR2 U20064 ( .A(n4337), .B(n4294), .Z(n4115) );
  NR2 U20065 ( .A(n4337), .B(n4294), .Z(n4116) );
  MUX41 U20066 ( .D0(n1237), .D1(n1223), .D2(n1229), .D3(n1216), .A(n4209), 
        .B(n4219), .Z(N178) );
  ND4 U20067 ( .A(n4174), .B(n4173), .C(n4172), .D(n4171), .Z(n1229) );
  MUX21L U20068 ( .A(n4163), .B(n4164), .S(n4335), .Z(n4174) );
  MUX21L U20069 ( .A(n4165), .B(n4166), .S(n4260), .Z(n4173) );
  MUX21L U20070 ( .A(n4170), .B(n4169), .S(n4295), .Z(n4171) );
  ND2 U20071 ( .A(n5234), .B(n4820), .Z(n1746) );
  MUX21L U20072 ( .A(n5278), .B(n4559), .S(n4906), .Z(n1741) );
  AN3 U20073 ( .A(n1727), .B(n4289), .C(n4252), .Z(n3732) );
  ND3 U20074 ( .A(n2047), .B(n2046), .C(n2045), .Z(n1727) );
  ND2 U20075 ( .A(n4446), .B(n4857), .Z(n2046) );
  ND2 U20076 ( .A(n5270), .B(n4858), .Z(n2047) );
  NR3 U20077 ( .A(n4259), .B(n4295), .C(n4195), .Z(n4163) );
  IVP U20078 ( .A(n1228), .Z(n4195) );
  AO7 U20079 ( .A(n4939), .B(n4377), .C(n3110), .Z(n1228) );
  ND2 U20080 ( .A(n5240), .B(n4582), .Z(n3110) );
  NR3 U20081 ( .A(n375), .B(n4334), .C(n4295), .Z(n4166) );
  ND2 U20082 ( .A(n4801), .B(n5188), .Z(n2883) );
  ND2 U20083 ( .A(n2656), .B(n2655), .Z(n1222) );
  AO7 U20084 ( .A(n4635), .B(n4881), .C(n2379), .Z(n1217) );
  ND2 U20085 ( .A(n2477), .B(n2476), .Z(n1218) );
  MUX21L U20086 ( .A(n4867), .B(n2249), .S(n4594), .Z(n1213) );
  ND2 U20087 ( .A(n2146), .B(n2145), .Z(n1211) );
  MUX21L U20088 ( .A(n4960), .B(n2321), .S(n5261), .Z(n1215) );
  AN3 U20089 ( .A(n4253), .B(n1225), .C(n4333), .Z(n4170) );
  ND2 U20090 ( .A(n2831), .B(n2830), .Z(n1225) );
  ND2 U20091 ( .A(n4563), .B(n4738), .Z(n2830) );
  MUX21L U20092 ( .A(n5281), .B(n2829), .S(n4930), .Z(n2831) );
  MUX41 U20093 ( .D0(n1726), .D1(n1710), .D2(n1718), .D3(n1702), .A(n4209), 
        .B(n4220), .Z(N125) );
  ND2 U20094 ( .A(n4954), .B(n5084), .Z(n1719) );
  MUX21L U20095 ( .A(n3407), .B(n4938), .S(n4588), .Z(n1723) );
  MUX21L U20096 ( .A(n4610), .B(n3287), .S(n4950), .Z(n1721) );
  AN3 U20097 ( .A(n5070), .B(n4289), .C(n4252), .Z(n3733) );
  ND2 U20098 ( .A(n4943), .B(n4387), .Z(n1226) );
  MUX21L U20099 ( .A(n5157), .B(n2240), .S(n4595), .Z(n1700) );
  ND2 U20100 ( .A(n2126), .B(n2125), .Z(n1697) );
  EO U20101 ( .A(n5227), .B(n4908), .Z(n1696) );
  MUX41 U20102 ( .D0(n1208), .D1(n1194), .D2(n1201), .D3(n1186), .A(n4210), 
        .B(n4219), .Z(N177) );
  NR3 U20103 ( .A(n378), .B(n4297), .C(n4268), .Z(n3675) );
  ND2 U20104 ( .A(n5260), .B(n4630), .Z(n2302) );
  MUX41 U20105 ( .D0(n1695), .D1(n1681), .D2(n1689), .D3(n1674), .A(LogIn2[47]), .B(n4220), .Z(N124) );
  NR2 U20106 ( .A(n4918), .B(n4429), .Z(n1205) );
  MUX21L U20107 ( .A(n4421), .B(n4921), .S(n5246), .Z(n1206) );
  ND2 U20108 ( .A(n3171), .B(n4438), .Z(n1202) );
  ND3 U20109 ( .A(n2493), .B(n2492), .C(n2491), .Z(n1190) );
  EO U20110 ( .A(n4898), .B(n4637), .Z(n1188) );
  MUX21L U20111 ( .A(n4891), .B(n2605), .S(n4622), .Z(n1192) );
  NR3 U20112 ( .A(n376), .B(n4292), .C(n4263), .Z(n3913) );
  ND2 U20113 ( .A(n4780), .B(n5118), .Z(n3486) );
  ND2 U20114 ( .A(n4499), .B(n4749), .Z(n1682) );
  MUX21L U20115 ( .A(n4819), .B(n5098), .S(n4556), .Z(n1688) );
  ND2 U20116 ( .A(n4947), .B(n2960), .Z(n1686) );
  AN3 U20117 ( .A(n1690), .B(n4251), .C(n4288), .Z(n3914) );
  NR2 U20118 ( .A(n4955), .B(n4585), .Z(n1690) );
  MUX41 U20119 ( .D0(n1181), .D1(n1166), .D2(n1173), .D3(n1160), .A(n4210), 
        .B(n4219), .Z(N176) );
  OR3 U20120 ( .A(n4627), .B(n5270), .C(n4909), .Z(n785) );
  NR2 U20121 ( .A(n4351), .B(n4188), .Z(n3685) );
  IVP U20122 ( .A(n1159), .Z(n4188) );
  AO4 U20123 ( .A(n4960), .B(n4632), .C(n5261), .D(n4632), .Z(n1159) );
  MUX41 U20124 ( .D0(n1666), .D1(n1648), .D2(n1657), .D3(n1640), .A(n4208), 
        .B(n4220), .Z(N123) );
  MUX21L U20125 ( .A(n4745), .B(n2777), .S(n4560), .Z(n1167) );
  EO U20126 ( .A(n5228), .B(n4947), .Z(n1169) );
  ND3 U20127 ( .A(n2834), .B(n2833), .C(n2832), .Z(n1168) );
  NR2 U20128 ( .A(n5257), .B(n4935), .Z(n1177) );
  NR3 U20129 ( .A(n4613), .B(n5252), .C(n4952), .Z(n1175) );
  AO7 U20130 ( .A(n4575), .B(n4772), .C(n5248), .Z(n1180) );
  ND3 U20131 ( .A(n3692), .B(n3691), .C(n3690), .Z(n1160) );
  MUX21L U20132 ( .A(n3688), .B(n3689), .S(n4351), .Z(n3691) );
  MUX21L U20133 ( .A(n3685), .B(n3684), .S(n4267), .Z(n3690) );
  MUX21L U20134 ( .A(n3686), .B(n3687), .S(n4297), .Z(n3692) );
  ND2 U20135 ( .A(n2304), .B(n2303), .Z(n1158) );
  ND2 U20136 ( .A(n5260), .B(n4631), .Z(n2304) );
  ND2 U20137 ( .A(n4962), .B(n4631), .Z(n2303) );
  NR3 U20138 ( .A(n380), .B(n4297), .C(n4268), .Z(n3637) );
  ND2 U20139 ( .A(n4963), .B(n4541), .Z(n2275) );
  ND2 U20140 ( .A(n2916), .B(n4397), .Z(n1652) );
  ND2 U20141 ( .A(n2991), .B(n2990), .Z(n1654) );
  ND2 U20142 ( .A(n2820), .B(n2819), .Z(n1651) );
  AN3 U20143 ( .A(n1182), .B(n4252), .C(n4288), .Z(n3676) );
  ND3 U20144 ( .A(n4854), .B(n5170), .C(n4454), .Z(n1182) );
  NR3 U20145 ( .A(n381), .B(n4350), .C(n4297), .Z(n3641) );
  ND2 U20146 ( .A(n4874), .B(n5149), .Z(n2313) );
  MUX41 U20147 ( .D0(n1157), .D1(n1143), .D2(n1149), .D3(n1138), .A(n4210), 
        .B(n4219), .Z(N175) );
  ND2 U20148 ( .A(n3696), .B(n3695), .Z(n1138) );
  NR2 U20149 ( .A(n4297), .B(n4409), .Z(n3684) );
  OR3 U20150 ( .A(n4625), .B(n5292), .C(n4970), .Z(n786) );
  ND2 U20151 ( .A(n4425), .B(n5116), .Z(n1154) );
  ND2 U20152 ( .A(n5259), .B(n4433), .Z(n1153) );
  ND2 U20153 ( .A(n5246), .B(n4921), .Z(n1155) );
  MUX41 U20154 ( .D0(n1634), .D1(n1616), .D2(n1625), .D3(n1608), .A(n4208), 
        .B(n4220), .Z(N122) );
  ND4 U20155 ( .A(n3655), .B(n3654), .C(n3653), .D(n3652), .Z(n1608) );
  NR3 U20156 ( .A(n4193), .B(n4336), .C(n4291), .Z(n3854) );
  IVP U20157 ( .A(n1148), .Z(n4193) );
  AO7 U20158 ( .A(n5240), .B(n4379), .C(n4940), .Z(n1148) );
  ND2 U20159 ( .A(n2739), .B(n2738), .Z(n1617) );
  MUX21L U20160 ( .A(n2866), .B(n5283), .S(n4565), .Z(n1620) );
  ND2 U20161 ( .A(n2822), .B(n2821), .Z(n1619) );
  AO7 U20162 ( .A(n4574), .B(n5127), .C(n4924), .Z(n1633) );
  MUX21L U20163 ( .A(n4427), .B(n4782), .S(n5244), .Z(n1631) );
  MUX21L U20164 ( .A(n5088), .B(n4586), .S(n4955), .Z(n1627) );
  NR2 U20165 ( .A(n4978), .B(n4634), .Z(n1139) );
  MUX41 U20166 ( .D0(n1136), .D1(n1123), .D2(n1127), .D3(n1121), .A(n4210), 
        .B(n4219), .Z(N174) );
  ND2 U20167 ( .A(n3698), .B(n3697), .Z(n1121) );
  AN3 U20168 ( .A(n1144), .B(n4251), .C(n4289), .Z(n3851) );
  ND2 U20169 ( .A(n4408), .B(n4741), .Z(n1144) );
  MUX41 U20170 ( .D0(n1603), .D1(n1586), .D2(n1595), .D3(n1580), .A(n4209), 
        .B(n4220), .Z(N121) );
  ND2 U20171 ( .A(n3661), .B(n3660), .Z(n1580) );
  ND4 U20172 ( .A(n4078), .B(n4077), .C(n4076), .D(n4075), .Z(n1586) );
  MUX21L U20173 ( .A(n4067), .B(n4068), .S(n4337), .Z(n4078) );
  MUX21L U20174 ( .A(n4071), .B(n4072), .S(n4341), .Z(n4076) );
  MUX21L U20175 ( .A(n4069), .B(n4070), .S(n4259), .Z(n4077) );
  AO7 U20176 ( .A(n5244), .B(n4782), .C(n4426), .Z(n1133) );
  ND2 U20177 ( .A(n3155), .B(n3154), .Z(n1128) );
  MUX21L U20178 ( .A(n3572), .B(n3571), .S(n4925), .Z(n1135) );
  AN3 U20179 ( .A(n1125), .B(n4331), .C(n4288), .Z(n3863) );
  AO7 U20180 ( .A(n5286), .B(n4947), .C(n4549), .Z(n1125) );
  ND2 U20181 ( .A(n3813), .B(n3812), .Z(n1123) );
  EO U20182 ( .A(n4290), .B(n4265), .Z(n3812) );
  MUX21L U20183 ( .A(n3811), .B(n3810), .S(n4265), .Z(n3813) );
  NR2 U20184 ( .A(n4353), .B(n760), .Z(n3811) );
  ND2 U20185 ( .A(n2741), .B(n2740), .Z(n1587) );
  MUX21L U20186 ( .A(n4747), .B(n2769), .S(n4560), .Z(n1588) );
  ND2 U20187 ( .A(n2854), .B(n2853), .Z(n1589) );
  NR2 U20188 ( .A(n4975), .B(n4619), .Z(n1584) );
  IVP U20189 ( .A(n1119), .Z(n4198) );
  ND2 U20190 ( .A(n3219), .B(n4478), .Z(n1112) );
  MUX21L U20191 ( .A(n5125), .B(n4417), .S(n4923), .Z(n1117) );
  MUX21L U20192 ( .A(n3749), .B(n3748), .S(n4208), .Z(n3751) );
  NR2 U20193 ( .A(n4222), .B(n384), .Z(n3748) );
  NR2 U20194 ( .A(n4222), .B(n4198), .Z(n3749) );
  ND2 U20195 ( .A(n2424), .B(n2423), .Z(n1581) );
  ND2 U20196 ( .A(n5266), .B(n4615), .Z(n2424) );
  ND2 U20197 ( .A(n4914), .B(n4615), .Z(n2423) );
  NR3 U20198 ( .A(n4573), .B(n4294), .C(n4261), .Z(n4067) );
  NR3 U20199 ( .A(n4637), .B(n4335), .C(n4264), .Z(n3859) );
  MUX21L U20200 ( .A(n3658), .B(n3659), .S(n4268), .Z(n3660) );
  NR3 U20201 ( .A(n4297), .B(n4351), .C(n4186), .Z(n3659) );
  ND3 U20202 ( .A(n4870), .B(n5154), .C(n4542), .Z(n1579) );
  MUX21L U20203 ( .A(n3870), .B(n3869), .S(n4291), .Z(n3874) );
  NR2 U20204 ( .A(n4335), .B(n2661), .Z(n3870) );
  NR2 U20205 ( .A(n4264), .B(n385), .Z(n3869) );
  MUX41 U20206 ( .D0(n1577), .D1(n1560), .D2(n1569), .D3(n1558), .A(n4209), 
        .B(n4220), .Z(N120) );
  AO7 U20207 ( .A(n764), .B(n3663), .C(n3662), .Z(n1558) );
  NR2 U20208 ( .A(n5248), .B(n4924), .Z(n1576) );
  ND2 U20209 ( .A(n4955), .B(n4586), .Z(n1571) );
  MUX21L U20210 ( .A(n5104), .B(n3340), .S(n4606), .Z(n1573) );
  ND3 U20211 ( .A(n3784), .B(n3783), .C(n3782), .Z(n1560) );
  MUX21L U20212 ( .A(n3777), .B(n4296), .S(n4353), .Z(n3783) );
  MUX21L U20213 ( .A(n3779), .B(n3778), .S(n4295), .Z(n3784) );
  MUX21L U20214 ( .A(n3780), .B(n3781), .S(n4295), .Z(n3782) );
  ND2 U20215 ( .A(n2426), .B(n2425), .Z(n1559) );
  ND2 U20216 ( .A(n5266), .B(n4615), .Z(n2426) );
  ND2 U20217 ( .A(n4914), .B(n4615), .Z(n2425) );
  OR3 U20218 ( .A(n4624), .B(n5292), .C(n4971), .Z(n787) );
  NR2 U20219 ( .A(n4353), .B(n760), .Z(n3779) );
  NR2 U20220 ( .A(n4291), .B(n4264), .Z(n3871) );
  AN3 U20221 ( .A(n1103), .B(n4250), .C(n4288), .Z(n3958) );
  AO4 U20222 ( .A(n4955), .B(n4586), .C(n5232), .D(n4586), .Z(n1103) );
  ND2 U20223 ( .A(n4062), .B(n4061), .Z(N119) );
  AO2 U20224 ( .A(n4222), .B(n1548), .C(n4222), .D(n4208), .Z(n4062) );
  MUX21L U20225 ( .A(n4060), .B(n1542), .S(n4208), .Z(n4061) );
  NR3 U20226 ( .A(n3514), .B(n4292), .C(n4262), .Z(n3957) );
  ND3 U20227 ( .A(n4571), .B(n5121), .C(n4922), .Z(n3514) );
  MUX21L U20228 ( .A(n3969), .B(n3968), .S(n4292), .Z(n3974) );
  NR2 U20229 ( .A(n4339), .B(n387), .Z(n3969) );
  NR3 U20230 ( .A(n4339), .B(n761), .C(n4262), .Z(n3968) );
  NR2 U20231 ( .A(n4222), .B(n4200), .Z(n4060) );
  IVP U20232 ( .A(n1557), .Z(n4200) );
  MUX21L U20233 ( .A(n4951), .B(n4482), .S(n5253), .Z(n1551) );
  NR2 U20234 ( .A(n4295), .B(n4266), .Z(n3777) );
  NR3 U20235 ( .A(n4193), .B(n4335), .C(n4290), .Z(n3832) );
  NR2 U20236 ( .A(n4266), .B(n4443), .Z(n3778) );
  NR2 U20237 ( .A(n4293), .B(n4185), .Z(n3967) );
  IVP U20238 ( .A(n1098), .Z(n4185) );
  AO4 U20239 ( .A(n4952), .B(n4612), .C(n5252), .D(n4612), .Z(n1098) );
  NR3 U20240 ( .A(n386), .B(n4290), .C(n4265), .Z(n3828) );
  ND2 U20241 ( .A(n4817), .B(n5100), .Z(n3044) );
  ND2 U20242 ( .A(n2428), .B(n2427), .Z(n1541) );
  ND2 U20243 ( .A(n5266), .B(n4615), .Z(n2428) );
  ND2 U20244 ( .A(n4914), .B(n4615), .Z(n2427) );
  NR2 U20245 ( .A(n4221), .B(n4199), .Z(n3741) );
  IVP U20246 ( .A(n1540), .Z(n4199) );
  AO7 U20247 ( .A(n5232), .B(n4436), .C(n4955), .Z(n1533) );
  AN3 U20248 ( .A(n4288), .B(n1099), .C(n4332), .Z(n3970) );
  NR2 U20249 ( .A(n4936), .B(n4605), .Z(n1099) );
  OR3 U20250 ( .A(n4551), .B(n5234), .C(n4945), .Z(n788) );
  NR2 U20251 ( .A(n4353), .B(n4579), .Z(n3786) );
  OR3 U20252 ( .A(n4563), .B(n5281), .C(n4930), .Z(n789) );
  AN3 U20253 ( .A(n4289), .B(n1529), .C(n4331), .Z(n3841) );
  ND2 U20254 ( .A(n2979), .B(n4392), .Z(n1529) );
  ND2 U20255 ( .A(n5233), .B(n4946), .Z(n2979) );
  ND3 U20256 ( .A(n3845), .B(n3844), .C(n3843), .Z(n1531) );
  MUX21L U20257 ( .A(n3837), .B(n3838), .S(n4265), .Z(n3844) );
  MUX21L U20258 ( .A(n3841), .B(n3842), .S(n4265), .Z(n3843) );
  MUX21L U20259 ( .A(n3840), .B(n3839), .S(n4290), .Z(n3845) );
  NR2 U20260 ( .A(n4334), .B(n4567), .Z(n3840) );
  NR2 U20261 ( .A(n4221), .B(n4201), .Z(n3740) );
  IVP U20262 ( .A(n1528), .Z(n4201) );
  AO3 U20263 ( .A(n4352), .B(n4186), .C(n4267), .D(n4296), .Z(n1528) );
  NR2 U20264 ( .A(n4339), .B(n4293), .Z(n3971) );
  NR2 U20265 ( .A(n4340), .B(n4186), .Z(n4012) );
  MUX21L U20266 ( .A(n4922), .B(n3518), .S(n5246), .Z(n1095) );
  ND2 U20267 ( .A(n4922), .B(n4420), .Z(n3518) );
  NR2 U20268 ( .A(n4335), .B(n4290), .Z(n3842) );
  NR2 U20269 ( .A(n4261), .B(n390), .Z(n3976) );
  ND2 U20270 ( .A(n4576), .B(n4771), .Z(n3580) );
  AO7 U20271 ( .A(n4590), .B(n4784), .C(n5113), .Z(n1524) );
  AO7 U20272 ( .A(n5257), .B(n4794), .C(n4606), .Z(n1523) );
  NR3 U20273 ( .A(n4583), .B(n5237), .C(n4953), .Z(n1520) );
  ND2 U20274 ( .A(n3903), .B(n3902), .Z(n1519) );
  NR2 U20275 ( .A(n4264), .B(n3901), .Z(n3903) );
  MUX21L U20276 ( .A(n1518), .B(n3900), .S(n4291), .Z(n3902) );
  NR2 U20277 ( .A(n4341), .B(n4292), .Z(n3901) );
  ND2 U20278 ( .A(n2980), .B(n4392), .Z(n1517) );
  ND2 U20279 ( .A(n5233), .B(n4946), .Z(n2980) );
  EO U20280 ( .A(n5227), .B(n4577), .Z(n790) );
  MUX21L U20281 ( .A(n4176), .B(n4175), .S(n4261), .Z(n4184) );
  NR2 U20282 ( .A(n4334), .B(n4186), .Z(n4175) );
  NR3 U20283 ( .A(n4334), .B(n393), .C(n4295), .Z(n4176) );
  AN3 U20284 ( .A(n4375), .B(n4251), .C(n4288), .Z(n3924) );
  MUX21L U20285 ( .A(n4179), .B(n4180), .S(n4334), .Z(n4182) );
  ND2 U20286 ( .A(n3278), .B(n3277), .Z(n1505) );
  ND2 U20287 ( .A(n4295), .B(n4259), .Z(n4181) );
  MUX21L U20288 ( .A(n3935), .B(n3934), .S(n4292), .Z(n3940) );
  NR3 U20289 ( .A(n4337), .B(n396), .C(n4263), .Z(n3934) );
  NR2 U20290 ( .A(n4337), .B(n765), .Z(n3935) );
  MUX21L U20291 ( .A(n3936), .B(n3937), .S(n4263), .Z(n3938) );
  NR2 U20292 ( .A(n4338), .B(n4292), .Z(n3937) );
  AN3 U20293 ( .A(n4288), .B(n1502), .C(n4332), .Z(n3936) );
  NR2 U20294 ( .A(n4935), .B(n4606), .Z(n1502) );
  MUX21L U20295 ( .A(n3943), .B(n3944), .S(n4292), .Z(n3945) );
  NR2 U20296 ( .A(n4262), .B(n398), .Z(n3944) );
  NR3 U20297 ( .A(n4263), .B(n4338), .C(n399), .Z(n3943) );
  MUX21L U20298 ( .A(n3950), .B(n3949), .S(n4292), .Z(n3951) );
  ND2 U20299 ( .A(n3947), .B(n1497), .Z(n3949) );
  ND2 U20300 ( .A(n3948), .B(n1499), .Z(n3950) );
  NR2 U20301 ( .A(n4338), .B(n4262), .Z(n3947) );
  NR2 U20302 ( .A(n4338), .B(n4262), .Z(n3948) );
  NR2 U20303 ( .A(n4222), .B(n413), .Z(n4064) );
  ND3 U20304 ( .A(n4340), .B(n842), .C(n4293), .Z(n4007) );
  MUX41 U20305 ( .D0(n1087), .D1(n1070), .D2(n1078), .D3(n1062), .A(n4210), 
        .B(n4219), .Z(N229) );
  MUX21L U20306 ( .A(n3790), .B(n3791), .S(n4295), .Z(n3799) );
  NR2 U20307 ( .A(n4353), .B(n760), .Z(n3791) );
  NR3 U20308 ( .A(n4353), .B(n780), .C(n4266), .Z(n3790) );
  ND2 U20309 ( .A(n4066), .B(n4065), .Z(N220) );
  AO2 U20310 ( .A(n4222), .B(n841), .C(n4222), .D(n4208), .Z(n4066) );
  MUX21L U20311 ( .A(n4064), .B(n839), .S(n4208), .Z(n4065) );
  ND3 U20312 ( .A(n3880), .B(n3879), .C(n3878), .Z(n841) );
  NR3 U20313 ( .A(n418), .B(n4347), .C(n4291), .Z(n3822) );
  ND2 U20314 ( .A(n4759), .B(n5199), .Z(n2497) );
  NR3 U20315 ( .A(n2661), .B(n4296), .C(n4267), .Z(n3710) );
  NR2 U20316 ( .A(n4340), .B(n4197), .Z(n4021) );
  IVP U20317 ( .A(n831), .Z(n4197) );
  AO4 U20318 ( .A(n4926), .B(n4576), .C(n5249), .D(n4576), .Z(n831) );
  NR2 U20319 ( .A(n4294), .B(n419), .Z(n4132) );
  ND2 U20320 ( .A(n5292), .B(n4970), .Z(n2660) );
  NR2 U20321 ( .A(n3761), .B(n3760), .Z(n3763) );
  NR2 U20322 ( .A(n4352), .B(n4296), .Z(n3761) );
  NR2 U20323 ( .A(n4296), .B(n780), .Z(n3760) );
  ND2 U20324 ( .A(n2955), .B(n2954), .Z(n984) );
  EO U20325 ( .A(n5221), .B(n4563), .Z(n982) );
  AO7 U20326 ( .A(n5277), .B(n4964), .C(n4472), .Z(n937) );
  ND2 U20327 ( .A(n2066), .B(n2065), .Z(n933) );
  ND3 U20328 ( .A(n2346), .B(n2345), .C(n2344), .Z(n939) );
  AN3 U20329 ( .A(n4290), .B(n1006), .C(n4333), .Z(n3821) );
  ND3 U20330 ( .A(n2575), .B(n2574), .C(n2573), .Z(n1006) );
  ND2 U20331 ( .A(n4974), .B(n4523), .Z(n2573) );
  ND2 U20332 ( .A(n4974), .B(n5289), .Z(n2575) );
  AN3 U20333 ( .A(n4288), .B(n767), .C(n4331), .Z(n3894) );
  MUX41 U20334 ( .D0(n1057), .D1(n1039), .D2(n1048), .D3(n1034), .A(n4210), 
        .B(n4219), .Z(N228) );
  ND4 U20335 ( .A(n4059), .B(n4058), .C(n4057), .D(n4056), .Z(n1034) );
  MUX41 U20336 ( .D0(n1027), .D1(n1009), .D2(n1018), .D3(n1003), .A(n4210), 
        .B(n4218), .Z(N227) );
  MUX41 U20337 ( .D0(n996), .D1(n980), .D2(n987), .D3(n972), .A(n4210), .B(
        n4218), .Z(N226) );
  MUX41 U20338 ( .D0(n964), .D1(n949), .D2(n957), .D3(n940), .A(n4210), .B(
        n4218), .Z(N225) );
  MUX41 U20339 ( .D0(n932), .D1(n915), .D2(n924), .D3(n906), .A(n4210), .B(
        n4218), .Z(N224) );
  MUX41 U20340 ( .D0(n876), .D1(n861), .D2(n867), .D3(n859), .A(n4210), .B(
        n4218), .Z(N222) );
  ND2 U20341 ( .A(n3763), .B(n3762), .Z(n861) );
  ND2 U20342 ( .A(n3729), .B(n3728), .Z(n859) );
  MUX21L U20343 ( .A(n4015), .B(n835), .S(n4261), .Z(n4020) );
  NR3 U20344 ( .A(n4584), .B(n5234), .C(n4957), .Z(n835) );
  MUX21L U20345 ( .A(n4134), .B(n4133), .S(n4258), .Z(n4135) );
  AN3 U20346 ( .A(n4290), .B(n1038), .C(n4334), .Z(n4134) );
  AN3 U20347 ( .A(n4333), .B(n4289), .C(n1035), .Z(n4133) );
  ND2 U20348 ( .A(n2553), .B(n2552), .Z(n1038) );
  MUX21L U20349 ( .A(n4048), .B(n4049), .S(n4341), .Z(n4059) );
  NR3 U20350 ( .A(n420), .B(n4294), .C(n4261), .Z(n4048) );
  ND2 U20351 ( .A(n4023), .B(n4022), .Z(n832) );
  AO6 U20352 ( .A(n4340), .B(n4293), .C(n4261), .Z(n4023) );
  MUX21L U20353 ( .A(n4021), .B(n830), .S(n4293), .Z(n4022) );
  ND2 U20354 ( .A(n3476), .B(n3475), .Z(n830) );
  AN3 U20355 ( .A(n882), .B(n4290), .C(n4331), .Z(n3794) );
  ND2 U20356 ( .A(n2586), .B(n4521), .Z(n882) );
  ND2 U20357 ( .A(n5290), .B(n4973), .Z(n2586) );
  AO4 U20358 ( .A(n4978), .B(n4635), .C(n5263), .D(n4635), .Z(n880) );
  NR3 U20359 ( .A(n5133), .B(n4296), .C(n4267), .Z(n3700) );
  NR2 U20360 ( .A(n4336), .B(n4294), .Z(n4127) );
  NR2 U20361 ( .A(n4336), .B(n4294), .Z(n4128) );
  NR2 U20362 ( .A(n4336), .B(n4978), .Z(n4130) );
  AN3 U20363 ( .A(n902), .B(n4252), .C(n4289), .Z(n3711) );
  ND3 U20364 ( .A(n4854), .B(n5170), .C(n4454), .Z(n902) );
  ND2 U20365 ( .A(n4291), .B(n833), .Z(n3816) );
  ND2 U20366 ( .A(n2590), .B(n4520), .Z(n833) );
  ND2 U20367 ( .A(n5290), .B(n4973), .Z(n2590) );
  ND2 U20368 ( .A(n4291), .B(n846), .Z(n3814) );
  ND2 U20369 ( .A(n2588), .B(n4521), .Z(n846) );
  ND2 U20370 ( .A(n5290), .B(n4973), .Z(n2588) );
  NR2 U20371 ( .A(n4336), .B(n4291), .Z(n3895) );
  AN3 U20372 ( .A(n1058), .B(n4252), .C(n4288), .Z(n3701) );
  ND2 U20373 ( .A(n4453), .B(n4855), .Z(n1058) );
  AN3 U20374 ( .A(n862), .B(n4251), .C(n4331), .Z(n3893) );
  ND3 U20375 ( .A(n4748), .B(n5197), .C(n4498), .Z(n862) );
  AN3 U20376 ( .A(n851), .B(n4332), .C(n4251), .Z(n3996) );
  ND3 U20377 ( .A(n4832), .B(n5089), .C(n4437), .Z(n851) );
  AN3 U20378 ( .A(n1980), .B(n4276), .C(n4333), .Z(n4156) );
  MUX21L U20379 ( .A(n3035), .B(n3034), .S(n5240), .Z(n1980) );
  ND2 U20380 ( .A(n4386), .B(n4815), .Z(n3035) );
  ND2 U20381 ( .A(n4943), .B(n4385), .Z(n3034) );
  AN3 U20382 ( .A(n1978), .B(n4276), .C(n4333), .Z(n4155) );
  NR2 U20383 ( .A(n4562), .B(n5193), .Z(n1978) );
  MUX21L U20384 ( .A(n4094), .B(n4093), .S(n4261), .Z(n4102) );
  NR2 U20385 ( .A(n4339), .B(n365), .Z(n4093) );
  AN3 U20386 ( .A(n1465), .B(n4309), .C(n4289), .Z(n4094) );
  AN3 U20387 ( .A(n1466), .B(n4277), .C(n4333), .Z(n4096) );
  MUX21L U20388 ( .A(n2671), .B(n5207), .S(n4970), .Z(n1466) );
  ND2 U20389 ( .A(n4625), .B(n5207), .Z(n2671) );
  IVP U20390 ( .A(n350), .Z(n4290) );
  IVP U20391 ( .A(n350), .Z(n4295) );
  IVP U20392 ( .A(n4276), .Z(n4306) );
  AN3 U20393 ( .A(n1409), .B(n4230), .C(n4331), .Z(n3881) );
  ND2 U20394 ( .A(n5235), .B(n3075), .Z(n1409) );
  ND2 U20395 ( .A(n4941), .B(n4579), .Z(n3075) );
  IVP U20396 ( .A(n4276), .Z(n4301) );
  IVP U20397 ( .A(n4280), .Z(n4292) );
  IVP U20398 ( .A(n4281), .Z(n4294) );
  IVP U20399 ( .A(n350), .Z(n4289) );
  IVP U20400 ( .A(n4276), .Z(n4302) );
  IVP U20401 ( .A(n4229), .Z(n4258) );
  IVP U20402 ( .A(n4224), .Z(n4253) );
  IVP U20403 ( .A(n4224), .Z(n4256) );
  IVP U20404 ( .A(n4310), .Z(n4335) );
  IVP U20405 ( .A(n4230), .Z(n4260) );
  IVP U20406 ( .A(n4312), .Z(n4334) );
  IVP U20407 ( .A(n4311), .Z(n4333) );
  IVP U20408 ( .A(n4223), .Z(n4257) );
  IVP U20409 ( .A(n4311), .Z(n4339) );
  IVP U20410 ( .A(n4312), .Z(n4350) );
  NR2 U20411 ( .A(n4335), .B(n4229), .Z(n4151) );
  IVP U20412 ( .A(n4286), .Z(n4291) );
  IVP U20413 ( .A(n4312), .Z(n4345) );
  IVP U20414 ( .A(n4312), .Z(n4346) );
  IVP U20415 ( .A(n4225), .Z(n4261) );
  IVP U20416 ( .A(n4312), .Z(n4349) );
  ND4 U20417 ( .A(n3992), .B(n3991), .C(n3990), .D(n3989), .Z(n1388) );
  ND4 U20418 ( .A(n1386), .B(n4293), .C(n4229), .D(n4316), .Z(n3989) );
  MUX21L U20419 ( .A(n3988), .B(n3987), .S(n4293), .Z(n3990) );
  MUX21L U20420 ( .A(n3985), .B(n3986), .S(n4293), .Z(n3991) );
  AN3 U20421 ( .A(n1387), .B(n4228), .C(n4332), .Z(n3985) );
  ND2 U20422 ( .A(n3507), .B(n3506), .Z(n1387) );
  ND3 U20423 ( .A(n4921), .B(n4423), .C(n5245), .Z(n3506) );
  MUX21L U20424 ( .A(n3504), .B(n3505), .S(n4921), .Z(n3507) );
  MUX21L U20425 ( .A(n3983), .B(n3984), .S(n4339), .Z(n3992) );
  AN3 U20426 ( .A(n1384), .B(n4281), .C(n4250), .Z(n3983) );
  AN3 U20427 ( .A(n1383), .B(n4281), .C(n4251), .Z(n3984) );
  ND2 U20428 ( .A(n4608), .B(n5072), .Z(n1384) );
  IVP U20429 ( .A(n4309), .Z(n4331) );
  IVP U20430 ( .A(n4225), .Z(n4264) );
  IVP U20431 ( .A(n4310), .Z(n4336) );
  IVP U20432 ( .A(n353), .Z(n4208) );
  AN3 U20433 ( .A(n1867), .B(n4316), .C(n4252), .Z(n4108) );
  MUX21L U20434 ( .A(n2393), .B(n5264), .S(n4636), .Z(n1867) );
  ND2 U20435 ( .A(n5264), .B(n4977), .Z(n2393) );
  AN3 U20436 ( .A(n1385), .B(n4226), .C(n4332), .Z(n3987) );
  MUX21L U20437 ( .A(n4543), .B(n4789), .S(n5259), .Z(n1385) );
  IVP U20438 ( .A(n4276), .Z(n4305) );
  IVP U20439 ( .A(n4282), .Z(n4293) );
  IVP U20440 ( .A(n4204), .Z(n4209) );
  IVP U20441 ( .A(n351), .Z(n4221) );
  IVP U20442 ( .A(n4223), .Z(n4251) );
  ND4 U20443 ( .A(n3673), .B(n3672), .C(n3671), .D(n3670), .Z(n1329) );
  ND4 U20444 ( .A(n1327), .B(n4297), .C(n4249), .D(n4329), .Z(n3670) );
  MUX21L U20445 ( .A(n3664), .B(n3665), .S(n4351), .Z(n3673) );
  MUX21L U20446 ( .A(n3666), .B(n3667), .S(n4351), .Z(n3672) );
  MUX21L U20447 ( .A(n3669), .B(n3668), .S(n4268), .Z(n3671) );
  NR3 U20448 ( .A(n369), .B(n4351), .C(n4297), .Z(n3669) );
  AN3 U20449 ( .A(n1325), .B(n4279), .C(n4332), .Z(n3668) );
  IVP U20450 ( .A(n4216), .Z(n4220) );
  IVP U20451 ( .A(n4225), .Z(n4262) );
  IVP U20452 ( .A(n4316), .Z(n4332) );
  AN3 U20453 ( .A(n1326), .B(n4224), .C(n4288), .Z(n3667) );
  MUX21L U20454 ( .A(n5162), .B(n2174), .S(n4967), .Z(n1326) );
  ND2 U20455 ( .A(n4463), .B(n5162), .Z(n2174) );
  IVP U20456 ( .A(n4224), .Z(n4254) );
  ND4 U20457 ( .A(n3776), .B(n3775), .C(n3774), .D(n3773), .Z(n1308) );
  ND4 U20458 ( .A(n1305), .B(n4296), .C(n4244), .D(n4325), .Z(n3773) );
  MUX21L U20459 ( .A(n3769), .B(n3770), .S(n4296), .Z(n3775) );
  MUX21L U20460 ( .A(n3767), .B(n3768), .S(n4352), .Z(n3776) );
  AN3 U20461 ( .A(n1870), .B(n4317), .C(n4289), .Z(n4105) );
  ND2 U20462 ( .A(n4894), .B(n5208), .Z(n1870) );
  AN3 U20463 ( .A(n1303), .B(n4282), .C(n4252), .Z(n3767) );
  ND2 U20464 ( .A(n2490), .B(n2489), .Z(n1303) );
  ND2 U20465 ( .A(n5287), .B(n4760), .Z(n2489) );
  MUX21L U20466 ( .A(n2488), .B(n4475), .S(n5286), .Z(n2490) );
  MUX21L U20467 ( .A(n3772), .B(n3771), .S(n4296), .Z(n3774) );
  NR3 U20468 ( .A(n4266), .B(n4353), .C(n4191), .Z(n3772) );
  AN3 U20469 ( .A(n1304), .B(n4226), .C(n4331), .Z(n3771) );
  IVP U20470 ( .A(n1307), .Z(n4191) );
  MUX21L U20471 ( .A(n4040), .B(n4041), .S(n4341), .Z(n4045) );
  AN3 U20472 ( .A(n4721), .B(n4285), .C(n4251), .Z(n4040) );
  ND2 U20473 ( .A(n2178), .B(n2177), .Z(n1297) );
  IVP U20474 ( .A(n4284), .Z(n4297) );
  IVP U20475 ( .A(n4310), .Z(n4337) );
  IVP U20476 ( .A(n4310), .Z(n4338) );
  IVP U20477 ( .A(n4223), .Z(n4252) );
  AN3 U20478 ( .A(n5070), .B(n4286), .C(n4253), .Z(n3664) );
  AN3 U20479 ( .A(n1302), .B(n4278), .C(n4252), .Z(n3768) );
  AO7 U20480 ( .A(n5267), .B(n4527), .C(n4915), .Z(n1302) );
  AN3 U20481 ( .A(n1306), .B(n4226), .C(n4331), .Z(n3769) );
  MUX21L U20482 ( .A(n5205), .B(n4757), .S(n4626), .Z(n1306) );
  AN3 U20483 ( .A(n1298), .B(n4314), .C(n4289), .Z(n4038) );
  ND2 U20484 ( .A(n2245), .B(n2244), .Z(n1298) );
  ND2 U20485 ( .A(n5276), .B(n4866), .Z(n2244) );
  MUX21L U20486 ( .A(n2243), .B(n4471), .S(n5276), .Z(n2245) );
  AN3 U20487 ( .A(n1299), .B(n4285), .C(n4332), .Z(n4042) );
  EN U20488 ( .A(n5222), .B(n4630), .Z(n1299) );
  IVP U20489 ( .A(n4226), .Z(n4268) );
  IVP U20490 ( .A(n4313), .Z(n4351) );
  IVP U20491 ( .A(n4311), .Z(n4344) );
  IVP U20492 ( .A(n4283), .Z(n4296) );
  IVP U20493 ( .A(n4312), .Z(n4348) );
  IVP U20494 ( .A(n4311), .Z(n4341) );
  IVP U20495 ( .A(n4217), .Z(n4219) );
  IVP U20496 ( .A(n4280), .Z(n4288) );
  AN3 U20497 ( .A(n1276), .B(n4277), .C(n4333), .Z(n4084) );
  ND2 U20498 ( .A(n2652), .B(n2651), .Z(n1276) );
  ND2 U20499 ( .A(n4971), .B(n5208), .Z(n2651) );
  MUX21L U20500 ( .A(n2650), .B(n4514), .S(n4971), .Z(n2652) );
  IVP U20501 ( .A(n4247), .Z(n4259) );
  IVP U20502 ( .A(n4226), .Z(n4266) );
  IVP U20503 ( .A(n4313), .Z(n4352) );
  IVP U20504 ( .A(n4313), .Z(n4353) );
  MUX21L U20505 ( .A(n4029), .B(n4028), .S(n4260), .Z(n4033) );
  AN3 U20506 ( .A(n1761), .B(n4314), .C(n4289), .Z(n4029) );
  EN U20507 ( .A(n5221), .B(n4964), .Z(n1761) );
  IVP U20508 ( .A(n4276), .Z(n4304) );
  IVP U20509 ( .A(n4311), .Z(n4340) );
  NR2 U20510 ( .A(n4341), .B(n4230), .Z(n4079) );
  ND4 U20511 ( .A(n4126), .B(n4125), .C(n4124), .D(n4123), .Z(n1250) );
  MUX21L U20512 ( .A(n4118), .B(n4117), .S(n4260), .Z(n4126) );
  MUX21L U20513 ( .A(n4120), .B(n4119), .S(n4258), .Z(n4125) );
  AO2 U20514 ( .A(n4116), .B(n4229), .C(n4115), .D(n1248), .Z(n4124) );
  AN3 U20515 ( .A(n4547), .B(n4277), .C(n4333), .Z(n4083) );
  MUX21L U20516 ( .A(n4143), .B(n4144), .S(n4336), .Z(n4148) );
  AN3 U20517 ( .A(n1253), .B(n4277), .C(n4253), .Z(n4143) );
  AN3 U20518 ( .A(n4899), .B(n4545), .C(n5227), .Z(n1254) );
  IVP U20519 ( .A(n4276), .Z(n4300) );
  IVP U20520 ( .A(n4224), .Z(n4255) );
  ND4 U20521 ( .A(n3739), .B(n3738), .C(n3737), .D(n3736), .Z(n1732) );
  ND4 U20522 ( .A(n1731), .B(n4296), .C(n4245), .D(n4326), .Z(n3736) );
  MUX21L U20523 ( .A(n3732), .B(n3733), .S(n4352), .Z(n3738) );
  MUX21L U20524 ( .A(n3735), .B(n3734), .S(n4296), .Z(n3737) );
  AN3 U20525 ( .A(n1256), .B(n4277), .C(n4334), .Z(n4145) );
  MUX21L U20526 ( .A(n4554), .B(n5234), .S(n4942), .Z(n1256) );
  AN3 U20527 ( .A(n1255), .B(n4313), .C(n4290), .Z(n4141) );
  MUX21L U20528 ( .A(n5235), .B(n4945), .S(n4551), .Z(n1255) );
  AN3 U20529 ( .A(n1247), .B(n4277), .C(n4333), .Z(n4119) );
  EO U20530 ( .A(n5224), .B(n4617), .Z(n1247) );
  MUX21L U20531 ( .A(n3730), .B(n3731), .S(n4352), .Z(n3739) );
  AN3 U20532 ( .A(n1729), .B(n4283), .C(n4252), .Z(n3730) );
  AN3 U20533 ( .A(n1728), .B(n4279), .C(n4252), .Z(n3731) );
  MUX21L U20534 ( .A(n4767), .B(n2136), .S(n5273), .Z(n1729) );
  AN3 U20535 ( .A(n1730), .B(n4225), .C(n4331), .Z(n3734) );
  ND2 U20536 ( .A(n2222), .B(n2221), .Z(n1730) );
  ND2 U20537 ( .A(n4595), .B(n4965), .Z(n2221) );
  MUX21L U20538 ( .A(n2220), .B(n5160), .S(n4966), .Z(n2222) );
  MUX21L U20539 ( .A(n4167), .B(n4168), .S(n4259), .Z(n4172) );
  AN3 U20540 ( .A(n1224), .B(n4313), .C(n4290), .Z(n4168) );
  ND2 U20541 ( .A(n3047), .B(n3046), .Z(n1227) );
  NR2 U20542 ( .A(n4260), .B(n4314), .Z(n4024) );
  AN3 U20543 ( .A(n5071), .B(n4315), .C(n4290), .Z(n4117) );
  IVP U20544 ( .A(n4312), .Z(n4347) );
  IVP U20545 ( .A(n4226), .Z(n4267) );
  NR2 U20546 ( .A(n4262), .B(n4284), .Z(n4164) );
  ND4 U20547 ( .A(n3921), .B(n3920), .C(n3919), .D(n3918), .Z(n1695) );
  ND4 U20548 ( .A(n1694), .B(n4292), .C(n4238), .D(n4320), .Z(n3918) );
  MUX21L U20549 ( .A(n3914), .B(n3915), .S(n4337), .Z(n3920) );
  MUX21L U20550 ( .A(n3912), .B(n3913), .S(n4337), .Z(n3921) );
  ND4 U20551 ( .A(n3683), .B(n3682), .C(n3681), .D(n3680), .Z(n1186) );
  ND4 U20552 ( .A(n1185), .B(n4297), .C(n4248), .D(n4328), .Z(n3680) );
  MUX21L U20553 ( .A(n3676), .B(n3677), .S(n4351), .Z(n3682) );
  MUX21L U20554 ( .A(n3674), .B(n3675), .S(n4351), .Z(n3683) );
  AN3 U20555 ( .A(n1692), .B(n4278), .C(n4251), .Z(n3912) );
  MUX21L U20556 ( .A(n3289), .B(n3288), .S(n5254), .Z(n1692) );
  ND2 U20557 ( .A(n4486), .B(n4844), .Z(n3289) );
  ND2 U20558 ( .A(n4610), .B(n4844), .Z(n3288) );
  AN3 U20559 ( .A(n1184), .B(n4224), .C(n4288), .Z(n3677) );
  AO7 U20560 ( .A(n5274), .B(n4967), .C(n4597), .Z(n1184) );
  MUX21L U20561 ( .A(n3917), .B(n3916), .S(n4263), .Z(n3919) );
  NR3 U20562 ( .A(n377), .B(n4337), .C(n4292), .Z(n3917) );
  AN3 U20563 ( .A(n1691), .B(n4278), .C(n4332), .Z(n3916) );
  MUX21L U20564 ( .A(n3679), .B(n3678), .S(n4268), .Z(n3681) );
  AN3 U20565 ( .A(n1183), .B(n4278), .C(n4331), .Z(n3678) );
  NR3 U20566 ( .A(n379), .B(n4351), .C(n4297), .Z(n3679) );
  NR2 U20567 ( .A(n4911), .B(n4602), .Z(n1183) );
  IVP U20568 ( .A(n4276), .Z(n4303) );
  AN3 U20569 ( .A(n1693), .B(n4248), .C(n4288), .Z(n3915) );
  AO7 U20570 ( .A(n4604), .B(n5107), .C(n3382), .Z(n1693) );
  ND2 U20571 ( .A(n5258), .B(n4936), .Z(n3382) );
  AN3 U20572 ( .A(n4547), .B(n4285), .C(n4253), .Z(n3674) );
  ND4 U20573 ( .A(n3645), .B(n3644), .C(n3643), .D(n3642), .Z(n1640) );
  MUX21L U20574 ( .A(n3641), .B(n3640), .S(n4268), .Z(n3643) );
  ND4 U20575 ( .A(n1639), .B(n4297), .C(n4241), .D(n4317), .Z(n3642) );
  MUX21L U20576 ( .A(n3636), .B(n3637), .S(n4350), .Z(n3645) );
  MUX21L U20577 ( .A(n3638), .B(n3639), .S(n4350), .Z(n3644) );
  AN3 U20578 ( .A(n1635), .B(n4253), .C(n4288), .Z(n3638) );
  AN3 U20579 ( .A(n1638), .B(n4223), .C(n4288), .Z(n3639) );
  ND3 U20580 ( .A(n4855), .B(n5170), .C(n4453), .Z(n1635) );
  IVP U20581 ( .A(n4311), .Z(n4343) );
  AN3 U20582 ( .A(n1637), .B(n4278), .C(n4253), .Z(n3636) );
  ND2 U20583 ( .A(n2166), .B(n2165), .Z(n1637) );
  ND2 U20584 ( .A(n5274), .B(n4598), .Z(n2166) );
  ND2 U20585 ( .A(n4968), .B(n4598), .Z(n2165) );
  AN3 U20586 ( .A(n1636), .B(n4287), .C(n4332), .Z(n3640) );
  AO4 U20587 ( .A(n4911), .B(n4602), .C(n5272), .D(n4602), .Z(n1636) );
  IVP U20588 ( .A(n4276), .Z(n4299) );
  IVP U20589 ( .A(n4207), .Z(n4210) );
  IVP U20590 ( .A(n4225), .Z(n4263) );
  NR2 U20591 ( .A(n4297), .B(n4248), .Z(n3689) );
  ND4 U20592 ( .A(n3858), .B(n3857), .C(n3856), .D(n3855), .Z(n1149) );
  MUX21L U20593 ( .A(n3854), .B(n3853), .S(n4265), .Z(n3856) );
  ND4 U20594 ( .A(n1147), .B(n4291), .C(n4240), .D(n4322), .Z(n3855) );
  MUX21L U20595 ( .A(n3851), .B(n3852), .S(n4335), .Z(n3857) );
  ND4 U20596 ( .A(n3809), .B(n3808), .C(n3807), .D(n3806), .Z(n1143) );
  ND3 U20597 ( .A(n1142), .B(n4325), .C(n4243), .Z(n3806) );
  MUX21L U20598 ( .A(n3804), .B(n3805), .S(n4266), .Z(n3807) );
  MUX21L U20599 ( .A(n3802), .B(n3803), .S(n4295), .Z(n3808) );
  AN3 U20600 ( .A(n1146), .B(n4228), .C(n4288), .Z(n3852) );
  ND2 U20601 ( .A(n2977), .B(n2976), .Z(n1146) );
  ND2 U20602 ( .A(n4946), .B(n4551), .Z(n2976) );
  MUX21L U20603 ( .A(n2975), .B(n4551), .S(n5231), .Z(n2977) );
  AN3 U20604 ( .A(n1141), .B(n4330), .C(n4289), .Z(n3804) );
  ND2 U20605 ( .A(n4975), .B(n4619), .Z(n1141) );
  MUX21L U20606 ( .A(n3849), .B(n3850), .S(n4334), .Z(n3858) );
  NR3 U20607 ( .A(n382), .B(n4290), .C(n4265), .Z(n3850) );
  AN3 U20608 ( .A(n1145), .B(n4280), .C(n4251), .Z(n3849) );
  MUX21L U20609 ( .A(n3800), .B(n3801), .S(n4353), .Z(n3809) );
  NR2 U20610 ( .A(n4295), .B(n4266), .Z(n3800) );
  AN3 U20611 ( .A(n1140), .B(n4279), .C(n4252), .Z(n3801) );
  ND2 U20612 ( .A(n2480), .B(n4473), .Z(n1140) );
  MUX21L U20613 ( .A(n3693), .B(n3694), .S(n4267), .Z(n3696) );
  AN3 U20614 ( .A(n4279), .B(n4318), .C(n4359), .Z(n3694) );
  ND2 U20615 ( .A(n2306), .B(n2305), .Z(n1137) );
  NR2 U20616 ( .A(n4267), .B(n4286), .Z(n3688) );
  ND4 U20617 ( .A(n3868), .B(n3867), .C(n3866), .D(n3865), .Z(n1127) );
  ND3 U20618 ( .A(n759), .B(n4285), .C(n4264), .Z(n3865) );
  MUX21L U20619 ( .A(n3859), .B(n3860), .S(n4290), .Z(n3868) );
  MUX21L U20620 ( .A(n3863), .B(n3864), .S(n4264), .Z(n3866) );
  ND3 U20621 ( .A(n1605), .B(n4287), .C(n4268), .Z(n3652) );
  ND2 U20622 ( .A(n2168), .B(n2167), .Z(n1605) );
  ND2 U20623 ( .A(n5274), .B(n4598), .Z(n2168) );
  ND2 U20624 ( .A(n4968), .B(n4598), .Z(n2167) );
  MUX21L U20625 ( .A(n3646), .B(n3647), .S(n4297), .Z(n3655) );
  NR3 U20626 ( .A(n383), .B(n4350), .C(n4268), .Z(n3646) );
  AN3 U20627 ( .A(n1604), .B(n4327), .C(n4253), .Z(n3647) );
  MUX21L U20628 ( .A(n3650), .B(n3651), .S(n4268), .Z(n3653) );
  NR2 U20629 ( .A(n4297), .B(n4329), .Z(n3651) );
  AN3 U20630 ( .A(n1606), .B(n4332), .C(n4288), .Z(n3650) );
  NR2 U20631 ( .A(n4968), .B(n4597), .Z(n1606) );
  MUX21L U20632 ( .A(n3648), .B(n3649), .S(n4350), .Z(n3654) );
  AN3 U20633 ( .A(n1607), .B(n4223), .C(n4288), .Z(n3648) );
  NR2 U20634 ( .A(n4297), .B(n755), .Z(n3649) );
  ND3 U20635 ( .A(n4869), .B(n5154), .C(n4543), .Z(n1607) );
  MUX21L U20636 ( .A(n3861), .B(n3862), .S(n4335), .Z(n3867) );
  AN3 U20637 ( .A(n1126), .B(n4228), .C(n4288), .Z(n3861) );
  NR2 U20638 ( .A(n4290), .B(n756), .Z(n3862) );
  ND2 U20639 ( .A(n3027), .B(n3026), .Z(n1126) );
  IVP U20640 ( .A(n4226), .Z(n4265) );
  AN3 U20641 ( .A(n4359), .B(n4279), .C(n4331), .Z(n3853) );
  AN3 U20642 ( .A(n1124), .B(n4313), .C(n4251), .Z(n3860) );
  NR2 U20643 ( .A(n4928), .B(n4560), .Z(n1124) );
  MUX21L U20644 ( .A(n4073), .B(n4074), .S(n4259), .Z(n4075) );
  AN3 U20645 ( .A(n1585), .B(n4277), .C(n4333), .Z(n4073) );
  AO4 U20646 ( .A(n4915), .B(n4616), .C(n5267), .D(n4616), .Z(n1582) );
  ND2 U20647 ( .A(n2481), .B(n4474), .Z(n1122) );
  ND2 U20648 ( .A(n5268), .B(n4917), .Z(n2481) );
  ND2 U20649 ( .A(n3751), .B(n3750), .Z(N173) );
  ND3 U20650 ( .A(n1110), .B(n4204), .C(n4221), .Z(n3750) );
  NR2 U20651 ( .A(n4353), .B(n4282), .Z(n3805) );
  ND3 U20652 ( .A(n4247), .B(n4286), .C(n1120), .Z(n3698) );
  AO7 U20653 ( .A(n5260), .B(n4963), .C(n4629), .Z(n1120) );
  ND2 U20654 ( .A(n4296), .B(n4248), .Z(n3695) );
  AO3 U20655 ( .A(n764), .B(n3875), .C(n3874), .D(n3873), .Z(n1110) );
  ND2 U20656 ( .A(n4240), .B(n4282), .Z(n3875) );
  MUX21L U20657 ( .A(n3871), .B(n3872), .S(n4336), .Z(n3873) );
  NR2 U20658 ( .A(n4290), .B(n4322), .Z(n3864) );
  ND2 U20659 ( .A(n4285), .B(n4326), .Z(n3758) );
  ND2 U20660 ( .A(n1109), .B(n4286), .Z(n3757) );
  AO4 U20661 ( .A(n4915), .B(n4617), .C(n5267), .D(n4617), .Z(n1109) );
  AN3 U20662 ( .A(n4547), .B(n4314), .C(n4289), .Z(n4069) );
  MUX21L U20663 ( .A(n3656), .B(n3657), .S(n4351), .Z(n3661) );
  NR2 U20664 ( .A(n4268), .B(n4287), .Z(n3657) );
  NR3 U20665 ( .A(n760), .B(n4297), .C(n4268), .Z(n3656) );
  ND2 U20666 ( .A(n4063), .B(n4203), .Z(N172) );
  MUX21L U20667 ( .A(n1108), .B(n1102), .S(n4222), .Z(n4063) );
  ND4 U20668 ( .A(n3965), .B(n3964), .C(n3963), .D(n3962), .Z(n1108) );
  ND4 U20669 ( .A(n1107), .B(n4292), .C(n4234), .D(n4318), .Z(n3962) );
  MUX21L U20670 ( .A(n3956), .B(n3957), .S(n4338), .Z(n3965) );
  MUX21L U20671 ( .A(n3958), .B(n3959), .S(n4338), .Z(n3964) );
  AN3 U20672 ( .A(n1583), .B(n4277), .C(n4252), .Z(n4071) );
  ND2 U20673 ( .A(n4525), .B(n4884), .Z(n1583) );
  MUX21L U20674 ( .A(n3961), .B(n3960), .S(n4262), .Z(n3963) );
  NR3 U20675 ( .A(n3523), .B(n4339), .C(n4292), .Z(n3961) );
  AN3 U20676 ( .A(n1104), .B(n4287), .C(n4332), .Z(n3960) );
  ND2 U20677 ( .A(n3753), .B(n3752), .Z(N171) );
  ND2 U20678 ( .A(n4222), .B(n4204), .Z(n3753) );
  NR2 U20679 ( .A(n4264), .B(n4287), .Z(n3872) );
  ND4 U20680 ( .A(n3836), .B(n3835), .C(n3834), .D(n3833), .Z(n1548) );
  MUX21L U20681 ( .A(n3832), .B(n3831), .S(n4265), .Z(n3834) );
  ND4 U20682 ( .A(n1547), .B(n4291), .C(n4242), .D(n4323), .Z(n3833) );
  MUX21L U20683 ( .A(n3827), .B(n3828), .S(n4334), .Z(n3836) );
  AN3 U20684 ( .A(n1106), .B(n4228), .C(n4288), .Z(n3959) );
  NR2 U20685 ( .A(n4605), .B(n4792), .Z(n1106) );
  AN3 U20686 ( .A(n1105), .B(n4287), .C(n4257), .Z(n3956) );
  AO7 U20687 ( .A(n5255), .B(n4949), .C(n4609), .Z(n1105) );
  ND3 U20688 ( .A(n4287), .B(n4328), .C(n4247), .Z(n3697) );
  ND2 U20689 ( .A(n1101), .B(n4204), .Z(n3752) );
  ND3 U20690 ( .A(n3974), .B(n3973), .C(n3972), .Z(n1101) );
  MUX21L U20691 ( .A(n3970), .B(n3971), .S(n4262), .Z(n3972) );
  MUX21L U20692 ( .A(n3966), .B(n3967), .S(n4262), .Z(n3973) );
  MUX21L U20693 ( .A(n3829), .B(n3830), .S(n4334), .Z(n3835) );
  AN3 U20694 ( .A(n1543), .B(n4251), .C(n4289), .Z(n3829) );
  AN3 U20695 ( .A(n1546), .B(n4227), .C(n4289), .Z(n3830) );
  NR2 U20696 ( .A(n4928), .B(n4560), .Z(n1543) );
  AO7 U20697 ( .A(n4186), .B(n3877), .C(n3876), .Z(n1102) );
  ND2 U20698 ( .A(n4239), .B(n4322), .Z(n3877) );
  ND2 U20699 ( .A(n4240), .B(n4282), .Z(n3876) );
  AN3 U20700 ( .A(n1545), .B(n4278), .C(n4251), .Z(n3827) );
  NR3 U20701 ( .A(n4565), .B(n5284), .C(n4933), .Z(n1545) );
  AN3 U20702 ( .A(n1100), .B(n4287), .C(n4332), .Z(n3966) );
  ND3 U20703 ( .A(n3517), .B(n3516), .C(n3515), .Z(n1100) );
  ND2 U20704 ( .A(n4420), .B(n4778), .Z(n3516) );
  ND2 U20705 ( .A(n5246), .B(n4778), .Z(n3517) );
  ND2 U20706 ( .A(n3789), .B(n3788), .Z(n1542) );
  MUX21L U20707 ( .A(n4243), .B(n3787), .S(n4295), .Z(n3788) );
  MUX21L U20708 ( .A(n3786), .B(n3785), .S(n4266), .Z(n3789) );
  ND2 U20709 ( .A(n3743), .B(n3742), .Z(N118) );
  ND3 U20710 ( .A(n1531), .B(n4207), .C(n4221), .Z(n3742) );
  MUX21L U20711 ( .A(n3741), .B(n3740), .S(n4208), .Z(n3743) );
  IVP U20712 ( .A(n4217), .Z(n4222) );
  AO3 U20713 ( .A(n4340), .B(n4014), .C(n4229), .D(n4013), .Z(n1097) );
  ND2 U20714 ( .A(n4281), .B(n1096), .Z(n4014) );
  MUX21L U20715 ( .A(n4011), .B(n4012), .S(n4293), .Z(n4013) );
  ND2 U20716 ( .A(n3578), .B(n3577), .Z(n1096) );
  AN3 U20717 ( .A(n1544), .B(n4278), .C(n4330), .Z(n3831) );
  ND3 U20718 ( .A(n4736), .B(n5190), .C(n4402), .Z(n1544) );
  ND2 U20719 ( .A(n4249), .B(n4287), .Z(n3662) );
  ND2 U20720 ( .A(n4249), .B(n4329), .Z(n3663) );
  MUX21L U20721 ( .A(n3745), .B(n3744), .S(n4221), .Z(N117) );
  ND2 U20722 ( .A(n1519), .B(n4207), .Z(n3744) );
  ND2 U20723 ( .A(n1527), .B(n4207), .Z(n3745) );
  ND2 U20724 ( .A(n3978), .B(n3977), .Z(n1094) );
  ND2 U20725 ( .A(n4293), .B(n4233), .Z(n3977) );
  MUX21L U20726 ( .A(n3976), .B(n3975), .S(n4339), .Z(n3978) );
  NR2 U20727 ( .A(n4262), .B(n4196), .Z(n3975) );
  AN3 U20728 ( .A(n1530), .B(n4281), .C(n4331), .Z(n3837) );
  ND2 U20729 ( .A(n4381), .B(n4822), .Z(n1530) );
  MUX21L U20730 ( .A(n3747), .B(n3746), .S(n4221), .Z(N116) );
  ND2 U20731 ( .A(n1511), .B(n4207), .Z(n3746) );
  ND2 U20732 ( .A(n1516), .B(n4206), .Z(n3747) );
  ND4 U20733 ( .A(n3931), .B(n3930), .C(n3929), .D(n3928), .Z(n1516) );
  ND4 U20734 ( .A(n1515), .B(n4292), .C(n4238), .D(n4320), .Z(n3928) );
  MUX21L U20735 ( .A(n3924), .B(n3925), .S(n4337), .Z(n3930) );
  MUX21L U20736 ( .A(n3927), .B(n3926), .S(n4263), .Z(n3929) );
  MUX21L U20737 ( .A(n3922), .B(n3923), .S(n4337), .Z(n3931) );
  NR3 U20738 ( .A(n391), .B(n4292), .C(n4263), .Z(n3923) );
  AN3 U20739 ( .A(n1513), .B(n4278), .C(n4251), .Z(n3922) );
  AN3 U20740 ( .A(n1512), .B(n4278), .C(n4332), .Z(n3926) );
  ND2 U20741 ( .A(n3276), .B(n3275), .Z(n1512) );
  ND2 U20742 ( .A(n5253), .B(n4611), .Z(n3276) );
  ND2 U20743 ( .A(n4950), .B(n4611), .Z(n3275) );
  AN3 U20744 ( .A(n1514), .B(n4233), .C(n4288), .Z(n3925) );
  MUX21L U20745 ( .A(n4606), .B(n3342), .S(n5257), .Z(n1514) );
  ND2 U20746 ( .A(n4606), .B(n4794), .Z(n3342) );
  ND4 U20747 ( .A(n4184), .B(n4183), .C(n4182), .D(n4181), .Z(n1509) );
  ND3 U20748 ( .A(n3848), .B(n3847), .C(n3846), .Z(n1511) );
  ND2 U20749 ( .A(n4241), .B(n4323), .Z(n3848) );
  ND2 U20750 ( .A(n4241), .B(n4284), .Z(n3846) );
  ND2 U20751 ( .A(n1510), .B(n4235), .Z(n3847) );
  ND2 U20752 ( .A(n3980), .B(n3979), .Z(n1092) );
  ND3 U20753 ( .A(n4232), .B(n4282), .C(n4339), .Z(n3979) );
  ND3 U20754 ( .A(n4233), .B(n4287), .C(n1091), .Z(n3980) );
  AO4 U20755 ( .A(n4925), .B(n4576), .C(n5249), .D(n4925), .Z(n1091) );
  MUX21L U20756 ( .A(n4177), .B(n4178), .S(n4295), .Z(n4183) );
  AN3 U20757 ( .A(n1508), .B(n4227), .C(n4333), .Z(n4177) );
  MUX21L U20758 ( .A(n4793), .B(n3343), .S(n4606), .Z(n1506) );
  ND3 U20759 ( .A(n3940), .B(n3939), .C(n3938), .Z(n1504) );
  ND3 U20760 ( .A(n4927), .B(n4410), .C(n5246), .Z(n1090) );
  MUX21L U20761 ( .A(n3932), .B(n3933), .S(n4263), .Z(n3939) );
  NR2 U20762 ( .A(n4292), .B(n4186), .Z(n3933) );
  AN3 U20763 ( .A(n1503), .B(n4287), .C(n4332), .Z(n3932) );
  ND2 U20764 ( .A(n3583), .B(n3582), .Z(n1089) );
  ND2 U20765 ( .A(n4413), .B(n5131), .Z(n3583) );
  AO2 U20766 ( .A(n3942), .B(n4338), .C(n3941), .D(n4338), .Z(n3946) );
  NR2 U20767 ( .A(n4263), .B(n4283), .Z(n3941) );
  NR2 U20768 ( .A(n4263), .B(n401), .Z(n3942) );
  ND2 U20769 ( .A(n3946), .B(n3945), .Z(n1501) );
  AN3 U20770 ( .A(n4202), .B(n4211), .C(n1500), .Z(n791) );
  NR2 U20771 ( .A(n4925), .B(n4576), .Z(n1088) );
  MUX21L U20772 ( .A(n4921), .B(n4571), .S(n5245), .Z(n1498) );
  MUX21L U20773 ( .A(n3953), .B(n3952), .S(n4338), .Z(n1496) );
  ND3 U20774 ( .A(n4237), .B(n4287), .C(n1495), .Z(n3952) );
  ND2 U20775 ( .A(n3548), .B(n4416), .Z(n1495) );
  EO U20776 ( .A(n5229), .B(n4924), .Z(n3548) );
  MUX21L U20777 ( .A(n3955), .B(n3954), .S(n4338), .Z(n1494) );
  ND3 U20778 ( .A(n4236), .B(n4280), .C(n1493), .Z(n3955) );
  MUX21L U20779 ( .A(n4575), .B(n3563), .S(n4924), .Z(n1493) );
  ND2 U20780 ( .A(n4574), .B(n5127), .Z(n3563) );
  ND3 U20781 ( .A(n4236), .B(n4287), .C(n1492), .Z(n3954) );
  AO4 U20782 ( .A(n4921), .B(n4571), .C(n5245), .D(n4571), .Z(n1492) );
  ND3 U20783 ( .A(n4237), .B(n4281), .C(n4415), .Z(n3953) );
  ND2 U20784 ( .A(n3622), .B(n3621), .Z(n1491) );
  EN U20785 ( .A(n5227), .B(n4578), .Z(n3622) );
  EO U20786 ( .A(n4901), .B(n4578), .Z(n3621) );
  MUX21L U20787 ( .A(n5248), .B(n4924), .S(n4575), .Z(n1490) );
  ND2 U20788 ( .A(n3565), .B(n3564), .Z(n1489) );
  ND2 U20789 ( .A(n4415), .B(n4773), .Z(n3565) );
  ND2 U20790 ( .A(n5248), .B(n4414), .Z(n3564) );
  AO4 U20791 ( .A(n4924), .B(n4575), .C(n5248), .D(n4575), .Z(n1488) );
  NR2 U20792 ( .A(n4925), .B(n4575), .Z(n1487) );
  NR2 U20793 ( .A(n4208), .B(n416), .Z(n3909) );
  ND2 U20794 ( .A(n4260), .B(n4284), .Z(n4018) );
  ND4 U20795 ( .A(n3708), .B(n3707), .C(n3706), .D(n3705), .Z(n1062) );
  MUX21L U20796 ( .A(n3699), .B(n3700), .S(n4351), .Z(n3708) );
  ND4 U20797 ( .A(n1061), .B(n4296), .C(n4247), .D(n4328), .Z(n3705) );
  MUX21L U20798 ( .A(n3701), .B(n3702), .S(n4352), .Z(n3707) );
  ND4 U20799 ( .A(n3799), .B(n3798), .C(n3797), .D(n3796), .Z(n884) );
  ND3 U20800 ( .A(n881), .B(n4325), .C(n4266), .Z(n3796) );
  MUX21L U20801 ( .A(n3792), .B(n3793), .S(n4295), .Z(n3798) );
  MUX21L U20802 ( .A(n3794), .B(n3795), .S(n4266), .Z(n3797) );
  ND4 U20803 ( .A(n4002), .B(n4001), .C(n4000), .D(n3999), .Z(n857) );
  ND4 U20804 ( .A(n855), .B(n4293), .C(n4231), .D(n4315), .Z(n3999) );
  MUX21L U20805 ( .A(n3993), .B(n3994), .S(n4339), .Z(n4002) );
  MUX21L U20806 ( .A(n3995), .B(n3996), .S(n4293), .Z(n4001) );
  AN3 U20807 ( .A(n856), .B(n4228), .C(n4332), .Z(n3995) );
  ND2 U20808 ( .A(n3546), .B(n3545), .Z(n856) );
  ND2 U20809 ( .A(n5247), .B(n4574), .Z(n3545) );
  EO U20810 ( .A(n4901), .B(n4574), .Z(n3546) );
  ND3 U20811 ( .A(n837), .B(n4315), .C(n4282), .Z(n4017) );
  ND2 U20812 ( .A(n3635), .B(n4410), .Z(n837) );
  EO U20813 ( .A(n5227), .B(n4938), .Z(n3635) );
  MUX41 U20814 ( .D0(n901), .D1(n884), .D2(n892), .D3(n879), .A(n4210), .B(
        n4218), .Z(N223) );
  AO3 U20815 ( .A(n4246), .B(n3724), .C(n3723), .D(n3722), .Z(n879) );
  MUX41 U20816 ( .D0(n857), .D1(n847), .D2(n850), .D3(n422), .A(n4209), .B(
        n4218), .Z(N221) );
  AO7 U20817 ( .A(n4324), .B(n3814), .C(n4243), .Z(n847) );
  ND4 U20818 ( .A(n3908), .B(n3907), .C(n3906), .D(n3905), .Z(n850) );
  MUX21L U20819 ( .A(n4005), .B(n4006), .S(n4340), .Z(n4009) );
  NR2 U20820 ( .A(n4261), .B(n4287), .Z(n4006) );
  NR3 U20821 ( .A(n4261), .B(n4293), .C(n417), .Z(n4005) );
  MUX21L U20822 ( .A(n4003), .B(n4004), .S(n4340), .Z(n4010) );
  NR2 U20823 ( .A(n4261), .B(n4186), .Z(n4004) );
  AN3 U20824 ( .A(n843), .B(n4287), .C(n4251), .Z(n4003) );
  MUX21L U20825 ( .A(n4016), .B(n4315), .S(n4260), .Z(n4019) );
  ND2 U20826 ( .A(n3474), .B(n3473), .Z(n836) );
  ND2 U20827 ( .A(n5244), .B(n4569), .Z(n3474) );
  MUX21L U20828 ( .A(n3704), .B(n3703), .S(n4267), .Z(n3706) );
  AN3 U20829 ( .A(n1059), .B(n4279), .C(n4331), .Z(n3703) );
  NR3 U20830 ( .A(n414), .B(n4352), .C(n4296), .Z(n3704) );
  ND2 U20831 ( .A(n2105), .B(n2104), .Z(n1059) );
  MUX21L U20832 ( .A(n3998), .B(n3997), .S(n4293), .Z(n4000) );
  AN3 U20833 ( .A(n854), .B(n4227), .C(n4332), .Z(n3997) );
  NR3 U20834 ( .A(n4261), .B(n4340), .C(n415), .Z(n3998) );
  AO4 U20835 ( .A(n4936), .B(n4604), .C(n5258), .D(n4604), .Z(n854) );
  ND2 U20836 ( .A(n3911), .B(n3910), .Z(N219) );
  ND2 U20837 ( .A(n834), .B(n4208), .Z(n3910) );
  MUX21L U20838 ( .A(n3909), .B(n4208), .S(n4222), .Z(n3911) );
  AO7 U20839 ( .A(n4324), .B(n3816), .C(n4242), .Z(n834) );
  NR2 U20840 ( .A(n3727), .B(n3726), .Z(n3729) );
  NR2 U20841 ( .A(n4267), .B(n4327), .Z(n3727) );
  NR2 U20842 ( .A(n4267), .B(n845), .Z(n3726) );
  ND4 U20843 ( .A(n4138), .B(n4137), .C(n4136), .D(n4135), .Z(n1039) );
  MUX21L U20844 ( .A(n4130), .B(n4129), .S(n4257), .Z(n4138) );
  AO2 U20845 ( .A(n4128), .B(n4230), .C(n4127), .D(n1037), .Z(n4136) );
  MUX21L U20846 ( .A(n4132), .B(n4131), .S(n4259), .Z(n4137) );
  ND4 U20847 ( .A(n3826), .B(n3825), .C(n3824), .D(n3823), .Z(n1009) );
  ND4 U20848 ( .A(n1005), .B(n4291), .C(n4265), .D(n4323), .Z(n3823) );
  MUX21L U20849 ( .A(n3817), .B(n3818), .S(n4353), .Z(n3826) );
  MUX21L U20850 ( .A(n3821), .B(n3822), .S(n4265), .Z(n3824) );
  ND4 U20851 ( .A(n3718), .B(n3717), .C(n3716), .D(n3715), .Z(n906) );
  ND4 U20852 ( .A(n4579), .B(n4296), .C(n4246), .D(n4327), .Z(n3715) );
  MUX21L U20853 ( .A(n3709), .B(n3710), .S(n4352), .Z(n3718) );
  MUX21L U20854 ( .A(n3711), .B(n3712), .S(n4352), .Z(n3717) );
  ND4 U20855 ( .A(n3899), .B(n3898), .C(n3897), .D(n3896), .Z(n867) );
  MUX21L U20856 ( .A(n3892), .B(n3893), .S(n4291), .Z(n3898) );
  ND3 U20857 ( .A(n866), .B(n4321), .C(n4279), .Z(n3896) );
  MUX21L U20858 ( .A(n3894), .B(n3895), .S(n4264), .Z(n3897) );
  AN3 U20859 ( .A(n1060), .B(n4246), .C(n4289), .Z(n3702) );
  ND2 U20860 ( .A(n2216), .B(n2215), .Z(n1060) );
  ND2 U20861 ( .A(n2212), .B(n5275), .Z(n2215) );
  MUX21L U20862 ( .A(n2213), .B(n2214), .S(n5275), .Z(n2216) );
  AN3 U20863 ( .A(n1036), .B(n4321), .C(n4290), .Z(n4129) );
  MUX21L U20864 ( .A(n2400), .B(n5265), .S(n4637), .Z(n1036) );
  ND2 U20865 ( .A(n5265), .B(n4883), .Z(n2400) );
  AN3 U20866 ( .A(n1007), .B(n4227), .C(n4290), .Z(n3817) );
  EO U20867 ( .A(n4903), .B(n4622), .Z(n1007) );
  AN3 U20868 ( .A(n905), .B(n4246), .C(n4289), .Z(n3712) );
  AO4 U20869 ( .A(n4967), .B(n4597), .C(n5275), .D(n4597), .Z(n905) );
  AN3 U20870 ( .A(n853), .B(n4287), .C(n4251), .Z(n3993) );
  ND2 U20871 ( .A(n3331), .B(n4489), .Z(n853) );
  ND2 U20872 ( .A(n5256), .B(n4934), .Z(n3331) );
  ND3 U20873 ( .A(n844), .B(n4232), .C(n4293), .Z(n4008) );
  ND2 U20874 ( .A(n3472), .B(n3471), .Z(n844) );
  ND2 U20875 ( .A(n5244), .B(n4569), .Z(n3472) );
  ND2 U20876 ( .A(n4920), .B(n4569), .Z(n3471) );
  ND3 U20877 ( .A(n3766), .B(n3765), .C(n3764), .Z(n829) );
  ND2 U20878 ( .A(n4244), .B(n4326), .Z(n3766) );
  ND2 U20879 ( .A(n4245), .B(n4285), .Z(n3764) );
  ND2 U20880 ( .A(n828), .B(n4244), .Z(n3765) );
  MUX21L U20881 ( .A(n4052), .B(n4053), .S(n4341), .Z(n4057) );
  AN3 U20882 ( .A(n1030), .B(n4277), .C(n4252), .Z(n4052) );
  ND3 U20883 ( .A(n2219), .B(n2218), .C(n2217), .Z(n1031) );
  MUX21L U20884 ( .A(n4054), .B(n4055), .S(n4259), .Z(n4056) );
  AN3 U20885 ( .A(n1033), .B(n4277), .C(n4333), .Z(n4054) );
  AO4 U20886 ( .A(n4912), .B(n4601), .C(n5272), .D(n4601), .Z(n1029) );
  MUX21L U20887 ( .A(n3819), .B(n3820), .S(n4291), .Z(n3825) );
  AN3 U20888 ( .A(n1008), .B(n4227), .C(n4330), .Z(n3819) );
  AN3 U20889 ( .A(n4330), .B(n4251), .C(n1004), .Z(n3820) );
  ND2 U20890 ( .A(n4970), .B(n4625), .Z(n1008) );
  MUX21L U20891 ( .A(n3714), .B(n3713), .S(n4267), .Z(n3716) );
  AN3 U20892 ( .A(n903), .B(n4278), .C(n4331), .Z(n3713) );
  NR3 U20893 ( .A(n421), .B(n4352), .C(n4296), .Z(n3714) );
  NR3 U20894 ( .A(n4601), .B(n5272), .C(n4912), .Z(n903) );
  MUX21L U20895 ( .A(n3719), .B(n3720), .S(n4296), .Z(n3723) );
  AN3 U20896 ( .A(n877), .B(n4310), .C(n4252), .Z(n3720) );
  NR2 U20897 ( .A(n4267), .B(n766), .Z(n3719) );
  NR3 U20898 ( .A(n4626), .B(n5270), .C(n4909), .Z(n877) );
  MUX21L U20899 ( .A(n3890), .B(n3891), .S(n4264), .Z(n3899) );
  AN3 U20900 ( .A(n864), .B(n4321), .C(n4288), .Z(n3890) );
  NR2 U20901 ( .A(n4291), .B(n4192), .Z(n3891) );
  AO4 U20902 ( .A(n4945), .B(n4552), .C(n5237), .D(n4552), .Z(n864) );
  MUX21L U20903 ( .A(n3904), .B(n4321), .S(n4264), .Z(n3905) );
  AN3 U20904 ( .A(n4290), .B(n767), .C(n4332), .Z(n3904) );
  ND2 U20905 ( .A(n3756), .B(n3755), .Z(N218) );
  MUX21L U20906 ( .A(n3754), .B(n4202), .S(n4222), .Z(n3756) );
  ND2 U20907 ( .A(n832), .B(n4202), .Z(n3755) );
  ND2 U20908 ( .A(n849), .B(n4280), .Z(n3907) );
  NR3 U20909 ( .A(n4555), .B(n5231), .C(n4942), .Z(n849) );
  AO2 U20910 ( .A(n848), .B(n4263), .C(n4263), .D(n4284), .Z(n3906) );
  NR3 U20911 ( .A(n4559), .B(n5278), .C(n4904), .Z(n848) );
  AN3 U20912 ( .A(n5221), .B(n4277), .C(n4334), .Z(n4131) );
  AN3 U20913 ( .A(n852), .B(n4287), .C(n4251), .Z(n3994) );
  AO7 U20914 ( .A(n5252), .B(n4952), .C(n4612), .Z(n852) );
  MUX21L U20915 ( .A(n3725), .B(n4246), .S(n4296), .Z(n3728) );
  AN3 U20916 ( .A(n858), .B(n4310), .C(n4252), .Z(n3725) );
  NR2 U20917 ( .A(n4913), .B(n4599), .Z(n858) );
  ND2 U20918 ( .A(n840), .B(n4238), .Z(n3879) );
  ND2 U20919 ( .A(n4947), .B(n4548), .Z(n840) );
  AO7 U20920 ( .A(n4324), .B(n3815), .C(n4242), .Z(n839) );
  ND2 U20921 ( .A(n4291), .B(n838), .Z(n3815) );
  ND2 U20922 ( .A(n2589), .B(n4520), .Z(n838) );
  ND2 U20923 ( .A(n5290), .B(n4973), .Z(n2589) );
  MUX21L U20924 ( .A(n4050), .B(n4051), .S(n4261), .Z(n4058) );
  AN3 U20925 ( .A(n1032), .B(n4314), .C(n4289), .Z(n4050) );
  ND2 U20926 ( .A(n4453), .B(n4855), .Z(n1028) );
  MUX21L U20927 ( .A(n3759), .B(n4283), .S(n4266), .Z(n3762) );
  AN3 U20928 ( .A(n4331), .B(n860), .C(n4289), .Z(n3759) );
  ND2 U20929 ( .A(n2587), .B(n4521), .Z(n860) );
  ND2 U20930 ( .A(n5290), .B(n4973), .Z(n2587) );
  ND3 U20931 ( .A(n4960), .B(n4632), .C(n5261), .Z(n845) );
  AN3 U20932 ( .A(n4900), .B(n4279), .C(n4252), .Z(n3699) );
  AN3 U20933 ( .A(n4734), .B(n4278), .C(n4251), .Z(n3818) );
  MUX21L U20934 ( .A(n3721), .B(n4285), .S(n4352), .Z(n3722) );
  AN3 U20935 ( .A(n4363), .B(n4225), .C(n4289), .Z(n3721) );
  AO7 U20936 ( .A(n4186), .B(n3982), .C(n3981), .Z(n827) );
  ND2 U20937 ( .A(n4231), .B(n4316), .Z(n3982) );
  IVP U20938 ( .A(n4276), .Z(n4298) );
  IVP U20939 ( .A(n4311), .Z(n4342) );
  AN3 U20940 ( .A(n904), .B(n4284), .C(n4252), .Z(n3709) );
  ND2 U20941 ( .A(n4462), .B(n4861), .Z(n904) );
  AN3 U20942 ( .A(n883), .B(n4227), .C(n4331), .Z(n3792) );
  ND3 U20943 ( .A(n4757), .B(n5204), .C(n4509), .Z(n883) );
  AN3 U20944 ( .A(n865), .B(n4228), .C(n4331), .Z(n3892) );
  ND3 U20945 ( .A(n4822), .B(n5096), .C(n4381), .Z(n865) );
  NR2 U20946 ( .A(n4353), .B(n4286), .Z(n3795) );
  ND2 U20947 ( .A(n878), .B(n4285), .Z(n3724) );
  ND2 U20948 ( .A(n4462), .B(n4862), .Z(n878) );
  ND2 U20949 ( .A(n4239), .B(n4280), .Z(n3878) );
  ND2 U20950 ( .A(n4239), .B(n4321), .Z(n3880) );
  ND2 U20951 ( .A(n4230), .B(n4283), .Z(n3981) );
  ND2 U20952 ( .A(n4279), .B(n4320), .Z(n3908) );
  IVP U20953 ( .A(LogIn2[44]), .Z(n4276) );
  IVP U20954 ( .A(n5296), .Z(n5301) );
  IVP U20955 ( .A(n5322), .Z(n5306) );
  IVP U20956 ( .A(n5297), .Z(n5298) );
  IVP U20957 ( .A(n5297), .Z(n5300) );
  IVP U20958 ( .A(n5296), .Z(n5303) );
  IVP U20959 ( .A(n5297), .Z(n5299) );
  IVP U20960 ( .A(n5296), .Z(n5302) );
  IVP U20961 ( .A(LogIn2[40]), .Z(n5305) );
  IVP U20962 ( .A(n5307), .Z(n5304) );
  IVP U20963 ( .A(n4308), .Z(n4277) );
  IVP U20964 ( .A(n4308), .Z(n4286) );
  IVP U20965 ( .A(n4307), .Z(n4279) );
  IVP U20966 ( .A(n4307), .Z(n4282) );
  IVP U20967 ( .A(n4296), .Z(n4278) );
  IVP U20968 ( .A(n4307), .Z(n4283) );
  IVP U20969 ( .A(n4307), .Z(n4284) );
  IVP U20970 ( .A(n4308), .Z(n4285) );
  IVP U20971 ( .A(n4308), .Z(n4287) );
  IVP U20972 ( .A(LogIn2[44]), .Z(n4280) );
  IVP U20973 ( .A(LogIn2[47]), .Z(n4204) );
  IVP U20974 ( .A(LogIn2[44]), .Z(n4281) );
  IVP U20975 ( .A(LogIn2[47]), .Z(n4207) );
  IVP U20976 ( .A(LogIn2[47]), .Z(n4203) );
  IVP U20977 ( .A(LogIn2[47]), .Z(n4206) );
  IVP U20978 ( .A(LogIn2[47]), .Z(n4202) );
  IVP U20979 ( .A(LogIn2[47]), .Z(n4205) );
  IVP U20980 ( .A(n5368), .Z(n5367) );
  IVP U20981 ( .A(n5368), .Z(n5366) );
  IVP U20982 ( .A(n5368), .Z(n5365) );
  IVP U20983 ( .A(n5370), .Z(n5363) );
  IVP U20984 ( .A(n5369), .Z(n5364) );
  IVP U20985 ( .A(n5371), .Z(n5362) );
  IVP U20986 ( .A(n5305), .Z(n5296) );
  IVP U20987 ( .A(n5306), .Z(n5297) );
  IVP U20988 ( .A(n4280), .Z(n4308) );
  IVP U20989 ( .A(n4281), .Z(n4307) );
  AO5 U20990 ( .A(n793), .B(n794), .C(n5379), .Z(n792) );
  FA1A U20991 ( .A(Term31[26]), .B(Term11[114]), .CI(
        \add_1_root_sub_1_root_add_55_2/carry[2] ), .CO(
        \add_1_root_sub_1_root_add_55_2/carry[3] ), .S(N280) );
  FA1A U20992 ( .A(Term31[24]), .B(Term11[112]), .CI(FractionBit[23]), .CO(
        \add_1_root_sub_1_root_add_55_2/carry[1] ), .S(N278) );
  FA1A U20993 ( .A(Term31[25]), .B(Term11[113]), .CI(
        \add_1_root_sub_1_root_add_55_2/carry[1] ), .CO(
        \add_1_root_sub_1_root_add_55_2/carry[2] ), .S(N279) );
  IV U20994 ( .A(n807), .Z(n808) );
  IV U20995 ( .A(n809), .Z(n810) );
  IV U20996 ( .A(n811), .Z(n812) );
  IV U20997 ( .A(n821), .Z(n822) );
  IV U20998 ( .A(n823), .Z(n824) );
  MUX81P U20999 ( .D0(n875), .D1(n871), .D2(n873), .D3(n869), .D4(n874), .D5(
        n870), .D6(n872), .D7(n868), .A(n4250), .B(n4306), .C(n4336), .Z(n876)
         );
  MUX81P U21000 ( .D0(n891), .D1(n4399), .D2(n889), .D3(n886), .D4(n890), .D5(
        n887), .D6(n888), .D7(n885), .A(n4254), .B(n4302), .C(n4353), .Z(n892)
         );
  MUX81P U21001 ( .D0(n900), .D1(n896), .D2(n898), .D3(n894), .D4(n899), .D5(
        n895), .D6(n897), .D7(n893), .A(n4254), .B(n4297), .C(n4341), .Z(n901)
         );
  MUX81P U21002 ( .D0(n914), .D1(n910), .D2(n912), .D3(n908), .D4(n913), .D5(
        n909), .D6(n911), .D7(n907), .A(n4254), .B(n4298), .C(n4341), .Z(n915)
         );
  MUX81P U21003 ( .D0(n923), .D1(n919), .D2(n921), .D3(n917), .D4(n922), .D5(
        n918), .D6(n920), .D7(n916), .A(n4254), .B(n4298), .C(n4341), .Z(n924)
         );
  MUX81P U21004 ( .D0(n931), .D1(n5269), .D2(n929), .D3(n926), .D4(n930), .D5(
        n927), .D6(n928), .D7(n925), .A(n4254), .B(n4298), .C(n4341), .Z(n932)
         );
  MUX81P U21005 ( .D0(n939), .D1(n935), .D2(n937), .D3(n933), .D4(n938), .D5(
        n934), .D6(n936), .D7(n4446), .A(n4254), .B(n4298), .C(n4341), .Z(n940) );
  MUX81P U21006 ( .D0(n948), .D1(n944), .D2(n946), .D3(n942), .D4(n947), .D5(
        n943), .D6(n945), .D7(n941), .A(n4254), .B(n4298), .C(n4342), .Z(n949)
         );
  MUX81P U21007 ( .D0(n5269), .D1(n953), .D2(n955), .D3(n951), .D4(n956), .D5(
        n952), .D6(n954), .D7(n950), .A(n4254), .B(n4298), .C(n4342), .Z(n957)
         );
  MUX81P U21008 ( .D0(n963), .D1(n767), .D2(n961), .D3(n958), .D4(n962), .D5(
        n959), .D6(n960), .D7(n5269), .A(n4254), .B(n4298), .C(n4342), .Z(n964) );
  MUX81P U21009 ( .D0(n971), .D1(n967), .D2(n969), .D3(n965), .D4(n970), .D5(
        n966), .D6(n968), .D7(n4858), .A(n4254), .B(n4298), .C(n4342), .Z(n972) );
  MUX81P U21010 ( .D0(n5268), .D1(n976), .D2(n978), .D3(n974), .D4(n979), .D5(
        n975), .D6(n977), .D7(n973), .A(n4254), .B(n4298), .C(n4342), .Z(n980)
         );
  MUX81P U21011 ( .D0(n767), .D1(n983), .D2(n985), .D3(n981), .D4(n986), .D5(
        n982), .D6(n984), .D7(n5268), .A(n4254), .B(n4298), .C(n4342), .Z(n987) );
  MUX81P U21012 ( .D0(n995), .D1(n991), .D2(n993), .D3(n989), .D4(n994), .D5(
        n990), .D6(n992), .D7(n988), .A(n4254), .B(n4298), .C(n4342), .Z(n996)
         );
  MUX81P U21013 ( .D0(n1002), .D1(n998), .D2(n1000), .D3(n997), .D4(n1001), 
        .D5(n5259), .D6(n999), .D7(n5176), .A(n4254), .B(n4298), .C(n4342), 
        .Z(n1003) );
  MUX81P U21014 ( .D0(n1017), .D1(n1013), .D2(n1015), .D3(n1011), .D4(n1016), 
        .D5(n1012), .D6(n1014), .D7(n1010), .A(n4255), .B(n4299), .C(n4342), 
        .Z(n1018) );
  MUX81P U21015 ( .D0(n1026), .D1(n1022), .D2(n1024), .D3(n1020), .D4(n1025), 
        .D5(n1021), .D6(n1023), .D7(n1019), .A(n4255), .B(n4299), .C(n4342), 
        .Z(n1027) );
  MUX81P U21016 ( .D0(n1047), .D1(n1043), .D2(n1045), .D3(n1041), .D4(n1046), 
        .D5(n1042), .D6(n1044), .D7(n1040), .A(n4255), .B(n4299), .C(n4342), 
        .Z(n1048) );
  MUX81P U21017 ( .D0(n1056), .D1(n1052), .D2(n1054), .D3(n1050), .D4(n1055), 
        .D5(n1051), .D6(n1053), .D7(n1049), .A(n4255), .B(n4299), .C(n4342), 
        .Z(n1057) );
  MUX81P U21018 ( .D0(n1069), .D1(n1066), .D2(n5268), .D3(n1064), .D4(n1068), 
        .D5(n1065), .D6(n1067), .D7(n1063), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1070) );
  MUX81P U21019 ( .D0(n1077), .D1(n1074), .D2(n1076), .D3(n1072), .D4(n781), 
        .D5(n1073), .D6(n1075), .D7(n1071), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1078) );
  MUX81P U21020 ( .D0(n1086), .D1(n1082), .D2(n1084), .D3(n1080), .D4(n1085), 
        .D5(n1081), .D6(n1083), .D7(n1079), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1087) );
  MUX81P U21021 ( .D0(n1118), .D1(n1114), .D2(n1116), .D3(n1112), .D4(n1117), 
        .D5(n1113), .D6(n1115), .D7(n1111), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1119) );
  MUX81P U21022 ( .D0(n1135), .D1(n1131), .D2(n1133), .D3(n1129), .D4(n1134), 
        .D5(n1130), .D6(n1132), .D7(n1128), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1136) );
  MUX81P U21023 ( .D0(n1156), .D1(n1152), .D2(n1154), .D3(n1151), .D4(n1155), 
        .D5(n5269), .D6(n1153), .D7(n1150), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1157) );
  MUX81P U21024 ( .D0(n4507), .D1(n4475), .D2(n1164), .D3(n1162), .D4(n1165), 
        .D5(n1163), .D6(n754), .D7(n1161), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1166) );
  MUX81P U21025 ( .D0(n1172), .D1(n4934), .D2(n1170), .D3(n1167), .D4(n1171), 
        .D5(n1168), .D6(n1169), .D7(n4502), .A(n4255), .B(n4299), .C(n4343), 
        .Z(n1173) );
  MUX81P U21026 ( .D0(n1180), .D1(n1176), .D2(n1178), .D3(n4934), .D4(n1179), 
        .D5(n1175), .D6(n1177), .D7(n1174), .A(n4255), .B(n4300), .C(n4343), 
        .Z(n1181) );
  MUX81P U21027 ( .D0(n4755), .D1(n1190), .D2(n1192), .D3(n1188), .D4(n1193), 
        .D5(n1189), .D6(n1191), .D7(n1187), .A(n4255), .B(n4300), .C(n4343), 
        .Z(n1194) );
  MUX81P U21028 ( .D0(n1200), .D1(n1197), .D2(n1198), .D3(n1195), .D4(n1199), 
        .D5(n1196), .D6(n5269), .D7(n4749), .A(n4255), .B(n4300), .C(n4343), 
        .Z(n1201) );
  MUX81P U21029 ( .D0(n1207), .D1(n1203), .D2(n1205), .D3(n5269), .D4(n1206), 
        .D5(n776), .D6(n1204), .D7(n1202), .A(n4255), .B(n4300), .C(n4343), 
        .Z(n1208) );
  MUX81P U21030 ( .D0(n1215), .D1(n1211), .D2(n1213), .D3(n1209), .D4(n1214), 
        .D5(n1210), .D6(n1212), .D7(n4445), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1216) );
  MUX81P U21031 ( .D0(n5177), .D1(n1219), .D2(n1221), .D3(n4976), .D4(n1222), 
        .D5(n1218), .D6(n1220), .D7(n1217), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1223) );
  MUX81P U21032 ( .D0(n1236), .D1(n1232), .D2(n1234), .D3(n1231), .D4(n1235), 
        .D5(n774), .D6(n1233), .D7(n1230), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1237) );
  MUX81P U21033 ( .D0(n1244), .D1(n1240), .D2(n1242), .D3(n1238), .D4(n1243), 
        .D5(n1239), .D6(n1241), .D7(n4859), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1245) );
  MUX81P U21034 ( .D0(n1264), .D1(n1261), .D2(n773), .D3(n1259), .D4(n1263), 
        .D5(n1260), .D6(n1262), .D7(n1258), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1265) );
  MUX81P U21035 ( .D0(n1272), .D1(n1268), .D2(n1270), .D3(n1266), .D4(n1271), 
        .D5(n1267), .D6(n1269), .D7(n5175), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1273) );
  MUX81P U21036 ( .D0(n1284), .D1(n1281), .D2(n1282), .D3(n1279), .D4(n1283), 
        .D5(n1280), .D6(n772), .D7(n1278), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1285) );
  MUX81P U21037 ( .D0(n1293), .D1(n1289), .D2(n1291), .D3(n1287), .D4(n1292), 
        .D5(n1288), .D6(n1290), .D7(n1286), .A(n4255), .B(n4300), .C(n4344), 
        .Z(n1294) );
  MUX81P U21038 ( .D0(n1316), .D1(n1312), .D2(n1314), .D3(n1310), .D4(n1315), 
        .D5(n1311), .D6(n1313), .D7(n1309), .A(n4256), .B(n4301), .C(n4344), 
        .Z(n1317) );
  MUX81P U21039 ( .D0(n4772), .D1(n1320), .D2(n1321), .D3(n4954), .D4(n1322), 
        .D5(n1319), .D6(n4591), .D7(n1318), .A(n4256), .B(n4301), .C(n4344), 
        .Z(n1323) );
  MUX81P U21040 ( .D0(n1337), .D1(n1333), .D2(n1335), .D3(n1331), .D4(n1336), 
        .D5(n1332), .D6(n1334), .D7(n1330), .A(n4256), .B(n4301), .C(n4344), 
        .Z(n1338) );
  MUX81P U21041 ( .D0(n1345), .D1(n1342), .D2(n1343), .D3(n1340), .D4(n1344), 
        .D5(n1341), .D6(n5268), .D7(n1339), .A(n4256), .B(n4301), .C(n4344), 
        .Z(n1346) );
  MUX81P U21042 ( .D0(n1353), .D1(n1350), .D2(n1352), .D3(n1348), .D4(n770), 
        .D5(n1349), .D6(n1351), .D7(n1347), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1354) );
  MUX81P U21043 ( .D0(n1362), .D1(n1358), .D2(n1360), .D3(n1356), .D4(n1361), 
        .D5(n1357), .D6(n1359), .D7(n1355), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1363) );
  MUX81P U21044 ( .D0(n1371), .D1(n1367), .D2(n1369), .D3(n1365), .D4(n1370), 
        .D5(n1366), .D6(n1368), .D7(n1364), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1372) );
  MUX81P U21045 ( .D0(n1380), .D1(n1376), .D2(n1378), .D3(n1374), .D4(n1379), 
        .D5(n1375), .D6(n1377), .D7(n1373), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1381) );
  MUX81P U21046 ( .D0(n1396), .D1(n1392), .D2(n1394), .D3(n1390), .D4(n1395), 
        .D5(n1391), .D6(n1393), .D7(n1389), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1397) );
  MUX81P U21047 ( .D0(n1405), .D1(n1401), .D2(n1403), .D3(n1399), .D4(n1404), 
        .D5(n1400), .D6(n1402), .D7(n1398), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1406) );
  MUX81P U21048 ( .D0(n1417), .D1(n1413), .D2(n1415), .D3(n1412), .D4(n1416), 
        .D5(n769), .D6(n1414), .D7(n1411), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1418) );
  MUX81P U21049 ( .D0(n1425), .D1(n1421), .D2(n1423), .D3(n1419), .D4(n1424), 
        .D5(n1420), .D6(n1422), .D7(n4859), .A(n4256), .B(n4301), .C(n4345), 
        .Z(n1426) );
  MUX81P U21050 ( .D0(n1434), .D1(n1430), .D2(n1432), .D3(n1428), .D4(n1433), 
        .D5(n1429), .D6(n1431), .D7(n1427), .A(n4256), .B(n4302), .C(n4345), 
        .Z(n1435) );
  MUX81P U21051 ( .D0(n1442), .D1(n1439), .D2(n759), .D3(n1437), .D4(n1441), 
        .D5(n1438), .D6(n1440), .D7(n1436), .A(n4256), .B(n4302), .C(n4345), 
        .Z(n1443) );
  MUX81P U21052 ( .D0(n1451), .D1(n1447), .D2(n1449), .D3(n1445), .D4(n1450), 
        .D5(n1446), .D6(n1448), .D7(n1444), .A(n4256), .B(n4302), .C(n4345), 
        .Z(n1452) );
  MUX81P U21053 ( .D0(n1460), .D1(n1456), .D2(n1458), .D3(n1454), .D4(n1459), 
        .D5(n1455), .D6(n1457), .D7(n1453), .A(n4256), .B(n4302), .C(n4345), 
        .Z(n1461) );
  MUX81P U21054 ( .D0(n1476), .D1(n1472), .D2(n1474), .D3(n1470), .D4(n1475), 
        .D5(n1471), .D6(n1473), .D7(n1469), .A(n4257), .B(n4302), .C(n4346), 
        .Z(n1477) );
  MUX81P U21055 ( .D0(n1485), .D1(n1481), .D2(n1483), .D3(n1479), .D4(n1484), 
        .D5(n1480), .D6(n1482), .D7(n1478), .A(n4256), .B(n4302), .C(n4346), 
        .Z(n1486) );
  MUX81P U21056 ( .D0(n1526), .D1(n1522), .D2(n1524), .D3(n4588), .D4(n1525), 
        .D5(n1521), .D6(n1523), .D7(n1520), .A(n4257), .B(n4302), .C(n4346), 
        .Z(n1527) );
  MUX81P U21057 ( .D0(n1539), .D1(n1535), .D2(n1537), .D3(n1533), .D4(n1538), 
        .D5(n1534), .D6(n1536), .D7(n1532), .A(n4256), .B(n4302), .C(n4346), 
        .Z(n1540) );
  MUX81P U21058 ( .D0(n1556), .D1(n1552), .D2(n1554), .D3(n1550), .D4(n1555), 
        .D5(n1551), .D6(n1553), .D7(n1549), .A(n4256), .B(n4302), .C(n4346), 
        .Z(n1557) );
  MUX81P U21059 ( .D0(n1568), .D1(n1564), .D2(n1566), .D3(n1562), .D4(n1567), 
        .D5(n1563), .D6(n1565), .D7(n1561), .A(n4257), .B(n4302), .C(n4346), 
        .Z(n1569) );
  MUX81P U21060 ( .D0(n1576), .D1(n779), .D2(n1574), .D3(n1571), .D4(n1575), 
        .D5(n1572), .D6(n1573), .D7(n1570), .A(n4257), .B(n4302), .C(n4346), 
        .Z(n1577) );
  MUX81P U21061 ( .D0(n1594), .D1(n1590), .D2(n1592), .D3(n1588), .D4(n1593), 
        .D5(n1589), .D6(n1591), .D7(n1587), .A(n4256), .B(n4303), .C(n4346), 
        .Z(n1595) );
  MUX81P U21062 ( .D0(n1602), .D1(n778), .D2(n1600), .D3(n1597), .D4(n1601), 
        .D5(n1598), .D6(n1599), .D7(n1596), .A(n4257), .B(n4303), .C(n4346), 
        .Z(n1603) );
  MUX81P U21063 ( .D0(n4756), .D1(n1612), .D2(n1614), .D3(n1610), .D4(n1615), 
        .D5(n1611), .D6(n1613), .D7(n1609), .A(n4257), .B(n4303), .C(n4346), 
        .Z(n1616) );
  MUX81P U21064 ( .D0(n1624), .D1(n1620), .D2(n1622), .D3(n1618), .D4(n1623), 
        .D5(n1619), .D6(n1621), .D7(n1617), .A(n4256), .B(n4303), .C(n4346), 
        .Z(n1625) );
  MUX81P U21065 ( .D0(n1633), .D1(n1629), .D2(n1631), .D3(n1627), .D4(n1632), 
        .D5(n1628), .D6(n1630), .D7(n1626), .A(n4257), .B(n4303), .C(n4346), 
        .Z(n1634) );
  MUX81P U21066 ( .D0(n1647), .D1(n4904), .D2(n1645), .D3(n1642), .D4(n1646), 
        .D5(n1643), .D6(n1644), .D7(n1641), .A(n4257), .B(n4303), .C(n4347), 
        .Z(n1648) );
  MUX81P U21067 ( .D0(n1656), .D1(n1652), .D2(n1654), .D3(n1650), .D4(n1655), 
        .D5(n1651), .D6(n1653), .D7(n1649), .A(n4256), .B(n4303), .C(n4347), 
        .Z(n1657) );
  MUX81P U21068 ( .D0(n1665), .D1(n1661), .D2(n1663), .D3(n1659), .D4(n1664), 
        .D5(n1660), .D6(n1662), .D7(n1658), .A(n4257), .B(n4303), .C(n4347), 
        .Z(n1666) );
  MUX81P U21069 ( .D0(n1673), .D1(n1669), .D2(n1671), .D3(n1667), .D4(n1672), 
        .D5(n1668), .D6(n1670), .D7(n4444), .A(n4257), .B(n4303), .C(n4347), 
        .Z(n1674) );
  MUX81P U21070 ( .D0(n1680), .D1(n5176), .D2(n1679), .D3(n1676), .D4(n4969), 
        .D5(n1677), .D6(n1678), .D7(n1675), .A(n4257), .B(n4303), .C(n4347), 
        .Z(n1681) );
  MUX81P U21071 ( .D0(n777), .D1(n1685), .D2(n1687), .D3(n1683), .D4(n1688), 
        .D5(n1684), .D6(n1686), .D7(n1682), .A(n4257), .B(n4303), .C(n4347), 
        .Z(n1689) );
  MUX81P U21072 ( .D0(n1701), .D1(n1698), .D2(n1700), .D3(n1696), .D4(n5268), 
        .D5(n1697), .D6(n1699), .D7(n4860), .A(n4257), .B(n4303), .C(n4347), 
        .Z(n1702) );
  MUX81P U21073 ( .D0(n1709), .D1(n4614), .D2(n1707), .D3(n1704), .D4(n1708), 
        .D5(n1705), .D6(n1706), .D7(n1703), .A(n4257), .B(n4304), .C(n4347), 
        .Z(n1710) );
  MUX81P U21074 ( .D0(n1717), .D1(n1713), .D2(n1715), .D3(n1711), .D4(n1716), 
        .D5(n1712), .D6(n1714), .D7(n775), .A(n4257), .B(n4304), .C(n4347), 
        .Z(n1718) );
  MUX81P U21075 ( .D0(n1725), .D1(n1721), .D2(n1723), .D3(n1719), .D4(n1724), 
        .D5(n1720), .D6(n1722), .D7(n5220), .A(n4257), .B(n4304), .C(n4347), 
        .Z(n1726) );
  MUX81P U21076 ( .D0(n1739), .D1(n4474), .D2(n1737), .D3(n1734), .D4(n1738), 
        .D5(n1735), .D6(n1736), .D7(n1733), .A(n4257), .B(n4304), .C(n4347), 
        .Z(n1740) );
  MUX81P U21077 ( .D0(n1747), .D1(n3408), .D2(n1745), .D3(n1742), .D4(n1746), 
        .D5(n1743), .D6(n1744), .D7(n1741), .A(n4257), .B(n4304), .C(n4348), 
        .Z(n1748) );
  MUX81P U21078 ( .D0(n1756), .D1(n1752), .D2(n1754), .D3(n1750), .D4(n1755), 
        .D5(n1751), .D6(n1753), .D7(n1749), .A(n4257), .B(n4304), .C(n4348), 
        .Z(n1757) );
  MUX81P U21079 ( .D0(n1770), .D1(n1766), .D2(n1768), .D3(n1764), .D4(n1769), 
        .D5(n1765), .D6(n1767), .D7(n5268), .A(n4256), .B(n4304), .C(n4348), 
        .Z(n1771) );
  MUX81P U21080 ( .D0(n1779), .D1(n1775), .D2(n1777), .D3(n1773), .D4(n1778), 
        .D5(n1774), .D6(n1776), .D7(n1772), .A(n4257), .B(n4304), .C(n4348), 
        .Z(n1780) );
  MUX81P U21081 ( .D0(n1788), .D1(n1784), .D2(n1786), .D3(n1782), .D4(n1787), 
        .D5(n1783), .D6(n1785), .D7(n1781), .A(n4257), .B(n4304), .C(n4348), 
        .Z(n1789) );
  MUX81P U21082 ( .D0(n1796), .D1(n1793), .D2(n5176), .D3(n1791), .D4(n1795), 
        .D5(n1792), .D6(n1794), .D7(n1790), .A(n4256), .B(n4304), .C(n4348), 
        .Z(n1797) );
  MUX81P U21083 ( .D0(n1805), .D1(n1801), .D2(n1803), .D3(n1799), .D4(n1804), 
        .D5(n1800), .D6(n1802), .D7(n1798), .A(n4254), .B(n4304), .C(n4348), 
        .Z(n1806) );
  MUX81P U21084 ( .D0(n1813), .D1(n1809), .D2(n1811), .D3(n1808), .D4(n1812), 
        .D5(n2878), .D6(n1810), .D7(n1807), .A(n4254), .B(n4304), .C(n4348), 
        .Z(n1814) );
  MUX81P U21085 ( .D0(n1821), .D1(n4908), .D2(n1819), .D3(n1816), .D4(n1820), 
        .D5(n1817), .D6(n1818), .D7(n1815), .A(n4254), .B(n4305), .C(n4348), 
        .Z(n1822) );
  MUX81P U21086 ( .D0(n1829), .D1(n1825), .D2(n1827), .D3(n1823), .D4(n1828), 
        .D5(n1824), .D6(n1826), .D7(n771), .A(n4254), .B(n4305), .C(n4348), 
        .Z(n1830) );
  MUX81P U21087 ( .D0(n1837), .D1(n1834), .D2(n1836), .D3(n1832), .D4(n4895), 
        .D5(n1833), .D6(n1835), .D7(n1831), .A(n4254), .B(n4305), .C(n4348), 
        .Z(n1838) );
  MUX81P U21088 ( .D0(n1846), .D1(n1842), .D2(n1844), .D3(n1840), .D4(n1845), 
        .D5(n1841), .D6(n1843), .D7(n1839), .A(n4254), .B(n4305), .C(n4348), 
        .Z(n1847) );
  MUX81P U21089 ( .D0(n1855), .D1(n1851), .D2(n1853), .D3(n1849), .D4(n1854), 
        .D5(n1850), .D6(n1852), .D7(n1848), .A(n4254), .B(n4305), .C(n4349), 
        .Z(n1856) );
  MUX81P U21090 ( .D0(n1864), .D1(n1860), .D2(n1862), .D3(n1858), .D4(n1863), 
        .D5(n1859), .D6(n1861), .D7(n1857), .A(n4254), .B(n4305), .C(n4349), 
        .Z(n1865) );
  MUX81P U21091 ( .D0(n1880), .D1(n1876), .D2(n1878), .D3(n1874), .D4(n1879), 
        .D5(n1875), .D6(n1877), .D7(n1873), .A(n4254), .B(n4305), .C(n4349), 
        .Z(n1881) );
  MUX81P U21092 ( .D0(n1889), .D1(n1885), .D2(n1887), .D3(n1883), .D4(n1888), 
        .D5(n1884), .D6(n1886), .D7(n1882), .A(n4253), .B(n4305), .C(n4349), 
        .Z(n1890) );
  MUX81P U21093 ( .D0(n1898), .D1(n1894), .D2(n1896), .D3(n1892), .D4(n1897), 
        .D5(n1893), .D6(n1895), .D7(n1891), .A(n4253), .B(n4305), .C(n4349), 
        .Z(n1899) );
  MUX81P U21094 ( .D0(n1907), .D1(n1903), .D2(n1905), .D3(n1901), .D4(n1906), 
        .D5(n1902), .D6(n1904), .D7(n1900), .A(n4253), .B(n4305), .C(n4349), 
        .Z(n1908) );
  MUX81P U21095 ( .D0(n1916), .D1(n1912), .D2(n1914), .D3(n1910), .D4(n1915), 
        .D5(n1911), .D6(n1913), .D7(n1909), .A(n4253), .B(n4305), .C(n4349), 
        .Z(n1917) );
  MUX81P U21096 ( .D0(n1925), .D1(n1921), .D2(n1923), .D3(n1919), .D4(n1924), 
        .D5(n1920), .D6(n1922), .D7(n1918), .A(n4253), .B(n4305), .C(n4349), 
        .Z(n1926) );
  MUX81P U21097 ( .D0(n1934), .D1(n1930), .D2(n1932), .D3(n1928), .D4(n1933), 
        .D5(n1929), .D6(n1931), .D7(n1927), .A(n4253), .B(n4306), .C(n4349), 
        .Z(n1935) );
  MUX81P U21098 ( .D0(n1943), .D1(n1939), .D2(n1941), .D3(n1937), .D4(n1942), 
        .D5(n1938), .D6(n1940), .D7(n1936), .A(n4253), .B(n4306), .C(n4349), 
        .Z(n1944) );
  MUX81P U21099 ( .D0(n5155), .D1(n771), .D2(n753), .D3(n1945), .D4(n1948), 
        .D5(n1946), .D6(n1947), .D7(n2893), .A(n4253), .B(n4306), .C(n4349), 
        .Z(n1949) );
  MUX81P U21100 ( .D0(n1957), .D1(n1953), .D2(n1955), .D3(n1951), .D4(n1956), 
        .D5(n1952), .D6(n1954), .D7(n1950), .A(n4253), .B(n4306), .C(n4349), 
        .Z(n1958) );
  MUX81P U21101 ( .D0(n1966), .D1(n1962), .D2(n1964), .D3(n1960), .D4(n1965), 
        .D5(n1961), .D6(n1963), .D7(n1959), .A(n4253), .B(n4306), .C(n4350), 
        .Z(n1967) );
  MUX81P U21102 ( .D0(n1975), .D1(n1971), .D2(n1973), .D3(n1969), .D4(n1974), 
        .D5(n1970), .D6(n1972), .D7(n1968), .A(n4253), .B(n4306), .C(n4350), 
        .Z(n1976) );
  MUX81P U21103 ( .D0(n1990), .D1(n1986), .D2(n1988), .D3(n1984), .D4(n1989), 
        .D5(n1985), .D6(n1987), .D7(n1983), .A(n4253), .B(n4306), .C(n4350), 
        .Z(n1991) );
  MUX81P U21104 ( .D0(n1999), .D1(n1995), .D2(n1997), .D3(n1993), .D4(n1998), 
        .D5(n1994), .D6(n1996), .D7(n1992), .A(n4253), .B(n4306), .C(n4350), 
        .Z(n2000) );
  MUX81P U21105 ( .D0(n2008), .D1(n2004), .D2(n2006), .D3(n2002), .D4(n2007), 
        .D5(n2003), .D6(n2005), .D7(n2001), .A(n4253), .B(n4306), .C(n4350), 
        .Z(n2009) );
  MUX81P U21106 ( .D0(n2016), .D1(n2013), .D2(n2015), .D3(n2011), .D4(n768), 
        .D5(n2012), .D6(n2014), .D7(n2010), .A(n4253), .B(n4306), .C(n4350), 
        .Z(n2017) );
  MUX81P U21107 ( .D0(n2025), .D1(n2021), .D2(n2023), .D3(n2019), .D4(n2024), 
        .D5(n2020), .D6(n2022), .D7(n2018), .A(n4253), .B(n4306), .C(n4350), 
        .Z(n2026) );
  AN2P U21108 ( .A(n4546), .B(n5227), .Z(n2039) );
  AN2P U21109 ( .A(n4903), .B(n4546), .Z(n2075) );
  AN2P U21110 ( .A(n5228), .B(n4546), .Z(n2094) );
  AN2P U21111 ( .A(n5228), .B(n4546), .Z(n2098) );
  AN2P U21112 ( .A(n5228), .B(n4902), .Z(n2102) );
  AN2P U21113 ( .A(n5228), .B(n4901), .Z(n2109) );
  AN2P U21114 ( .A(n4901), .B(n4545), .Z(n2115) );
  AN2P U21115 ( .A(n5229), .B(n4900), .Z(n2141) );
  AN2P U21116 ( .A(n5229), .B(n4900), .Z(n2150) );
  AN2P U21117 ( .A(n5229), .B(n4900), .Z(n2153) );
  AN2P U21118 ( .A(n5229), .B(n4547), .Z(n2175) );
  AN2P U21119 ( .A(n5229), .B(n4544), .Z(n2179) );
  AN2P U21120 ( .A(n4903), .B(n4545), .Z(n2214) );
  AN2P U21121 ( .A(n4901), .B(n4546), .Z(n2243) );
  AN2P U21122 ( .A(n5221), .B(n4546), .Z(n2270) );
  AN2P U21123 ( .A(n5221), .B(n4900), .Z(n2284) );
  AN2P U21124 ( .A(n4899), .B(n4545), .Z(n2318) );
  AN2P U21125 ( .A(n4544), .B(n4898), .Z(n2331) );
  AN2P U21126 ( .A(n5223), .B(n4545), .Z(n2366) );
  AN2P U21127 ( .A(n5223), .B(n4897), .Z(n2373) );
  AN2P U21128 ( .A(n5223), .B(n4897), .Z(n2376) );
  AN2P U21129 ( .A(n5224), .B(n4898), .Z(n2402) );
  AN2P U21130 ( .A(n4899), .B(n4546), .Z(n2409) );
  AN2P U21131 ( .A(n4545), .B(n5224), .Z(n2430) );
  AN2P U21132 ( .A(n4899), .B(n5224), .Z(n2446) );
  AN2P U21133 ( .A(n5224), .B(n4545), .Z(n2453) );
  AN2P U21134 ( .A(n4545), .B(n5225), .Z(n2458) );
  AN2P U21135 ( .A(n5225), .B(n4898), .Z(n2468) );
  AN2P U21136 ( .A(n4547), .B(n5225), .Z(n2482) );
  AN2P U21137 ( .A(n4897), .B(n4546), .Z(n2488) );
  AN2P U21138 ( .A(n4897), .B(n4545), .Z(n2512) );
  AN2P U21139 ( .A(n5226), .B(n4900), .Z(n2537) );
  AN2P U21140 ( .A(n5226), .B(n4900), .Z(n2542) );
  AN2P U21141 ( .A(n5226), .B(n4545), .Z(n2546) );
  AN2P U21142 ( .A(n5226), .B(n4901), .Z(n2550) );
  AN2P U21143 ( .A(n5226), .B(n4902), .Z(n2565) );
  AN2P U21144 ( .A(n4902), .B(n4545), .Z(n2570) );
  AN2P U21145 ( .A(n4901), .B(n4546), .Z(n2613) );
  AN2P U21146 ( .A(n4902), .B(n4546), .Z(n2626) );
  AN2P U21147 ( .A(n5224), .B(n4902), .Z(n2631) );
  AN2P U21148 ( .A(n5226), .B(n4547), .Z(n2645) );
  AN2P U21149 ( .A(n5226), .B(n4547), .Z(n2650) );
  AN2P U21150 ( .A(n4903), .B(n4547), .Z(n2661) );
  AN2P U21151 ( .A(n4902), .B(n4547), .Z(n2674) );
  AN2P U21152 ( .A(n5225), .B(n4547), .Z(n2701) );
  AN2P U21153 ( .A(n4546), .B(n5224), .Z(n2717) );
  AN2P U21154 ( .A(n5224), .B(n4902), .Z(n2723) );
  AN2P U21155 ( .A(n4902), .B(n5224), .Z(n2731) );
  AN2P U21156 ( .A(n5223), .B(n4545), .Z(n2761) );
  AN2P U21157 ( .A(n5223), .B(n4545), .Z(n2765) );
  AN2P U21158 ( .A(n4903), .B(n4545), .Z(n2772) );
  AN2P U21159 ( .A(n4903), .B(n4545), .Z(n2778) );
  AN2P U21160 ( .A(n4900), .B(n4545), .Z(n2844) );
  AN2P U21161 ( .A(n5229), .B(n4899), .Z(n2856) );
  AN2P U21162 ( .A(n5229), .B(n4898), .Z(n2878) );
  AN2P U21163 ( .A(n4898), .B(n4546), .Z(n2890) );
  AN2P U21164 ( .A(n5229), .B(n4898), .Z(n2893) );
  AN2P U21165 ( .A(n5229), .B(n4898), .Z(n2899) );
  AN2P U21166 ( .A(n4546), .B(n5228), .Z(n2919) );
  AN2P U21167 ( .A(n4547), .B(n5228), .Z(n2928) );
  AN2P U21168 ( .A(n4547), .B(n5228), .Z(n2934) );
  AN2P U21169 ( .A(n4900), .B(n4545), .Z(n2951) );
  AN2P U21170 ( .A(n4898), .B(n4544), .Z(n2992) );
  AN2P U21171 ( .A(n5228), .B(n4545), .Z(n2998) );
  AN2P U21172 ( .A(n5228), .B(n4897), .Z(n3007) );
  AN2P U21173 ( .A(n4897), .B(n4547), .Z(n3065) );
  AN2P U21174 ( .A(n5221), .B(n4898), .Z(n3071) );
  AN2P U21175 ( .A(n5222), .B(n4547), .Z(n3085) );
  AN2P U21176 ( .A(n5223), .B(n4546), .Z(n3094) );
  AN2P U21177 ( .A(n5223), .B(n4899), .Z(n3111) );
  AN2P U21178 ( .A(n5224), .B(n4899), .Z(n3127) );
  AN2P U21179 ( .A(n4899), .B(n5225), .Z(n3141) );
  AN2P U21180 ( .A(n4545), .B(n4901), .Z(n3192) );
  AN2P U21181 ( .A(n5226), .B(n4901), .Z(n3197) );
  AN2P U21182 ( .A(n5226), .B(n4901), .Z(n3202) );
  AN2P U21183 ( .A(n4901), .B(n4545), .Z(n3209) );
  AN2P U21184 ( .A(n4902), .B(n5226), .Z(n3225) );
  AN2P U21185 ( .A(n4902), .B(n5226), .Z(n3232) );
  AN2P U21186 ( .A(n5226), .B(n4545), .Z(n3242) );
  AN2P U21187 ( .A(n4544), .B(n4903), .Z(n3257) );
  AN2P U21188 ( .A(n5225), .B(n4545), .Z(n3293) );
  AN2P U21189 ( .A(n5224), .B(n4545), .Z(n3306) );
  AN2P U21190 ( .A(n5223), .B(n4546), .Z(n3352) );
  AN2P U21191 ( .A(n5223), .B(n4546), .Z(n3362) );
  AN2P U21192 ( .A(n4546), .B(n4897), .Z(n3377) );
  AN2P U21193 ( .A(n5222), .B(n4546), .Z(n3404) );
  AN2P U21194 ( .A(n5222), .B(n4898), .Z(n3408) );
  AN2P U21195 ( .A(n5222), .B(n4546), .Z(n3421) );
  AN2P U21196 ( .A(n4899), .B(n5222), .Z(n3430) );
  AN2P U21197 ( .A(n5221), .B(n4899), .Z(n3434) );
  AN2P U21198 ( .A(n4546), .B(n4899), .Z(n3440) );
  AN2P U21199 ( .A(n4899), .B(n4546), .Z(n3445) );
  AN2P U21200 ( .A(n5221), .B(n4899), .Z(n3451) );
  AN2P U21201 ( .A(n5230), .B(n4544), .Z(n3504) );
  AN2P U21202 ( .A(n5229), .B(n4544), .Z(n3523) );
  AN2P U21203 ( .A(n5228), .B(n4902), .Z(n3554) );
  AN2P U21204 ( .A(n4903), .B(n5228), .Z(n3590) );
  AN2P U21205 ( .A(n4903), .B(n4546), .Z(n3600) );
  AN2P U21206 ( .A(n4902), .B(n4546), .Z(n3612) );
  AN2P U21207 ( .A(n4288), .B(n1579), .Z(n3658) );
  AN2P U21208 ( .A(n1158), .B(n4331), .Z(n3686) );
  AN2P U21209 ( .A(n4331), .B(n1137), .Z(n3693) );
  AN2P U21210 ( .A(n4208), .B(n829), .Z(n3754) );
  AN2P U21211 ( .A(n4252), .B(n1559), .Z(n3781) );
  AN2P U21212 ( .A(n1541), .B(n4290), .Z(n3785) );
  AN2P U21213 ( .A(n4331), .B(n4252), .Z(n3787) );
  AN2P U21214 ( .A(n880), .B(n4252), .Z(n3793) );
  AN2P U21215 ( .A(n1139), .B(n4252), .Z(n3803) );
  AN2P U21216 ( .A(n4330), .B(n1122), .Z(n3810) );
  AN2P U21217 ( .A(n4331), .B(n1517), .Z(n3900) );
  OR2 U21218 ( .A(n404), .B(n3951), .Z(n1500) );
  AN2P U21219 ( .A(n4332), .B(n1095), .Z(n4011) );
  AN2P U21220 ( .A(n4332), .B(n4288), .Z(n4015) );
  AN2P U21221 ( .A(n4288), .B(n836), .Z(n4016) );
  AN2P U21222 ( .A(n4332), .B(n4251), .Z(n4025) );
  AN2P U21223 ( .A(n1758), .B(n4289), .Z(n4028) );
  AN2P U21224 ( .A(n1760), .B(n4332), .Z(n4030) );
  AN2P U21225 ( .A(n4332), .B(n1759), .Z(n4031) );
  AN2P U21226 ( .A(n4289), .B(n4251), .Z(n4037) );
  AN2P U21227 ( .A(n1295), .B(n4289), .Z(n4039) );
  AN2P U21228 ( .A(n4289), .B(n1297), .Z(n4041) );
  AN2P U21229 ( .A(n4332), .B(n1296), .Z(n4043) );
  AN2P U21230 ( .A(n4289), .B(n4251), .Z(n4049) );
  AN2P U21231 ( .A(n1028), .B(n4289), .Z(n4051) );
  AN2P U21232 ( .A(n4289), .B(n1031), .Z(n4053) );
  AN2P U21233 ( .A(n4333), .B(n1029), .Z(n4055) );
  AN2P U21234 ( .A(n4289), .B(n4252), .Z(n4068) );
  AN2P U21235 ( .A(n1581), .B(n4289), .Z(n4070) );
  AN2P U21236 ( .A(n4289), .B(n1584), .Z(n4072) );
  AN2P U21237 ( .A(n4333), .B(n1582), .Z(n4074) );
  AN2P U21238 ( .A(n1274), .B(n4289), .Z(n4085) );
  AN2P U21239 ( .A(n1868), .B(n4333), .Z(n4107) );
  AN2P U21240 ( .A(n4334), .B(n1869), .Z(n4110) );
  AN2P U21241 ( .A(n4290), .B(n4252), .Z(n4140) );
  AN2P U21242 ( .A(n1251), .B(n4290), .Z(n4142) );
  AN2P U21243 ( .A(n4290), .B(n1254), .Z(n4144) );
  AN2P U21244 ( .A(n4333), .B(n1252), .Z(n4146) );
  AN2P U21245 ( .A(n1977), .B(n4289), .Z(n4157) );
  AN2P U21246 ( .A(n1226), .B(n4290), .Z(n4165) );
  AN2P U21247 ( .A(n1227), .B(n4333), .Z(n4167) );
  AN2P U21248 ( .A(n5071), .B(n4333), .Z(n4169) );
  AN2P U21249 ( .A(n1506), .B(n4333), .Z(n4178) );
  AN2P U21250 ( .A(n1507), .B(n4289), .Z(n4179) );
  AN2P U21251 ( .A(n4254), .B(n1505), .Z(n4180) );
  IVA U21252 ( .A(n4218), .Z(n4211) );
  IVA U21253 ( .A(n4218), .Z(n4212) );
  IVA U21254 ( .A(n4218), .Z(n4213) );
  IVA U21255 ( .A(n4222), .Z(n4214) );
  IVA U21256 ( .A(n4222), .Z(n4215) );
  IVA U21257 ( .A(LogIn2[46]), .Z(n4216) );
  IVA U21258 ( .A(LogIn2[46]), .Z(n4217) );
  IVA U21259 ( .A(n4215), .Z(n4218) );
  IVA U21260 ( .A(n4270), .Z(n4223) );
  IVA U21261 ( .A(n4270), .Z(n4224) );
  IVA U21262 ( .A(n4275), .Z(n4225) );
  IVA U21263 ( .A(n4250), .Z(n4226) );
  IVA U21264 ( .A(n4263), .Z(n4227) );
  IVA U21265 ( .A(n4275), .Z(n4228) );
  IVA U21266 ( .A(LogIn2[45]), .Z(n4229) );
  IVA U21267 ( .A(LogIn2[45]), .Z(n4230) );
  IVA U21268 ( .A(n4272), .Z(n4231) );
  IVA U21269 ( .A(n4271), .Z(n4232) );
  IVA U21270 ( .A(n4271), .Z(n4233) );
  IVA U21271 ( .A(n4271), .Z(n4234) );
  IVA U21272 ( .A(n4271), .Z(n4235) );
  IVA U21273 ( .A(n4271), .Z(n4236) );
  IVA U21274 ( .A(n4271), .Z(n4237) );
  IVA U21275 ( .A(n4272), .Z(n4238) );
  IVA U21276 ( .A(n4272), .Z(n4239) );
  IVA U21277 ( .A(n4272), .Z(n4240) );
  IVA U21278 ( .A(n4273), .Z(n4241) );
  IVA U21279 ( .A(n4273), .Z(n4242) );
  IVA U21280 ( .A(n4273), .Z(n4243) );
  IVA U21281 ( .A(n4274), .Z(n4244) );
  IVA U21282 ( .A(n4274), .Z(n4245) );
  IVA U21283 ( .A(n4274), .Z(n4246) );
  IVA U21284 ( .A(n4275), .Z(n4247) );
  IVA U21285 ( .A(n4275), .Z(n4248) );
  IVA U21286 ( .A(n4275), .Z(n4249) );
  IV U21287 ( .A(n4223), .Z(n4250) );
  IVA U21288 ( .A(n4269), .Z(n4270) );
  IVA U21289 ( .A(n4227), .Z(n4271) );
  IVA U21290 ( .A(n4227), .Z(n4272) );
  IVA U21291 ( .A(n4227), .Z(n4273) );
  IVA U21292 ( .A(n4231), .Z(n4274) );
  IVA U21293 ( .A(n4230), .Z(n4275) );
  IVA U21294 ( .A(n4340), .Z(n4309) );
  IVA U21295 ( .A(LogIn2[43]), .Z(n4310) );
  IVA U21296 ( .A(LogIn2[43]), .Z(n4311) );
  IVA U21297 ( .A(LogIn2[43]), .Z(n4312) );
  IVA U21298 ( .A(n4358), .Z(n4313) );
  IVA U21299 ( .A(n4330), .Z(n4314) );
  IVA U21300 ( .A(n4354), .Z(n4315) );
  IVA U21301 ( .A(n4354), .Z(n4316) );
  IVA U21302 ( .A(n4354), .Z(n4317) );
  IVA U21303 ( .A(n4355), .Z(n4318) );
  IVA U21304 ( .A(n4355), .Z(n4319) );
  IVA U21305 ( .A(n4355), .Z(n4320) );
  IVA U21306 ( .A(n4356), .Z(n4321) );
  IVA U21307 ( .A(n4356), .Z(n4322) );
  IVA U21308 ( .A(n4356), .Z(n4323) );
  IVA U21309 ( .A(n4357), .Z(n4324) );
  IVA U21310 ( .A(n4357), .Z(n4325) );
  IVA U21311 ( .A(n4357), .Z(n4326) );
  IVA U21312 ( .A(n4358), .Z(n4327) );
  IVA U21313 ( .A(n4358), .Z(n4328) );
  IVA U21314 ( .A(n4358), .Z(n4329) );
  IV U21315 ( .A(n4309), .Z(n4330) );
  IVA U21316 ( .A(n4309), .Z(n4354) );
  IVA U21317 ( .A(n4328), .Z(n4355) );
  IVA U21318 ( .A(n4327), .Z(n4356) );
  IVA U21319 ( .A(n4314), .Z(n4357) );
  IVA U21320 ( .A(n4309), .Z(n4358) );
  IVA U21321 ( .A(n4659), .Z(n4359) );
  IVA U21322 ( .A(n4659), .Z(n4360) );
  IVA U21323 ( .A(n4660), .Z(n4361) );
  IVA U21324 ( .A(n4660), .Z(n4362) );
  IVA U21325 ( .A(n4660), .Z(n4363) );
  IVA U21326 ( .A(n4661), .Z(n4364) );
  IVA U21327 ( .A(n4661), .Z(n4365) );
  IVA U21328 ( .A(n4661), .Z(n4366) );
  IVA U21329 ( .A(n4662), .Z(n4367) );
  IVA U21330 ( .A(n4662), .Z(n4368) );
  IVA U21331 ( .A(n4662), .Z(n4369) );
  IVA U21332 ( .A(n4663), .Z(n4370) );
  IVA U21333 ( .A(n4663), .Z(n4371) );
  IVA U21334 ( .A(n4663), .Z(n4372) );
  IVA U21335 ( .A(n4664), .Z(n4373) );
  IVA U21336 ( .A(n4664), .Z(n4374) );
  IVA U21337 ( .A(n4664), .Z(n4375) );
  IVA U21338 ( .A(n4665), .Z(n4376) );
  IVA U21339 ( .A(n4665), .Z(n4377) );
  IVA U21340 ( .A(n4665), .Z(n4378) );
  IVA U21341 ( .A(n4666), .Z(n4379) );
  IVA U21342 ( .A(n4666), .Z(n4380) );
  IVA U21343 ( .A(n4666), .Z(n4381) );
  IVA U21344 ( .A(n4667), .Z(n4382) );
  IVA U21345 ( .A(n4667), .Z(n4383) );
  IVA U21346 ( .A(n4667), .Z(n4384) );
  IVA U21347 ( .A(n4668), .Z(n4385) );
  IVA U21348 ( .A(n4668), .Z(n4386) );
  IVA U21349 ( .A(n4668), .Z(n4387) );
  IVA U21350 ( .A(n4669), .Z(n4388) );
  IVA U21351 ( .A(n4669), .Z(n4389) );
  IVA U21352 ( .A(n4669), .Z(n4390) );
  IVA U21353 ( .A(n4670), .Z(n4391) );
  IVA U21354 ( .A(n4670), .Z(n4392) );
  IVA U21355 ( .A(n4670), .Z(n4393) );
  IVA U21356 ( .A(n4671), .Z(n4394) );
  IVA U21357 ( .A(n4671), .Z(n4395) );
  IVA U21358 ( .A(n4671), .Z(n4396) );
  IVA U21359 ( .A(n4672), .Z(n4397) );
  IVA U21360 ( .A(n4672), .Z(n4398) );
  IVA U21361 ( .A(n4672), .Z(n4399) );
  IVA U21362 ( .A(n4673), .Z(n4400) );
  IVA U21363 ( .A(n4673), .Z(n4401) );
  IVA U21364 ( .A(n4673), .Z(n4402) );
  IVA U21365 ( .A(n4674), .Z(n4403) );
  IVA U21366 ( .A(n4674), .Z(n4404) );
  IVA U21367 ( .A(n4674), .Z(n4405) );
  IVA U21368 ( .A(n4675), .Z(n4406) );
  IVA U21369 ( .A(n4675), .Z(n4407) );
  IVA U21370 ( .A(n4675), .Z(n4408) );
  IVA U21371 ( .A(n4676), .Z(n4409) );
  IVA U21372 ( .A(n4676), .Z(n4410) );
  IVA U21373 ( .A(n4676), .Z(n4411) );
  IVA U21374 ( .A(n4677), .Z(n4412) );
  IVA U21375 ( .A(n4677), .Z(n4413) );
  IVA U21376 ( .A(n4677), .Z(n4414) );
  IVA U21377 ( .A(n4678), .Z(n4415) );
  IVA U21378 ( .A(n4678), .Z(n4416) );
  IVA U21379 ( .A(n4678), .Z(n4417) );
  IVA U21380 ( .A(n4679), .Z(n4418) );
  IVA U21381 ( .A(n4679), .Z(n4419) );
  IVA U21382 ( .A(n4679), .Z(n4420) );
  IVA U21383 ( .A(n4680), .Z(n4421) );
  IVA U21384 ( .A(n4680), .Z(n4422) );
  IVA U21385 ( .A(n4680), .Z(n4423) );
  IVA U21386 ( .A(n4681), .Z(n4424) );
  IVA U21387 ( .A(n4681), .Z(n4425) );
  IVA U21388 ( .A(n4681), .Z(n4426) );
  IVA U21389 ( .A(n4682), .Z(n4427) );
  IVA U21390 ( .A(n4682), .Z(n4428) );
  IVA U21391 ( .A(n4682), .Z(n4429) );
  IVA U21392 ( .A(n4683), .Z(n4430) );
  IVA U21393 ( .A(n4683), .Z(n4431) );
  IVA U21394 ( .A(n4683), .Z(n4432) );
  IVA U21395 ( .A(n4684), .Z(n4433) );
  IVA U21396 ( .A(n4684), .Z(n4434) );
  IVA U21397 ( .A(n4684), .Z(n4435) );
  IVA U21398 ( .A(n4685), .Z(n4436) );
  IVA U21399 ( .A(n4685), .Z(n4437) );
  IVA U21400 ( .A(n4685), .Z(n4438) );
  IVA U21401 ( .A(n4686), .Z(n4439) );
  IVA U21402 ( .A(n4686), .Z(n4440) );
  IVA U21403 ( .A(n4686), .Z(n4441) );
  IVA U21404 ( .A(n4687), .Z(n4442) );
  IVA U21405 ( .A(n4687), .Z(n4443) );
  IVA U21406 ( .A(n4687), .Z(n4444) );
  IVA U21407 ( .A(n4688), .Z(n4445) );
  IVA U21408 ( .A(n4688), .Z(n4446) );
  IVA U21409 ( .A(n4688), .Z(n4447) );
  IVA U21410 ( .A(n4689), .Z(n4448) );
  IVA U21411 ( .A(n4689), .Z(n4449) );
  IVA U21412 ( .A(n4689), .Z(n4450) );
  IVA U21413 ( .A(n4690), .Z(n4451) );
  IVA U21414 ( .A(n4690), .Z(n4452) );
  IVA U21415 ( .A(n4690), .Z(n4453) );
  IVA U21416 ( .A(n4691), .Z(n4454) );
  IVA U21417 ( .A(n4691), .Z(n4455) );
  IVA U21418 ( .A(n4691), .Z(n4456) );
  IVA U21419 ( .A(n4692), .Z(n4457) );
  IVA U21420 ( .A(n4692), .Z(n4458) );
  IVA U21421 ( .A(n4692), .Z(n4459) );
  IVA U21422 ( .A(n4693), .Z(n4460) );
  IVA U21423 ( .A(n4693), .Z(n4461) );
  IVA U21424 ( .A(n4693), .Z(n4462) );
  IVA U21425 ( .A(n4694), .Z(n4463) );
  IVA U21426 ( .A(n4694), .Z(n4464) );
  IVA U21427 ( .A(n4694), .Z(n4465) );
  IVA U21428 ( .A(n4695), .Z(n4466) );
  IVA U21429 ( .A(n4695), .Z(n4467) );
  IVA U21430 ( .A(n4695), .Z(n4468) );
  IVA U21431 ( .A(n4696), .Z(n4469) );
  IVA U21432 ( .A(n4696), .Z(n4470) );
  IVA U21433 ( .A(n4696), .Z(n4471) );
  IVA U21434 ( .A(n4697), .Z(n4472) );
  IVA U21435 ( .A(n4697), .Z(n4473) );
  IVA U21436 ( .A(n4697), .Z(n4474) );
  IVA U21437 ( .A(n4698), .Z(n4475) );
  IVA U21438 ( .A(n4698), .Z(n4476) );
  IVA U21439 ( .A(n4698), .Z(n4477) );
  IVA U21440 ( .A(n4699), .Z(n4478) );
  IVA U21441 ( .A(n4699), .Z(n4479) );
  IVA U21442 ( .A(n4699), .Z(n4480) );
  IVA U21443 ( .A(n4700), .Z(n4481) );
  IVA U21444 ( .A(n4700), .Z(n4482) );
  IVA U21445 ( .A(n4700), .Z(n4483) );
  IVA U21446 ( .A(n4701), .Z(n4484) );
  IVA U21447 ( .A(n4701), .Z(n4485) );
  IVA U21448 ( .A(n4701), .Z(n4486) );
  IVA U21449 ( .A(n4702), .Z(n4487) );
  IVA U21450 ( .A(n4702), .Z(n4488) );
  IVA U21451 ( .A(n4702), .Z(n4489) );
  IVA U21452 ( .A(n4703), .Z(n4490) );
  IVA U21453 ( .A(n4703), .Z(n4491) );
  IVA U21454 ( .A(n4703), .Z(n4492) );
  IVA U21455 ( .A(n4704), .Z(n4493) );
  IVA U21456 ( .A(n4704), .Z(n4494) );
  IVA U21457 ( .A(n4704), .Z(n4495) );
  IVA U21458 ( .A(n4705), .Z(n4496) );
  IVA U21459 ( .A(n4705), .Z(n4497) );
  IVA U21460 ( .A(n4705), .Z(n4498) );
  IVA U21461 ( .A(n4706), .Z(n4499) );
  IVA U21462 ( .A(n4706), .Z(n4500) );
  IVA U21463 ( .A(n4706), .Z(n4501) );
  IVA U21464 ( .A(n4707), .Z(n4502) );
  IVA U21465 ( .A(n4707), .Z(n4503) );
  IVA U21466 ( .A(n4707), .Z(n4504) );
  IVA U21467 ( .A(n4708), .Z(n4505) );
  IVA U21468 ( .A(n4708), .Z(n4506) );
  IVA U21469 ( .A(n4708), .Z(n4507) );
  IVA U21470 ( .A(n4709), .Z(n4508) );
  IVA U21471 ( .A(n4709), .Z(n4509) );
  IVA U21472 ( .A(n4709), .Z(n4510) );
  IVA U21473 ( .A(n4710), .Z(n4511) );
  IVA U21474 ( .A(n4710), .Z(n4512) );
  IVA U21475 ( .A(n4710), .Z(n4513) );
  IVA U21476 ( .A(n4711), .Z(n4514) );
  IVA U21477 ( .A(n4711), .Z(n4515) );
  IVA U21478 ( .A(n4711), .Z(n4516) );
  IVA U21479 ( .A(n4712), .Z(n4517) );
  IVA U21480 ( .A(n4712), .Z(n4518) );
  IVA U21481 ( .A(n4712), .Z(n4519) );
  IVA U21482 ( .A(n4713), .Z(n4520) );
  IVA U21483 ( .A(n4713), .Z(n4521) );
  IVA U21484 ( .A(n4713), .Z(n4522) );
  IVA U21485 ( .A(n4714), .Z(n4523) );
  IVA U21486 ( .A(n4714), .Z(n4524) );
  IVA U21487 ( .A(n4714), .Z(n4525) );
  IVA U21488 ( .A(n4715), .Z(n4526) );
  IVA U21489 ( .A(n4715), .Z(n4527) );
  IVA U21490 ( .A(n4715), .Z(n4528) );
  IVA U21491 ( .A(n4716), .Z(n4529) );
  IVA U21492 ( .A(n4716), .Z(n4530) );
  IVA U21493 ( .A(n4716), .Z(n4531) );
  IVA U21494 ( .A(n4717), .Z(n4532) );
  IVA U21495 ( .A(n4717), .Z(n4533) );
  IVA U21496 ( .A(n4717), .Z(n4534) );
  IVA U21497 ( .A(n4718), .Z(n4535) );
  IVA U21498 ( .A(n4718), .Z(n4536) );
  IVA U21499 ( .A(n4718), .Z(n4537) );
  IVA U21500 ( .A(n4719), .Z(n4538) );
  IVA U21501 ( .A(n4719), .Z(n4539) );
  IVA U21502 ( .A(n4719), .Z(n4540) );
  IVA U21503 ( .A(n4720), .Z(n4541) );
  IVA U21504 ( .A(n4720), .Z(n4542) );
  IVA U21505 ( .A(n4720), .Z(n4543) );
  IV U21506 ( .A(n4367), .Z(n4544) );
  IVA U21507 ( .A(n4666), .Z(n4638) );
  IVA U21508 ( .A(n4667), .Z(n4639) );
  IVA U21509 ( .A(n4665), .Z(n4640) );
  IVA U21510 ( .A(n4696), .Z(n4641) );
  IVA U21511 ( .A(LogIn2[42]), .Z(n4642) );
  IVA U21512 ( .A(LogIn2[42]), .Z(n4643) );
  IVA U21513 ( .A(LogIn2[42]), .Z(n4644) );
  IVA U21514 ( .A(LogIn2[42]), .Z(n4645) );
  IVA U21515 ( .A(LogIn2[42]), .Z(n4646) );
  IVA U21516 ( .A(LogIn2[42]), .Z(n4647) );
  IVA U21517 ( .A(n4709), .Z(n4648) );
  IVA U21518 ( .A(n4719), .Z(n4649) );
  IVA U21519 ( .A(n4667), .Z(n4650) );
  IVA U21520 ( .A(n4673), .Z(n4651) );
  IVA U21521 ( .A(n4701), .Z(n4652) );
  IVA U21522 ( .A(LogIn2[42]), .Z(n4653) );
  IVA U21523 ( .A(n4666), .Z(n4654) );
  IVA U21524 ( .A(LogIn2[42]), .Z(n4655) );
  IVA U21525 ( .A(n4694), .Z(n4656) );
  IVA U21526 ( .A(LogIn2[42]), .Z(n4657) );
  IVA U21527 ( .A(LogIn2[42]), .Z(n4658) );
  IVA U21528 ( .A(n4658), .Z(n4659) );
  IVA U21529 ( .A(n4658), .Z(n4660) );
  IVA U21530 ( .A(n4658), .Z(n4661) );
  IVA U21531 ( .A(n4657), .Z(n4662) );
  IVA U21532 ( .A(n4657), .Z(n4663) );
  IVA U21533 ( .A(n4657), .Z(n4664) );
  IVA U21534 ( .A(n4656), .Z(n4665) );
  IVA U21535 ( .A(n4656), .Z(n4666) );
  IVA U21536 ( .A(n4656), .Z(n4667) );
  IVA U21537 ( .A(n4655), .Z(n4668) );
  IVA U21538 ( .A(n4655), .Z(n4669) );
  IVA U21539 ( .A(n4655), .Z(n4670) );
  IVA U21540 ( .A(n4654), .Z(n4671) );
  IVA U21541 ( .A(n4654), .Z(n4672) );
  IVA U21542 ( .A(n4654), .Z(n4673) );
  IVA U21543 ( .A(n4653), .Z(n4674) );
  IVA U21544 ( .A(n4653), .Z(n4675) );
  IVA U21545 ( .A(n4653), .Z(n4676) );
  IVA U21546 ( .A(n4652), .Z(n4677) );
  IVA U21547 ( .A(n4652), .Z(n4678) );
  IVA U21548 ( .A(n4652), .Z(n4679) );
  IVA U21549 ( .A(n4651), .Z(n4680) );
  IVA U21550 ( .A(n4651), .Z(n4681) );
  IVA U21551 ( .A(n4651), .Z(n4682) );
  IVA U21552 ( .A(n4650), .Z(n4683) );
  IVA U21553 ( .A(n4650), .Z(n4684) );
  IVA U21554 ( .A(n4650), .Z(n4685) );
  IVA U21555 ( .A(n4649), .Z(n4686) );
  IVA U21556 ( .A(n4649), .Z(n4687) );
  IVA U21557 ( .A(n4649), .Z(n4688) );
  IVA U21558 ( .A(n4648), .Z(n4689) );
  IVA U21559 ( .A(n4648), .Z(n4690) );
  IVA U21560 ( .A(n4648), .Z(n4691) );
  IVA U21561 ( .A(n4647), .Z(n4692) );
  IVA U21562 ( .A(n4647), .Z(n4693) );
  IVA U21563 ( .A(n4647), .Z(n4694) );
  IVA U21564 ( .A(n4646), .Z(n4695) );
  IVA U21565 ( .A(n4646), .Z(n4696) );
  IVA U21566 ( .A(n4646), .Z(n4697) );
  IVA U21567 ( .A(n4645), .Z(n4698) );
  IVA U21568 ( .A(n4645), .Z(n4699) );
  IVA U21569 ( .A(n4645), .Z(n4700) );
  IVA U21570 ( .A(n4644), .Z(n4701) );
  IVA U21571 ( .A(n4644), .Z(n4702) );
  IVA U21572 ( .A(n4644), .Z(n4703) );
  IVA U21573 ( .A(n4643), .Z(n4704) );
  IVA U21574 ( .A(n4643), .Z(n4705) );
  IVA U21575 ( .A(n4643), .Z(n4706) );
  IVA U21576 ( .A(n4642), .Z(n4707) );
  IVA U21577 ( .A(n4642), .Z(n4708) );
  IVA U21578 ( .A(n4642), .Z(n4709) );
  IVA U21579 ( .A(n4641), .Z(n4710) );
  IVA U21580 ( .A(n4641), .Z(n4711) );
  IVA U21581 ( .A(n4641), .Z(n4712) );
  IVA U21582 ( .A(n4640), .Z(n4713) );
  IVA U21583 ( .A(n4640), .Z(n4714) );
  IVA U21584 ( .A(n4640), .Z(n4715) );
  IVA U21585 ( .A(n4639), .Z(n4716) );
  IVA U21586 ( .A(n4639), .Z(n4717) );
  IVA U21587 ( .A(n4639), .Z(n4718) );
  IVA U21588 ( .A(n4638), .Z(n4719) );
  IVA U21589 ( .A(n4638), .Z(n4720) );
  IVA U21590 ( .A(n4999), .Z(n4721) );
  IVA U21591 ( .A(n4999), .Z(n4722) );
  IVA U21592 ( .A(n5000), .Z(n4723) );
  IVA U21593 ( .A(n5000), .Z(n4724) );
  IVA U21594 ( .A(n5000), .Z(n4725) );
  IVA U21595 ( .A(n5001), .Z(n4726) );
  IVA U21596 ( .A(n5001), .Z(n4727) );
  IVA U21597 ( .A(n5001), .Z(n4728) );
  IVA U21598 ( .A(n5002), .Z(n4729) );
  IVA U21599 ( .A(n5002), .Z(n4730) );
  IVA U21600 ( .A(n5002), .Z(n4731) );
  IVA U21601 ( .A(n5003), .Z(n4732) );
  IVA U21602 ( .A(n5003), .Z(n4733) );
  IVA U21603 ( .A(n5003), .Z(n4734) );
  IVA U21604 ( .A(n5004), .Z(n4735) );
  IVA U21605 ( .A(n5004), .Z(n4736) );
  IVA U21606 ( .A(n5004), .Z(n4737) );
  IVA U21607 ( .A(n5005), .Z(n4738) );
  IVA U21608 ( .A(n5005), .Z(n4739) );
  IVA U21609 ( .A(n5005), .Z(n4740) );
  IVA U21610 ( .A(n5006), .Z(n4741) );
  IVA U21611 ( .A(n5006), .Z(n4742) );
  IVA U21612 ( .A(n5006), .Z(n4743) );
  IVA U21613 ( .A(n5007), .Z(n4744) );
  IVA U21614 ( .A(n5007), .Z(n4745) );
  IVA U21615 ( .A(n5007), .Z(n4746) );
  IVA U21616 ( .A(n5008), .Z(n4747) );
  IVA U21617 ( .A(n5008), .Z(n4748) );
  IVA U21618 ( .A(n5008), .Z(n4749) );
  IVA U21619 ( .A(n5009), .Z(n4750) );
  IVA U21620 ( .A(n5009), .Z(n4751) );
  IVA U21621 ( .A(n5009), .Z(n4752) );
  IVA U21622 ( .A(n5010), .Z(n4753) );
  IVA U21623 ( .A(n5010), .Z(n4754) );
  IVA U21624 ( .A(n5010), .Z(n4755) );
  IVA U21625 ( .A(n5011), .Z(n4756) );
  IVA U21626 ( .A(n5011), .Z(n4757) );
  IVA U21627 ( .A(n5011), .Z(n4758) );
  IVA U21628 ( .A(n5012), .Z(n4759) );
  IVA U21629 ( .A(n5012), .Z(n4760) );
  IVA U21630 ( .A(n5012), .Z(n4761) );
  IVA U21631 ( .A(n5013), .Z(n4762) );
  IVA U21632 ( .A(n5013), .Z(n4763) );
  IVA U21633 ( .A(n5013), .Z(n4764) );
  IVA U21634 ( .A(n5014), .Z(n4765) );
  IVA U21635 ( .A(n5014), .Z(n4766) );
  IVA U21636 ( .A(n5014), .Z(n4767) );
  IVA U21637 ( .A(n5015), .Z(n4768) );
  IVA U21638 ( .A(n5015), .Z(n4769) );
  IVA U21639 ( .A(n5015), .Z(n4770) );
  IVA U21640 ( .A(n5016), .Z(n4771) );
  IVA U21641 ( .A(n5016), .Z(n4772) );
  IVA U21642 ( .A(n5016), .Z(n4773) );
  IVA U21643 ( .A(n5017), .Z(n4774) );
  IVA U21644 ( .A(n5017), .Z(n4775) );
  IVA U21645 ( .A(n5017), .Z(n4776) );
  IVA U21646 ( .A(n5018), .Z(n4777) );
  IVA U21647 ( .A(n5018), .Z(n4778) );
  IVA U21648 ( .A(n5018), .Z(n4779) );
  IVA U21649 ( .A(n5019), .Z(n4780) );
  IVA U21650 ( .A(n5019), .Z(n4781) );
  IVA U21651 ( .A(n5019), .Z(n4782) );
  IVA U21652 ( .A(n5020), .Z(n4783) );
  IVA U21653 ( .A(n5020), .Z(n4784) );
  IVA U21654 ( .A(n5020), .Z(n4785) );
  IVA U21655 ( .A(n5021), .Z(n4786) );
  IVA U21656 ( .A(n5021), .Z(n4787) );
  IVA U21657 ( .A(n5021), .Z(n4788) );
  IVA U21658 ( .A(n5022), .Z(n4789) );
  IVA U21659 ( .A(n5022), .Z(n4790) );
  IVA U21660 ( .A(n5022), .Z(n4791) );
  IVA U21661 ( .A(n5023), .Z(n4792) );
  IVA U21662 ( .A(n5023), .Z(n4793) );
  IVA U21663 ( .A(n5023), .Z(n4794) );
  IVA U21664 ( .A(n5024), .Z(n4795) );
  IVA U21665 ( .A(n5024), .Z(n4796) );
  IVA U21666 ( .A(n5024), .Z(n4797) );
  IVA U21667 ( .A(n5025), .Z(n4798) );
  IVA U21668 ( .A(n5025), .Z(n4799) );
  IVA U21669 ( .A(n5025), .Z(n4800) );
  IVA U21670 ( .A(n5026), .Z(n4801) );
  IVA U21671 ( .A(n5026), .Z(n4802) );
  IVA U21672 ( .A(n5026), .Z(n4803) );
  IVA U21673 ( .A(n5027), .Z(n4804) );
  IVA U21674 ( .A(n5027), .Z(n4805) );
  IVA U21675 ( .A(n5027), .Z(n4806) );
  IVA U21676 ( .A(n5028), .Z(n4807) );
  IVA U21677 ( .A(n5028), .Z(n4808) );
  IVA U21678 ( .A(n5028), .Z(n4809) );
  IVA U21679 ( .A(n5029), .Z(n4810) );
  IVA U21680 ( .A(n5029), .Z(n4811) );
  IVA U21681 ( .A(n5029), .Z(n4812) );
  IVA U21682 ( .A(n5030), .Z(n4813) );
  IVA U21683 ( .A(n5030), .Z(n4814) );
  IVA U21684 ( .A(n5030), .Z(n4815) );
  IVA U21685 ( .A(n5031), .Z(n4816) );
  IVA U21686 ( .A(n5031), .Z(n4817) );
  IVA U21687 ( .A(n5031), .Z(n4818) );
  IVA U21688 ( .A(n5032), .Z(n4819) );
  IVA U21689 ( .A(n5032), .Z(n4820) );
  IVA U21690 ( .A(n5032), .Z(n4821) );
  IVA U21691 ( .A(n5033), .Z(n4822) );
  IVA U21692 ( .A(n5033), .Z(n4823) );
  IVA U21693 ( .A(n5033), .Z(n4824) );
  IVA U21694 ( .A(n5034), .Z(n4825) );
  IVA U21695 ( .A(n5034), .Z(n4826) );
  IVA U21696 ( .A(n5034), .Z(n4827) );
  IVA U21697 ( .A(n5035), .Z(n4828) );
  IVA U21698 ( .A(n5035), .Z(n4829) );
  IVA U21699 ( .A(n5035), .Z(n4830) );
  IVA U21700 ( .A(n5036), .Z(n4831) );
  IVA U21701 ( .A(n5036), .Z(n4832) );
  IVA U21702 ( .A(n5036), .Z(n4833) );
  IVA U21703 ( .A(n5037), .Z(n4834) );
  IVA U21704 ( .A(n5037), .Z(n4835) );
  IVA U21705 ( .A(n5037), .Z(n4836) );
  IVA U21706 ( .A(n5038), .Z(n4837) );
  IVA U21707 ( .A(n5038), .Z(n4838) );
  IVA U21708 ( .A(n5038), .Z(n4839) );
  IVA U21709 ( .A(n5039), .Z(n4840) );
  IVA U21710 ( .A(n5039), .Z(n4841) );
  IVA U21711 ( .A(n5039), .Z(n4842) );
  IVA U21712 ( .A(n5040), .Z(n4843) );
  IVA U21713 ( .A(n5040), .Z(n4844) );
  IVA U21714 ( .A(n5040), .Z(n4845) );
  IVA U21715 ( .A(n5041), .Z(n4846) );
  IVA U21716 ( .A(n5041), .Z(n4847) );
  IVA U21717 ( .A(n5041), .Z(n4848) );
  IVA U21718 ( .A(n5042), .Z(n4849) );
  IVA U21719 ( .A(n5042), .Z(n4850) );
  IVA U21720 ( .A(n5042), .Z(n4851) );
  IVA U21721 ( .A(n5043), .Z(n4852) );
  IVA U21722 ( .A(n5043), .Z(n4853) );
  IVA U21723 ( .A(n5043), .Z(n4854) );
  IVA U21724 ( .A(n5044), .Z(n4855) );
  IVA U21725 ( .A(n5044), .Z(n4856) );
  IVA U21726 ( .A(n5044), .Z(n4857) );
  IVA U21727 ( .A(n5045), .Z(n4858) );
  IVA U21728 ( .A(n5045), .Z(n4859) );
  IVA U21729 ( .A(n5045), .Z(n4860) );
  IVA U21730 ( .A(n5046), .Z(n4861) );
  IVA U21731 ( .A(n5046), .Z(n4862) );
  IVA U21732 ( .A(n5046), .Z(n4863) );
  IVA U21733 ( .A(n5047), .Z(n4864) );
  IVA U21734 ( .A(n5047), .Z(n4865) );
  IVA U21735 ( .A(n5047), .Z(n4866) );
  IVA U21736 ( .A(n5048), .Z(n4867) );
  IVA U21737 ( .A(n5048), .Z(n4868) );
  IVA U21738 ( .A(n5048), .Z(n4869) );
  IVA U21739 ( .A(n5049), .Z(n4870) );
  IVA U21740 ( .A(n5049), .Z(n4871) );
  IVA U21741 ( .A(n5049), .Z(n4872) );
  IVA U21742 ( .A(n5050), .Z(n4873) );
  IVA U21743 ( .A(n5050), .Z(n4874) );
  IVA U21744 ( .A(n5050), .Z(n4875) );
  IVA U21745 ( .A(n5051), .Z(n4876) );
  IVA U21746 ( .A(n5051), .Z(n4877) );
  IVA U21747 ( .A(n5051), .Z(n4878) );
  IVA U21748 ( .A(n5052), .Z(n4879) );
  IVA U21749 ( .A(n5052), .Z(n4880) );
  IVA U21750 ( .A(n5052), .Z(n4881) );
  IVA U21751 ( .A(n5053), .Z(n4882) );
  IVA U21752 ( .A(n5053), .Z(n4883) );
  IVA U21753 ( .A(n5053), .Z(n4884) );
  IVA U21754 ( .A(n5054), .Z(n4885) );
  IVA U21755 ( .A(n5054), .Z(n4886) );
  IVA U21756 ( .A(n5054), .Z(n4887) );
  IVA U21757 ( .A(n5055), .Z(n4888) );
  IVA U21758 ( .A(n5055), .Z(n4889) );
  IVA U21759 ( .A(n5055), .Z(n4890) );
  IVA U21760 ( .A(n5056), .Z(n4891) );
  IVA U21761 ( .A(n5056), .Z(n4892) );
  IVA U21762 ( .A(n5056), .Z(n4893) );
  IVA U21763 ( .A(n5057), .Z(n4894) );
  IVA U21764 ( .A(n5057), .Z(n4895) );
  IVA U21765 ( .A(n5057), .Z(n4896) );
  IVA U21766 ( .A(n5043), .Z(n4979) );
  IVA U21767 ( .A(LogIn2[41]), .Z(n4980) );
  IVA U21768 ( .A(n5006), .Z(n4981) );
  IVA U21769 ( .A(n5004), .Z(n4982) );
  IVA U21770 ( .A(LogIn2[41]), .Z(n4983) );
  IVA U21771 ( .A(LogIn2[41]), .Z(n4984) );
  IVA U21772 ( .A(n5004), .Z(n4985) );
  IVA U21773 ( .A(n5004), .Z(n4986) );
  IVA U21774 ( .A(n5045), .Z(n4987) );
  IVA U21775 ( .A(n4999), .Z(n4988) );
  IVA U21776 ( .A(LogIn2[41]), .Z(n4989) );
  IVA U21777 ( .A(n5049), .Z(n4990) );
  IVA U21778 ( .A(LogIn2[41]), .Z(n4991) );
  IVA U21779 ( .A(LogIn2[41]), .Z(n4992) );
  IVA U21780 ( .A(n5012), .Z(n4993) );
  IVA U21781 ( .A(LogIn2[41]), .Z(n4994) );
  IVA U21782 ( .A(n5057), .Z(n4995) );
  IVA U21783 ( .A(LogIn2[41]), .Z(n4996) );
  IVA U21784 ( .A(LogIn2[41]), .Z(n4997) );
  IVA U21785 ( .A(LogIn2[41]), .Z(n4998) );
  IVA U21786 ( .A(n4998), .Z(n4999) );
  IVA U21787 ( .A(n4998), .Z(n5000) );
  IVA U21788 ( .A(n4998), .Z(n5001) );
  IVA U21789 ( .A(n4997), .Z(n5002) );
  IVA U21790 ( .A(n4997), .Z(n5003) );
  IVA U21791 ( .A(n4997), .Z(n5004) );
  IVA U21792 ( .A(n4996), .Z(n5005) );
  IVA U21793 ( .A(n4996), .Z(n5006) );
  IVA U21794 ( .A(n4996), .Z(n5007) );
  IVA U21795 ( .A(n4995), .Z(n5008) );
  IVA U21796 ( .A(n4995), .Z(n5009) );
  IVA U21797 ( .A(n4995), .Z(n5010) );
  IVA U21798 ( .A(n4994), .Z(n5011) );
  IVA U21799 ( .A(n4994), .Z(n5012) );
  IVA U21800 ( .A(n4994), .Z(n5013) );
  IVA U21801 ( .A(n4993), .Z(n5014) );
  IVA U21802 ( .A(n4993), .Z(n5015) );
  IVA U21803 ( .A(n4993), .Z(n5016) );
  IVA U21804 ( .A(n4992), .Z(n5017) );
  IVA U21805 ( .A(n4992), .Z(n5018) );
  IVA U21806 ( .A(n4992), .Z(n5019) );
  IVA U21807 ( .A(n4991), .Z(n5020) );
  IVA U21808 ( .A(n4991), .Z(n5021) );
  IVA U21809 ( .A(n4991), .Z(n5022) );
  IVA U21810 ( .A(n4990), .Z(n5023) );
  IVA U21811 ( .A(n4990), .Z(n5024) );
  IVA U21812 ( .A(n4990), .Z(n5025) );
  IVA U21813 ( .A(n4989), .Z(n5026) );
  IVA U21814 ( .A(n4989), .Z(n5027) );
  IVA U21815 ( .A(n4989), .Z(n5028) );
  IVA U21816 ( .A(n4988), .Z(n5029) );
  IVA U21817 ( .A(n4988), .Z(n5030) );
  IVA U21818 ( .A(n4988), .Z(n5031) );
  IVA U21819 ( .A(n4987), .Z(n5032) );
  IVA U21820 ( .A(n4987), .Z(n5033) );
  IVA U21821 ( .A(n4987), .Z(n5034) );
  IVA U21822 ( .A(n4986), .Z(n5035) );
  IVA U21823 ( .A(n4986), .Z(n5036) );
  IVA U21824 ( .A(n4986), .Z(n5037) );
  IVA U21825 ( .A(n4985), .Z(n5038) );
  IVA U21826 ( .A(n4985), .Z(n5039) );
  IVA U21827 ( .A(n4985), .Z(n5040) );
  IVA U21828 ( .A(n4984), .Z(n5041) );
  IVA U21829 ( .A(n4984), .Z(n5042) );
  IVA U21830 ( .A(n4984), .Z(n5043) );
  IVA U21831 ( .A(n4983), .Z(n5044) );
  IVA U21832 ( .A(n4983), .Z(n5045) );
  IVA U21833 ( .A(n4983), .Z(n5046) );
  IVA U21834 ( .A(n4982), .Z(n5047) );
  IVA U21835 ( .A(n4982), .Z(n5048) );
  IVA U21836 ( .A(n4982), .Z(n5049) );
  IVA U21837 ( .A(n4981), .Z(n5050) );
  IVA U21838 ( .A(n4981), .Z(n5051) );
  IVA U21839 ( .A(n4981), .Z(n5052) );
  IVA U21840 ( .A(n4980), .Z(n5053) );
  IVA U21841 ( .A(n4980), .Z(n5054) );
  IVA U21842 ( .A(n4980), .Z(n5055) );
  IVA U21843 ( .A(n4979), .Z(n5056) );
  IVA U21844 ( .A(n4979), .Z(n5057) );
  IVA U21845 ( .A(n5307), .Z(n5058) );
  IVA U21846 ( .A(n5308), .Z(n5059) );
  IVA U21847 ( .A(n5308), .Z(n5060) );
  IVA U21848 ( .A(n5308), .Z(n5061) );
  IVA U21849 ( .A(n5309), .Z(n5062) );
  IVA U21850 ( .A(n5309), .Z(n5063) );
  IVA U21851 ( .A(n5309), .Z(n5064) );
  IVA U21852 ( .A(n5310), .Z(n5065) );
  IVA U21853 ( .A(n5310), .Z(n5066) );
  IVA U21854 ( .A(n5310), .Z(n5067) );
  IVA U21855 ( .A(n5311), .Z(n5068) );
  IVA U21856 ( .A(n5311), .Z(n5069) );
  IVA U21857 ( .A(n5311), .Z(n5070) );
  IVA U21858 ( .A(n5312), .Z(n5071) );
  IVA U21859 ( .A(n5312), .Z(n5072) );
  IVA U21860 ( .A(n5312), .Z(n5073) );
  IVA U21861 ( .A(n5313), .Z(n5074) );
  IVA U21862 ( .A(n5313), .Z(n5075) );
  IVA U21863 ( .A(n5313), .Z(n5076) );
  IVA U21864 ( .A(n5314), .Z(n5077) );
  IVA U21865 ( .A(n5314), .Z(n5078) );
  IVA U21866 ( .A(n5314), .Z(n5079) );
  IVA U21867 ( .A(n5315), .Z(n5080) );
  IVA U21868 ( .A(n5315), .Z(n5081) );
  IVA U21869 ( .A(n5315), .Z(n5082) );
  IVA U21870 ( .A(n5316), .Z(n5083) );
  IVA U21871 ( .A(n5316), .Z(n5084) );
  IVA U21872 ( .A(n5316), .Z(n5085) );
  IVA U21873 ( .A(n5317), .Z(n5086) );
  IVA U21874 ( .A(n5317), .Z(n5087) );
  IVA U21875 ( .A(n5317), .Z(n5088) );
  IVA U21876 ( .A(n5318), .Z(n5089) );
  IVA U21877 ( .A(n5318), .Z(n5090) );
  IVA U21878 ( .A(n5318), .Z(n5091) );
  IVA U21879 ( .A(n5319), .Z(n5092) );
  IVA U21880 ( .A(n5319), .Z(n5093) );
  IVA U21881 ( .A(n5319), .Z(n5094) );
  IVA U21882 ( .A(n5320), .Z(n5095) );
  IVA U21883 ( .A(n5320), .Z(n5096) );
  IVA U21884 ( .A(n5320), .Z(n5097) );
  IVA U21885 ( .A(n5321), .Z(n5098) );
  IVA U21886 ( .A(n5321), .Z(n5099) );
  IVA U21887 ( .A(n5321), .Z(n5100) );
  IVA U21888 ( .A(n5322), .Z(n5101) );
  IVA U21889 ( .A(n5322), .Z(n5102) );
  IVA U21890 ( .A(n5322), .Z(n5103) );
  IVA U21891 ( .A(n5323), .Z(n5104) );
  IVA U21892 ( .A(n5323), .Z(n5105) );
  IVA U21893 ( .A(n5323), .Z(n5106) );
  IVA U21894 ( .A(n5324), .Z(n5107) );
  IVA U21895 ( .A(n5324), .Z(n5108) );
  IVA U21896 ( .A(n5324), .Z(n5109) );
  IVA U21897 ( .A(n5325), .Z(n5110) );
  IVA U21898 ( .A(n5325), .Z(n5111) );
  IVA U21899 ( .A(n5325), .Z(n5112) );
  IVA U21900 ( .A(n5326), .Z(n5113) );
  IVA U21901 ( .A(n5326), .Z(n5114) );
  IVA U21902 ( .A(n5326), .Z(n5115) );
  IVA U21903 ( .A(n5327), .Z(n5116) );
  IVA U21904 ( .A(n5327), .Z(n5117) );
  IVA U21905 ( .A(n5327), .Z(n5118) );
  IVA U21906 ( .A(n5328), .Z(n5119) );
  IVA U21907 ( .A(n5328), .Z(n5120) );
  IVA U21908 ( .A(n5328), .Z(n5121) );
  IVA U21909 ( .A(n5329), .Z(n5122) );
  IVA U21910 ( .A(n5329), .Z(n5123) );
  IVA U21911 ( .A(n5329), .Z(n5124) );
  IVA U21912 ( .A(n5330), .Z(n5125) );
  IVA U21913 ( .A(n5330), .Z(n5126) );
  IVA U21914 ( .A(n5330), .Z(n5127) );
  IVA U21915 ( .A(n5331), .Z(n5128) );
  IVA U21916 ( .A(n5331), .Z(n5129) );
  IVA U21917 ( .A(n5331), .Z(n5130) );
  IVA U21918 ( .A(n5332), .Z(n5131) );
  IVA U21919 ( .A(n5332), .Z(n5132) );
  IVA U21920 ( .A(n5332), .Z(n5133) );
  IVA U21921 ( .A(n5333), .Z(n5134) );
  IVA U21922 ( .A(n5333), .Z(n5135) );
  IVA U21923 ( .A(n5333), .Z(n5136) );
  IVA U21924 ( .A(n5334), .Z(n5137) );
  IVA U21925 ( .A(n5334), .Z(n5138) );
  IVA U21926 ( .A(n5334), .Z(n5139) );
  IVA U21927 ( .A(n5335), .Z(n5140) );
  IVA U21928 ( .A(n5335), .Z(n5141) );
  IVA U21929 ( .A(n5335), .Z(n5142) );
  IVA U21930 ( .A(n5336), .Z(n5143) );
  IVA U21931 ( .A(n5336), .Z(n5144) );
  IVA U21932 ( .A(n5336), .Z(n5145) );
  IVA U21933 ( .A(n5337), .Z(n5146) );
  IVA U21934 ( .A(n5337), .Z(n5147) );
  IVA U21935 ( .A(n5337), .Z(n5148) );
  IVA U21936 ( .A(n5338), .Z(n5149) );
  IVA U21937 ( .A(n5338), .Z(n5150) );
  IVA U21938 ( .A(n5338), .Z(n5151) );
  IVA U21939 ( .A(n5339), .Z(n5152) );
  IVA U21940 ( .A(n5339), .Z(n5153) );
  IVA U21941 ( .A(n5339), .Z(n5154) );
  IVA U21942 ( .A(n5340), .Z(n5155) );
  IVA U21943 ( .A(n5340), .Z(n5156) );
  IVA U21944 ( .A(n5340), .Z(n5157) );
  IVA U21945 ( .A(n5341), .Z(n5158) );
  IVA U21946 ( .A(n5341), .Z(n5159) );
  IVA U21947 ( .A(n5341), .Z(n5160) );
  IVA U21948 ( .A(n5342), .Z(n5161) );
  IVA U21949 ( .A(n5342), .Z(n5162) );
  IVA U21950 ( .A(n5342), .Z(n5163) );
  IVA U21951 ( .A(n5343), .Z(n5164) );
  IVA U21952 ( .A(n5343), .Z(n5165) );
  IVA U21953 ( .A(n5343), .Z(n5166) );
  IVA U21954 ( .A(n5344), .Z(n5167) );
  IVA U21955 ( .A(n5344), .Z(n5168) );
  IVA U21956 ( .A(n5344), .Z(n5169) );
  IVA U21957 ( .A(n5345), .Z(n5170) );
  IVA U21958 ( .A(n5345), .Z(n5171) );
  IVA U21959 ( .A(n5345), .Z(n5172) );
  IVA U21960 ( .A(n5346), .Z(n5173) );
  IVA U21961 ( .A(n5346), .Z(n5174) );
  IVA U21962 ( .A(n5346), .Z(n5175) );
  IVA U21963 ( .A(n5347), .Z(n5176) );
  IVA U21964 ( .A(n5347), .Z(n5177) );
  IVA U21965 ( .A(n5347), .Z(n5178) );
  IVA U21966 ( .A(n5348), .Z(n5179) );
  IVA U21967 ( .A(n5348), .Z(n5180) );
  IVA U21968 ( .A(n5348), .Z(n5181) );
  IVA U21969 ( .A(n5349), .Z(n5182) );
  IVA U21970 ( .A(n5349), .Z(n5183) );
  IVA U21971 ( .A(n5349), .Z(n5184) );
  IVA U21972 ( .A(n5350), .Z(n5185) );
  IVA U21973 ( .A(n5350), .Z(n5186) );
  IVA U21974 ( .A(n5350), .Z(n5187) );
  IVA U21975 ( .A(n5351), .Z(n5188) );
  IVA U21976 ( .A(n5351), .Z(n5189) );
  IVA U21977 ( .A(n5351), .Z(n5190) );
  IVA U21978 ( .A(n5352), .Z(n5191) );
  IVA U21979 ( .A(n5352), .Z(n5192) );
  IVA U21980 ( .A(n5352), .Z(n5193) );
  IVA U21981 ( .A(n5353), .Z(n5194) );
  IVA U21982 ( .A(n5353), .Z(n5195) );
  IVA U21983 ( .A(n5353), .Z(n5196) );
  IVA U21984 ( .A(n5354), .Z(n5197) );
  IVA U21985 ( .A(n5354), .Z(n5198) );
  IVA U21986 ( .A(n5354), .Z(n5199) );
  IVA U21987 ( .A(n5355), .Z(n5200) );
  IVA U21988 ( .A(n5355), .Z(n5201) );
  IVA U21989 ( .A(n5355), .Z(n5202) );
  IVA U21990 ( .A(n5356), .Z(n5203) );
  IVA U21991 ( .A(n5356), .Z(n5204) );
  IVA U21992 ( .A(n5356), .Z(n5205) );
  IVA U21993 ( .A(n5357), .Z(n5206) );
  IVA U21994 ( .A(n5357), .Z(n5207) );
  IVA U21995 ( .A(n5357), .Z(n5208) );
  IVA U21996 ( .A(n5358), .Z(n5209) );
  IVA U21997 ( .A(n5358), .Z(n5210) );
  IVA U21998 ( .A(n5358), .Z(n5211) );
  IVA U21999 ( .A(n5359), .Z(n5212) );
  IVA U22000 ( .A(n5359), .Z(n5213) );
  IVA U22001 ( .A(n5359), .Z(n5214) );
  IVA U22002 ( .A(n5360), .Z(n5215) );
  IVA U22003 ( .A(n5360), .Z(n5216) );
  IVA U22004 ( .A(n5360), .Z(n5217) );
  IVA U22005 ( .A(n5361), .Z(n5218) );
  IVA U22006 ( .A(n5361), .Z(n5219) );
  IVA U22007 ( .A(n5361), .Z(n5220) );
  IVA U22008 ( .A(n5105), .Z(n5307) );
  IVA U22009 ( .A(n352), .Z(n5308) );
  IVA U22010 ( .A(n5113), .Z(n5309) );
  IVA U22011 ( .A(n352), .Z(n5310) );
  IVA U22012 ( .A(n352), .Z(n5311) );
  IVA U22013 ( .A(n5306), .Z(n5312) );
  IVA U22014 ( .A(n5306), .Z(n5313) );
  IVA U22015 ( .A(n5306), .Z(n5314) );
  IVA U22016 ( .A(n5306), .Z(n5315) );
  IVA U22017 ( .A(n5306), .Z(n5316) );
  IVA U22018 ( .A(n5107), .Z(n5317) );
  IVA U22019 ( .A(n5103), .Z(n5318) );
  IVA U22020 ( .A(n5101), .Z(n5319) );
  IVA U22021 ( .A(n5110), .Z(n5320) );
  IVA U22022 ( .A(n5115), .Z(n5321) );
  IVA U22023 ( .A(n5305), .Z(n5322) );
  IVA U22024 ( .A(n5305), .Z(n5323) );
  IVA U22025 ( .A(n5305), .Z(n5324) );
  IVA U22026 ( .A(n5305), .Z(n5325) );
  IVA U22027 ( .A(n5305), .Z(n5326) );
  IVA U22028 ( .A(n5304), .Z(n5327) );
  IVA U22029 ( .A(n5304), .Z(n5328) );
  IVA U22030 ( .A(n5304), .Z(n5329) );
  IVA U22031 ( .A(n5304), .Z(n5330) );
  IVA U22032 ( .A(n5304), .Z(n5331) );
  IVA U22033 ( .A(n5303), .Z(n5332) );
  IVA U22034 ( .A(n5303), .Z(n5333) );
  IVA U22035 ( .A(n5303), .Z(n5334) );
  IVA U22036 ( .A(n5303), .Z(n5335) );
  IVA U22037 ( .A(n5303), .Z(n5336) );
  IVA U22038 ( .A(n5302), .Z(n5337) );
  IVA U22039 ( .A(n5302), .Z(n5338) );
  IVA U22040 ( .A(n5302), .Z(n5339) );
  IVA U22041 ( .A(n5302), .Z(n5340) );
  IVA U22042 ( .A(n5302), .Z(n5341) );
  IVA U22043 ( .A(n5301), .Z(n5342) );
  IVA U22044 ( .A(n5301), .Z(n5343) );
  IVA U22045 ( .A(n5301), .Z(n5344) );
  IVA U22046 ( .A(n5301), .Z(n5345) );
  IVA U22047 ( .A(n5301), .Z(n5346) );
  IVA U22048 ( .A(n5300), .Z(n5347) );
  IVA U22049 ( .A(n5300), .Z(n5348) );
  IVA U22050 ( .A(n5300), .Z(n5349) );
  IVA U22051 ( .A(n5300), .Z(n5350) );
  IVA U22052 ( .A(n5300), .Z(n5351) );
  IVA U22053 ( .A(n5299), .Z(n5352) );
  IVA U22054 ( .A(n5299), .Z(n5353) );
  IVA U22055 ( .A(n5299), .Z(n5354) );
  IVA U22056 ( .A(n5299), .Z(n5355) );
  IVA U22057 ( .A(n5299), .Z(n5356) );
  IVA U22058 ( .A(n5298), .Z(n5357) );
  IVA U22059 ( .A(n5298), .Z(n5358) );
  IVA U22060 ( .A(n5298), .Z(n5359) );
  IVA U22061 ( .A(n5298), .Z(n5360) );
  IVA U22062 ( .A(n5298), .Z(n5361) );
  IVA U22063 ( .A(n5388), .Z(n5368) );
  IVA U22064 ( .A(n5388), .Z(n5369) );
  IVA U22065 ( .A(n5388), .Z(n5370) );
  IVA U22066 ( .A(n5388), .Z(n5371) );
  IVA U22067 ( .A(reset), .Z(n5388) );
  AO5 U22068 ( .A(Term1[103]), .B(Term3[15]), .C(n412), .Z(n5386) );
  IVA U22069 ( .A(n5386), .Z(n5372) );
  AO5 U22070 ( .A(Term1[104]), .B(Term3[16]), .C(n5372), .Z(n5385) );
  IVA U22071 ( .A(n5385), .Z(n5373) );
  AO5 U22072 ( .A(Term1[105]), .B(Term3[17]), .C(n5373), .Z(n5384) );
  IVA U22073 ( .A(n5384), .Z(n5374) );
  AO5 U22074 ( .A(Term1[106]), .B(Term3[18]), .C(n5374), .Z(n5383) );
  IVA U22075 ( .A(n5383), .Z(n5375) );
  AO5 U22076 ( .A(Term1[107]), .B(Term3[19]), .C(n5375), .Z(n5382) );
  IVA U22077 ( .A(n5382), .Z(n5376) );
  AO5 U22078 ( .A(Term1[108]), .B(Term3[20]), .C(n5376), .Z(n5381) );
  IVA U22079 ( .A(n5381), .Z(n5377) );
  AO5 U22080 ( .A(Term1[109]), .B(Term3[21]), .C(n5377), .Z(n5380) );
  IVA U22081 ( .A(n5380), .Z(n5378) );
  AO5 U22082 ( .A(Term1[110]), .B(Term3[22]), .C(n5378), .Z(n5379) );
  EN3P U22083 ( .A(Term1[111]), .B(Term3[23]), .C(n5379), .Z(N252) );
  EN3P U22084 ( .A(Term1[110]), .B(Term3[22]), .C(n5380), .Z(N251) );
  EN3P U22085 ( .A(Term1[109]), .B(Term3[21]), .C(n5381), .Z(N250) );
  EN3P U22086 ( .A(Term1[108]), .B(Term3[20]), .C(n5382), .Z(N249) );
  EN3P U22087 ( .A(Term1[107]), .B(Term3[19]), .C(n5383), .Z(N248) );
  EN3P U22088 ( .A(Term1[106]), .B(Term3[18]), .C(n5384), .Z(N247) );
  EN3P U22089 ( .A(Term1[105]), .B(Term3[17]), .C(n5385), .Z(N246) );
  EN3P U22090 ( .A(Term1[104]), .B(Term3[16]), .C(n5386), .Z(N245) );
  EO U22091 ( .A(Term3[15]), .B(Term1[103]), .Z(n5387) );
  EO U22092 ( .A(n412), .B(n5387), .Z(N244) );
  EO U22093 ( .A(Term3[14]), .B(Term1[102]), .Z(N243) );
  EO U22094 ( .A(Term11[118]), .B(\add_1_root_sub_1_root_add_55_2/carry[6] ), 
        .Z(N284) );
  AN2 U22095 ( .A(\add_1_root_sub_1_root_add_55_2/carry[5] ), .B(Term11[117]), 
        .Z(\add_1_root_sub_1_root_add_55_2/carry[6] ) );
  EO U22096 ( .A(Term11[117]), .B(\add_1_root_sub_1_root_add_55_2/carry[5] ), 
        .Z(N283) );
  AN2 U22097 ( .A(\add_1_root_sub_1_root_add_55_2/carry[4] ), .B(Term11[116]), 
        .Z(\add_1_root_sub_1_root_add_55_2/carry[5] ) );
  EO U22098 ( .A(Term11[116]), .B(\add_1_root_sub_1_root_add_55_2/carry[4] ), 
        .Z(N282) );
  AN2 U22099 ( .A(\add_1_root_sub_1_root_add_55_2/carry[3] ), .B(Term11[115]), 
        .Z(\add_1_root_sub_1_root_add_55_2/carry[4] ) );
  EO U22100 ( .A(Term11[115]), .B(\add_1_root_sub_1_root_add_55_2/carry[3] ), 
        .Z(N281) );
endmodule

