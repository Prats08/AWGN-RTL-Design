/* Module to calculate sin of the input signal (16,16) bits 

Func - 	0 for sine
	1 for Cosine

Latency = 1 clock cycle

*/

module SinBlock(input clk, input reset, input func, input [15:0] x, output reg [15:0] sinValue);

reg [14:0] Coeff[16384];
reg [13:0] Address;

always @(posedge clk)
begin
	if(!reset)
	begin

		case( {func, x[15:14]} )

		// Sine Calculation
	
		3'b000 : begin
				sinValue[15] <= 1'b0;
				Address = x[13:0];
				sinValue [14:0] <= Coeff [Address];  
			end

		3'b001 : begin
				sinValue[15] <= 1'b0;
				Address = (14'b1111_1111_1111_11 - x[13:0]);
				sinValue [14:0] <= Coeff [Address];
			end
	
		3'b010 : begin
				sinValue[15] <= 1'b1;
				Address = x[13:0];
				sinValue [14:0] <= Coeff [Address];
			end
	
		3'b011 : begin
				sinValue[15] <= 1'b1;
				Address = (14'b1111_1111_1111_11 - x[13:0]);
				sinValue [14:0] <= Coeff [Address];
			end

		// Cosine Calculation

		3'b100 : begin
				sinValue[15] <= 1'b0;
				Address = (14'b1111_1111_1111_11 - x[13:0]);
				sinValue [14:0] <= Coeff [Address];
			end

		3'b101 : begin
				sinValue[15] <= 1'b1;
				Address = x[13:0];
				sinValue [14:0] <= Coeff [Address];  
			end

		3'b110 : begin
				sinValue[15] <= 1'b1;
				Address = (14'b1111_1111_1111_11 - x[13:0]);
				sinValue [14:0] <= Coeff [Address];
			end
	
		3'b111 : begin
				sinValue[15] <= 1'b0;
				Address = x[13:0];
				sinValue [14:0] <= Coeff [Address];
			end	

		endcase
	end // reset

	else
	begin

		Coeff[0] <= 15'b000000000000000;
		Coeff[1] <= 15'b000000000000011;
		Coeff[2] <= 15'b000000000000110;
		Coeff[3] <= 15'b000000000001001;
		Coeff[4] <= 15'b000000000001101;
		Coeff[5] <= 15'b000000000010000;
		Coeff[6] <= 15'b000000000010011;
		Coeff[7] <= 15'b000000000010110;
		Coeff[8] <= 15'b000000000011001;
		Coeff[9] <= 15'b000000000011100;
		Coeff[10] <= 15'b000000000011111;
		Coeff[11] <= 15'b000000000100011;
		Coeff[12] <= 15'b000000000100110;
		Coeff[13] <= 15'b000000000101001;
		Coeff[14] <= 15'b000000000101100;
		Coeff[15] <= 15'b000000000101111;
		Coeff[16] <= 15'b000000000110010;
		Coeff[17] <= 15'b000000000110101;
		Coeff[18] <= 15'b000000000111001;
		Coeff[19] <= 15'b000000000111100;
		Coeff[20] <= 15'b000000000111111;
		Coeff[21] <= 15'b000000001000010;
		Coeff[22] <= 15'b000000001000101;
		Coeff[23] <= 15'b000000001001000;
		Coeff[24] <= 15'b000000001001011;
		Coeff[25] <= 15'b000000001001111;
		Coeff[26] <= 15'b000000001010010;
		Coeff[27] <= 15'b000000001010101;
		Coeff[28] <= 15'b000000001011000;
		Coeff[29] <= 15'b000000001011011;
		Coeff[30] <= 15'b000000001011110;
		Coeff[31] <= 15'b000000001100001;
		Coeff[32] <= 15'b000000001100101;
		Coeff[33] <= 15'b000000001101000;
		Coeff[34] <= 15'b000000001101011;
		Coeff[35] <= 15'b000000001101110;
		Coeff[36] <= 15'b000000001110001;
		Coeff[37] <= 15'b000000001110100;
		Coeff[38] <= 15'b000000001110111;
		Coeff[39] <= 15'b000000001111011;
		Coeff[40] <= 15'b000000001111110;
		Coeff[41] <= 15'b000000010000001;
		Coeff[42] <= 15'b000000010000100;
		Coeff[43] <= 15'b000000010000111;
		Coeff[44] <= 15'b000000010001010;
		Coeff[45] <= 15'b000000010001101;
		Coeff[46] <= 15'b000000010010001;
		Coeff[47] <= 15'b000000010010100;
		Coeff[48] <= 15'b000000010010111;
		Coeff[49] <= 15'b000000010011010;
		Coeff[50] <= 15'b000000010011101;
		Coeff[51] <= 15'b000000010100000;
		Coeff[52] <= 15'b000000010100011;
		Coeff[53] <= 15'b000000010100111;
		Coeff[54] <= 15'b000000010101010;
		Coeff[55] <= 15'b000000010101101;
		Coeff[56] <= 15'b000000010110000;
		Coeff[57] <= 15'b000000010110011;
		Coeff[58] <= 15'b000000010110110;
		Coeff[59] <= 15'b000000010111001;
		Coeff[60] <= 15'b000000010111100;
		Coeff[61] <= 15'b000000011000000;
		Coeff[62] <= 15'b000000011000011;
		Coeff[63] <= 15'b000000011000110;
		Coeff[64] <= 15'b000000011001001;
		Coeff[65] <= 15'b000000011001100;
		Coeff[66] <= 15'b000000011001111;
		Coeff[67] <= 15'b000000011010010;
		Coeff[68] <= 15'b000000011010110;
		Coeff[69] <= 15'b000000011011001;
		Coeff[70] <= 15'b000000011011100;
		Coeff[71] <= 15'b000000011011111;
		Coeff[72] <= 15'b000000011100010;
		Coeff[73] <= 15'b000000011100101;
		Coeff[74] <= 15'b000000011101000;
		Coeff[75] <= 15'b000000011101100;
		Coeff[76] <= 15'b000000011101111;
		Coeff[77] <= 15'b000000011110010;
		Coeff[78] <= 15'b000000011110101;
		Coeff[79] <= 15'b000000011111000;
		Coeff[80] <= 15'b000000011111011;
		Coeff[81] <= 15'b000000011111110;
		Coeff[82] <= 15'b000000100000010;
		Coeff[83] <= 15'b000000100000101;
		Coeff[84] <= 15'b000000100001000;
		Coeff[85] <= 15'b000000100001011;
		Coeff[86] <= 15'b000000100001110;
		Coeff[87] <= 15'b000000100010001;
		Coeff[88] <= 15'b000000100010100;
		Coeff[89] <= 15'b000000100011000;
		Coeff[90] <= 15'b000000100011011;
		Coeff[91] <= 15'b000000100011110;
		Coeff[92] <= 15'b000000100100001;
		Coeff[93] <= 15'b000000100100100;
		Coeff[94] <= 15'b000000100100111;
		Coeff[95] <= 15'b000000100101010;
		Coeff[96] <= 15'b000000100101110;
		Coeff[97] <= 15'b000000100110001;
		Coeff[98] <= 15'b000000100110100;
		Coeff[99] <= 15'b000000100110111;
		Coeff[100] <= 15'b000000100111010;
		Coeff[101] <= 15'b000000100111101;
		Coeff[102] <= 15'b000000101000000;
		Coeff[103] <= 15'b000000101000100;
		Coeff[104] <= 15'b000000101000111;
		Coeff[105] <= 15'b000000101001010;
		Coeff[106] <= 15'b000000101001101;
		Coeff[107] <= 15'b000000101010000;
		Coeff[108] <= 15'b000000101010011;
		Coeff[109] <= 15'b000000101010110;
		Coeff[110] <= 15'b000000101011010;
		Coeff[111] <= 15'b000000101011101;
		Coeff[112] <= 15'b000000101100000;
		Coeff[113] <= 15'b000000101100011;
		Coeff[114] <= 15'b000000101100110;
		Coeff[115] <= 15'b000000101101001;
		Coeff[116] <= 15'b000000101101100;
		Coeff[117] <= 15'b000000101110000;
		Coeff[118] <= 15'b000000101110011;
		Coeff[119] <= 15'b000000101110110;
		Coeff[120] <= 15'b000000101111001;
		Coeff[121] <= 15'b000000101111100;
		Coeff[122] <= 15'b000000101111111;
		Coeff[123] <= 15'b000000110000010;
		Coeff[124] <= 15'b000000110000110;
		Coeff[125] <= 15'b000000110001001;
		Coeff[126] <= 15'b000000110001100;
		Coeff[127] <= 15'b000000110001111;
		Coeff[128] <= 15'b000000110010010;
		Coeff[129] <= 15'b000000110010101;
		Coeff[130] <= 15'b000000110011000;
		Coeff[131] <= 15'b000000110011100;
		Coeff[132] <= 15'b000000110011111;
		Coeff[133] <= 15'b000000110100010;
		Coeff[134] <= 15'b000000110100101;
		Coeff[135] <= 15'b000000110101000;
		Coeff[136] <= 15'b000000110101011;
		Coeff[137] <= 15'b000000110101110;
		Coeff[138] <= 15'b000000110110010;
		Coeff[139] <= 15'b000000110110101;
		Coeff[140] <= 15'b000000110111000;
		Coeff[141] <= 15'b000000110111011;
		Coeff[142] <= 15'b000000110111110;
		Coeff[143] <= 15'b000000111000001;
		Coeff[144] <= 15'b000000111000100;
		Coeff[145] <= 15'b000000111001000;
		Coeff[146] <= 15'b000000111001011;
		Coeff[147] <= 15'b000000111001110;
		Coeff[148] <= 15'b000000111010001;
		Coeff[149] <= 15'b000000111010100;
		Coeff[150] <= 15'b000000111010111;
		Coeff[151] <= 15'b000000111011010;
		Coeff[152] <= 15'b000000111011110;
		Coeff[153] <= 15'b000000111100001;
		Coeff[154] <= 15'b000000111100100;
		Coeff[155] <= 15'b000000111100111;
		Coeff[156] <= 15'b000000111101010;
		Coeff[157] <= 15'b000000111101101;
		Coeff[158] <= 15'b000000111110000;
		Coeff[159] <= 15'b000000111110011;
		Coeff[160] <= 15'b000000111110111;
		Coeff[161] <= 15'b000000111111010;
		Coeff[162] <= 15'b000000111111101;
		Coeff[163] <= 15'b000001000000000;
		Coeff[164] <= 15'b000001000000011;
		Coeff[165] <= 15'b000001000000110;
		Coeff[166] <= 15'b000001000001001;
		Coeff[167] <= 15'b000001000001101;
		Coeff[168] <= 15'b000001000010000;
		Coeff[169] <= 15'b000001000010011;
		Coeff[170] <= 15'b000001000010110;
		Coeff[171] <= 15'b000001000011001;
		Coeff[172] <= 15'b000001000011100;
		Coeff[173] <= 15'b000001000011111;
		Coeff[174] <= 15'b000001000100011;
		Coeff[175] <= 15'b000001000100110;
		Coeff[176] <= 15'b000001000101001;
		Coeff[177] <= 15'b000001000101100;
		Coeff[178] <= 15'b000001000101111;
		Coeff[179] <= 15'b000001000110010;
		Coeff[180] <= 15'b000001000110101;
		Coeff[181] <= 15'b000001000111001;
		Coeff[182] <= 15'b000001000111100;
		Coeff[183] <= 15'b000001000111111;
		Coeff[184] <= 15'b000001001000010;
		Coeff[185] <= 15'b000001001000101;
		Coeff[186] <= 15'b000001001001000;
		Coeff[187] <= 15'b000001001001011;
		Coeff[188] <= 15'b000001001001111;
		Coeff[189] <= 15'b000001001010010;
		Coeff[190] <= 15'b000001001010101;
		Coeff[191] <= 15'b000001001011000;
		Coeff[192] <= 15'b000001001011011;
		Coeff[193] <= 15'b000001001011110;
		Coeff[194] <= 15'b000001001100001;
		Coeff[195] <= 15'b000001001100101;
		Coeff[196] <= 15'b000001001101000;
		Coeff[197] <= 15'b000001001101011;
		Coeff[198] <= 15'b000001001101110;
		Coeff[199] <= 15'b000001001110001;
		Coeff[200] <= 15'b000001001110100;
		Coeff[201] <= 15'b000001001110111;
		Coeff[202] <= 15'b000001001111011;
		Coeff[203] <= 15'b000001001111110;
		Coeff[204] <= 15'b000001010000001;
		Coeff[205] <= 15'b000001010000100;
		Coeff[206] <= 15'b000001010000111;
		Coeff[207] <= 15'b000001010001010;
		Coeff[208] <= 15'b000001010001101;
		Coeff[209] <= 15'b000001010010001;
		Coeff[210] <= 15'b000001010010100;
		Coeff[211] <= 15'b000001010010111;
		Coeff[212] <= 15'b000001010011010;
		Coeff[213] <= 15'b000001010011101;
		Coeff[214] <= 15'b000001010100000;
		Coeff[215] <= 15'b000001010100011;
		Coeff[216] <= 15'b000001010100111;
		Coeff[217] <= 15'b000001010101010;
		Coeff[218] <= 15'b000001010101101;
		Coeff[219] <= 15'b000001010110000;
		Coeff[220] <= 15'b000001010110011;
		Coeff[221] <= 15'b000001010110110;
		Coeff[222] <= 15'b000001010111001;
		Coeff[223] <= 15'b000001010111101;
		Coeff[224] <= 15'b000001011000000;
		Coeff[225] <= 15'b000001011000011;
		Coeff[226] <= 15'b000001011000110;
		Coeff[227] <= 15'b000001011001001;
		Coeff[228] <= 15'b000001011001100;
		Coeff[229] <= 15'b000001011001111;
		Coeff[230] <= 15'b000001011010011;
		Coeff[231] <= 15'b000001011010110;
		Coeff[232] <= 15'b000001011011001;
		Coeff[233] <= 15'b000001011011100;
		Coeff[234] <= 15'b000001011011111;
		Coeff[235] <= 15'b000001011100010;
		Coeff[236] <= 15'b000001011100101;
		Coeff[237] <= 15'b000001011101000;
		Coeff[238] <= 15'b000001011101100;
		Coeff[239] <= 15'b000001011101111;
		Coeff[240] <= 15'b000001011110010;
		Coeff[241] <= 15'b000001011110101;
		Coeff[242] <= 15'b000001011111000;
		Coeff[243] <= 15'b000001011111011;
		Coeff[244] <= 15'b000001011111110;
		Coeff[245] <= 15'b000001100000010;
		Coeff[246] <= 15'b000001100000101;
		Coeff[247] <= 15'b000001100001000;
		Coeff[248] <= 15'b000001100001011;
		Coeff[249] <= 15'b000001100001110;
		Coeff[250] <= 15'b000001100010001;
		Coeff[251] <= 15'b000001100010100;
		Coeff[252] <= 15'b000001100011000;
		Coeff[253] <= 15'b000001100011011;
		Coeff[254] <= 15'b000001100011110;
		Coeff[255] <= 15'b000001100100001;
		Coeff[256] <= 15'b000001100100100;
		Coeff[257] <= 15'b000001100100111;
		Coeff[258] <= 15'b000001100101010;
		Coeff[259] <= 15'b000001100101110;
		Coeff[260] <= 15'b000001100110001;
		Coeff[261] <= 15'b000001100110100;
		Coeff[262] <= 15'b000001100110111;
		Coeff[263] <= 15'b000001100111010;
		Coeff[264] <= 15'b000001100111101;
		Coeff[265] <= 15'b000001101000000;
		Coeff[266] <= 15'b000001101000100;
		Coeff[267] <= 15'b000001101000111;
		Coeff[268] <= 15'b000001101001010;
		Coeff[269] <= 15'b000001101001101;
		Coeff[270] <= 15'b000001101010000;
		Coeff[271] <= 15'b000001101010011;
		Coeff[272] <= 15'b000001101010110;
		Coeff[273] <= 15'b000001101011010;
		Coeff[274] <= 15'b000001101011101;
		Coeff[275] <= 15'b000001101100000;
		Coeff[276] <= 15'b000001101100011;
		Coeff[277] <= 15'b000001101100110;
		Coeff[278] <= 15'b000001101101001;
		Coeff[279] <= 15'b000001101101100;
		Coeff[280] <= 15'b000001101110000;
		Coeff[281] <= 15'b000001101110011;
		Coeff[282] <= 15'b000001101110110;
		Coeff[283] <= 15'b000001101111001;
		Coeff[284] <= 15'b000001101111100;
		Coeff[285] <= 15'b000001101111111;
		Coeff[286] <= 15'b000001110000010;
		Coeff[287] <= 15'b000001110000110;
		Coeff[288] <= 15'b000001110001001;
		Coeff[289] <= 15'b000001110001100;
		Coeff[290] <= 15'b000001110001111;
		Coeff[291] <= 15'b000001110010010;
		Coeff[292] <= 15'b000001110010101;
		Coeff[293] <= 15'b000001110011000;
		Coeff[294] <= 15'b000001110011100;
		Coeff[295] <= 15'b000001110011111;
		Coeff[296] <= 15'b000001110100010;
		Coeff[297] <= 15'b000001110100101;
		Coeff[298] <= 15'b000001110101000;
		Coeff[299] <= 15'b000001110101011;
		Coeff[300] <= 15'b000001110101110;
		Coeff[301] <= 15'b000001110110001;
		Coeff[302] <= 15'b000001110110101;
		Coeff[303] <= 15'b000001110111000;
		Coeff[304] <= 15'b000001110111011;
		Coeff[305] <= 15'b000001110111110;
		Coeff[306] <= 15'b000001111000001;
		Coeff[307] <= 15'b000001111000100;
		Coeff[308] <= 15'b000001111000111;
		Coeff[309] <= 15'b000001111001011;
		Coeff[310] <= 15'b000001111001110;
		Coeff[311] <= 15'b000001111010001;
		Coeff[312] <= 15'b000001111010100;
		Coeff[313] <= 15'b000001111010111;
		Coeff[314] <= 15'b000001111011010;
		Coeff[315] <= 15'b000001111011101;
		Coeff[316] <= 15'b000001111100001;
		Coeff[317] <= 15'b000001111100100;
		Coeff[318] <= 15'b000001111100111;
		Coeff[319] <= 15'b000001111101010;
		Coeff[320] <= 15'b000001111101101;
		Coeff[321] <= 15'b000001111110000;
		Coeff[322] <= 15'b000001111110011;
		Coeff[323] <= 15'b000001111110111;
		Coeff[324] <= 15'b000001111111010;
		Coeff[325] <= 15'b000001111111101;
		Coeff[326] <= 15'b000010000000000;
		Coeff[327] <= 15'b000010000000011;
		Coeff[328] <= 15'b000010000000110;
		Coeff[329] <= 15'b000010000001001;
		Coeff[330] <= 15'b000010000001101;
		Coeff[331] <= 15'b000010000010000;
		Coeff[332] <= 15'b000010000010011;
		Coeff[333] <= 15'b000010000010110;
		Coeff[334] <= 15'b000010000011001;
		Coeff[335] <= 15'b000010000011100;
		Coeff[336] <= 15'b000010000011111;
		Coeff[337] <= 15'b000010000100011;
		Coeff[338] <= 15'b000010000100110;
		Coeff[339] <= 15'b000010000101001;
		Coeff[340] <= 15'b000010000101100;
		Coeff[341] <= 15'b000010000101111;
		Coeff[342] <= 15'b000010000110010;
		Coeff[343] <= 15'b000010000110101;
		Coeff[344] <= 15'b000010000111001;
		Coeff[345] <= 15'b000010000111100;
		Coeff[346] <= 15'b000010000111111;
		Coeff[347] <= 15'b000010001000010;
		Coeff[348] <= 15'b000010001000101;
		Coeff[349] <= 15'b000010001001000;
		Coeff[350] <= 15'b000010001001011;
		Coeff[351] <= 15'b000010001001110;
		Coeff[352] <= 15'b000010001010010;
		Coeff[353] <= 15'b000010001010101;
		Coeff[354] <= 15'b000010001011000;
		Coeff[355] <= 15'b000010001011011;
		Coeff[356] <= 15'b000010001011110;
		Coeff[357] <= 15'b000010001100001;
		Coeff[358] <= 15'b000010001100100;
		Coeff[359] <= 15'b000010001101000;
		Coeff[360] <= 15'b000010001101011;
		Coeff[361] <= 15'b000010001101110;
		Coeff[362] <= 15'b000010001110001;
		Coeff[363] <= 15'b000010001110100;
		Coeff[364] <= 15'b000010001110111;
		Coeff[365] <= 15'b000010001111010;
		Coeff[366] <= 15'b000010001111110;
		Coeff[367] <= 15'b000010010000001;
		Coeff[368] <= 15'b000010010000100;
		Coeff[369] <= 15'b000010010000111;
		Coeff[370] <= 15'b000010010001010;
		Coeff[371] <= 15'b000010010001101;
		Coeff[372] <= 15'b000010010010000;
		Coeff[373] <= 15'b000010010010100;
		Coeff[374] <= 15'b000010010010111;
		Coeff[375] <= 15'b000010010011010;
		Coeff[376] <= 15'b000010010011101;
		Coeff[377] <= 15'b000010010100000;
		Coeff[378] <= 15'b000010010100011;
		Coeff[379] <= 15'b000010010100110;
		Coeff[380] <= 15'b000010010101010;
		Coeff[381] <= 15'b000010010101101;
		Coeff[382] <= 15'b000010010110000;
		Coeff[383] <= 15'b000010010110011;
		Coeff[384] <= 15'b000010010110110;
		Coeff[385] <= 15'b000010010111001;
		Coeff[386] <= 15'b000010010111100;
		Coeff[387] <= 15'b000010011000000;
		Coeff[388] <= 15'b000010011000011;
		Coeff[389] <= 15'b000010011000110;
		Coeff[390] <= 15'b000010011001001;
		Coeff[391] <= 15'b000010011001100;
		Coeff[392] <= 15'b000010011001111;
		Coeff[393] <= 15'b000010011010010;
		Coeff[394] <= 15'b000010011010101;
		Coeff[395] <= 15'b000010011011001;
		Coeff[396] <= 15'b000010011011100;
		Coeff[397] <= 15'b000010011011111;
		Coeff[398] <= 15'b000010011100010;
		Coeff[399] <= 15'b000010011100101;
		Coeff[400] <= 15'b000010011101000;
		Coeff[401] <= 15'b000010011101011;
		Coeff[402] <= 15'b000010011101111;
		Coeff[403] <= 15'b000010011110010;
		Coeff[404] <= 15'b000010011110101;
		Coeff[405] <= 15'b000010011111000;
		Coeff[406] <= 15'b000010011111011;
		Coeff[407] <= 15'b000010011111110;
		Coeff[408] <= 15'b000010100000001;
		Coeff[409] <= 15'b000010100000101;
		Coeff[410] <= 15'b000010100001000;
		Coeff[411] <= 15'b000010100001011;
		Coeff[412] <= 15'b000010100001110;
		Coeff[413] <= 15'b000010100010001;
		Coeff[414] <= 15'b000010100010100;
		Coeff[415] <= 15'b000010100010111;
		Coeff[416] <= 15'b000010100011011;
		Coeff[417] <= 15'b000010100011110;
		Coeff[418] <= 15'b000010100100001;
		Coeff[419] <= 15'b000010100100100;
		Coeff[420] <= 15'b000010100100111;
		Coeff[421] <= 15'b000010100101010;
		Coeff[422] <= 15'b000010100101101;
		Coeff[423] <= 15'b000010100110001;
		Coeff[424] <= 15'b000010100110100;
		Coeff[425] <= 15'b000010100110111;
		Coeff[426] <= 15'b000010100111010;
		Coeff[427] <= 15'b000010100111101;
		Coeff[428] <= 15'b000010101000000;
		Coeff[429] <= 15'b000010101000011;
		Coeff[430] <= 15'b000010101000111;
		Coeff[431] <= 15'b000010101001010;
		Coeff[432] <= 15'b000010101001101;
		Coeff[433] <= 15'b000010101010000;
		Coeff[434] <= 15'b000010101010011;
		Coeff[435] <= 15'b000010101010110;
		Coeff[436] <= 15'b000010101011001;
		Coeff[437] <= 15'b000010101011100;
		Coeff[438] <= 15'b000010101100000;
		Coeff[439] <= 15'b000010101100011;
		Coeff[440] <= 15'b000010101100110;
		Coeff[441] <= 15'b000010101101001;
		Coeff[442] <= 15'b000010101101100;
		Coeff[443] <= 15'b000010101101111;
		Coeff[444] <= 15'b000010101110010;
		Coeff[445] <= 15'b000010101110110;
		Coeff[446] <= 15'b000010101111001;
		Coeff[447] <= 15'b000010101111100;
		Coeff[448] <= 15'b000010101111111;
		Coeff[449] <= 15'b000010110000010;
		Coeff[450] <= 15'b000010110000101;
		Coeff[451] <= 15'b000010110001000;
		Coeff[452] <= 15'b000010110001100;
		Coeff[453] <= 15'b000010110001111;
		Coeff[454] <= 15'b000010110010010;
		Coeff[455] <= 15'b000010110010101;
		Coeff[456] <= 15'b000010110011000;
		Coeff[457] <= 15'b000010110011011;
		Coeff[458] <= 15'b000010110011110;
		Coeff[459] <= 15'b000010110100010;
		Coeff[460] <= 15'b000010110100101;
		Coeff[461] <= 15'b000010110101000;
		Coeff[462] <= 15'b000010110101011;
		Coeff[463] <= 15'b000010110101110;
		Coeff[464] <= 15'b000010110110001;
		Coeff[465] <= 15'b000010110110100;
		Coeff[466] <= 15'b000010110110111;
		Coeff[467] <= 15'b000010110111011;
		Coeff[468] <= 15'b000010110111110;
		Coeff[469] <= 15'b000010111000001;
		Coeff[470] <= 15'b000010111000100;
		Coeff[471] <= 15'b000010111000111;
		Coeff[472] <= 15'b000010111001010;
		Coeff[473] <= 15'b000010111001101;
		Coeff[474] <= 15'b000010111010001;
		Coeff[475] <= 15'b000010111010100;
		Coeff[476] <= 15'b000010111010111;
		Coeff[477] <= 15'b000010111011010;
		Coeff[478] <= 15'b000010111011101;
		Coeff[479] <= 15'b000010111100000;
		Coeff[480] <= 15'b000010111100011;
		Coeff[481] <= 15'b000010111100111;
		Coeff[482] <= 15'b000010111101010;
		Coeff[483] <= 15'b000010111101101;
		Coeff[484] <= 15'b000010111110000;
		Coeff[485] <= 15'b000010111110011;
		Coeff[486] <= 15'b000010111110110;
		Coeff[487] <= 15'b000010111111001;
		Coeff[488] <= 15'b000010111111101;
		Coeff[489] <= 15'b000011000000000;
		Coeff[490] <= 15'b000011000000011;
		Coeff[491] <= 15'b000011000000110;
		Coeff[492] <= 15'b000011000001001;
		Coeff[493] <= 15'b000011000001100;
		Coeff[494] <= 15'b000011000001111;
		Coeff[495] <= 15'b000011000010011;
		Coeff[496] <= 15'b000011000010110;
		Coeff[497] <= 15'b000011000011001;
		Coeff[498] <= 15'b000011000011100;
		Coeff[499] <= 15'b000011000011111;
		Coeff[500] <= 15'b000011000100010;
		Coeff[501] <= 15'b000011000100101;
		Coeff[502] <= 15'b000011000101000;
		Coeff[503] <= 15'b000011000101100;
		Coeff[504] <= 15'b000011000101111;
		Coeff[505] <= 15'b000011000110010;
		Coeff[506] <= 15'b000011000110101;
		Coeff[507] <= 15'b000011000111000;
		Coeff[508] <= 15'b000011000111011;
		Coeff[509] <= 15'b000011000111110;
		Coeff[510] <= 15'b000011001000010;
		Coeff[511] <= 15'b000011001000101;
		Coeff[512] <= 15'b000011001001000;
		Coeff[513] <= 15'b000011001001011;
		Coeff[514] <= 15'b000011001001110;
		Coeff[515] <= 15'b000011001010001;
		Coeff[516] <= 15'b000011001010100;
		Coeff[517] <= 15'b000011001011000;
		Coeff[518] <= 15'b000011001011011;
		Coeff[519] <= 15'b000011001011110;
		Coeff[520] <= 15'b000011001100001;
		Coeff[521] <= 15'b000011001100100;
		Coeff[522] <= 15'b000011001100111;
		Coeff[523] <= 15'b000011001101010;
		Coeff[524] <= 15'b000011001101110;
		Coeff[525] <= 15'b000011001110001;
		Coeff[526] <= 15'b000011001110100;
		Coeff[527] <= 15'b000011001110111;
		Coeff[528] <= 15'b000011001111010;
		Coeff[529] <= 15'b000011001111101;
		Coeff[530] <= 15'b000011010000000;
		Coeff[531] <= 15'b000011010000011;
		Coeff[532] <= 15'b000011010000111;
		Coeff[533] <= 15'b000011010001010;
		Coeff[534] <= 15'b000011010001101;
		Coeff[535] <= 15'b000011010010000;
		Coeff[536] <= 15'b000011010010011;
		Coeff[537] <= 15'b000011010010110;
		Coeff[538] <= 15'b000011010011001;
		Coeff[539] <= 15'b000011010011101;
		Coeff[540] <= 15'b000011010100000;
		Coeff[541] <= 15'b000011010100011;
		Coeff[542] <= 15'b000011010100110;
		Coeff[543] <= 15'b000011010101001;
		Coeff[544] <= 15'b000011010101100;
		Coeff[545] <= 15'b000011010101111;
		Coeff[546] <= 15'b000011010110011;
		Coeff[547] <= 15'b000011010110110;
		Coeff[548] <= 15'b000011010111001;
		Coeff[549] <= 15'b000011010111100;
		Coeff[550] <= 15'b000011010111111;
		Coeff[551] <= 15'b000011011000010;
		Coeff[552] <= 15'b000011011000101;
		Coeff[553] <= 15'b000011011001000;
		Coeff[554] <= 15'b000011011001100;
		Coeff[555] <= 15'b000011011001111;
		Coeff[556] <= 15'b000011011010010;
		Coeff[557] <= 15'b000011011010101;
		Coeff[558] <= 15'b000011011011000;
		Coeff[559] <= 15'b000011011011011;
		Coeff[560] <= 15'b000011011011110;
		Coeff[561] <= 15'b000011011100010;
		Coeff[562] <= 15'b000011011100101;
		Coeff[563] <= 15'b000011011101000;
		Coeff[564] <= 15'b000011011101011;
		Coeff[565] <= 15'b000011011101110;
		Coeff[566] <= 15'b000011011110001;
		Coeff[567] <= 15'b000011011110100;
		Coeff[568] <= 15'b000011011111000;
		Coeff[569] <= 15'b000011011111011;
		Coeff[570] <= 15'b000011011111110;
		Coeff[571] <= 15'b000011100000001;
		Coeff[572] <= 15'b000011100000100;
		Coeff[573] <= 15'b000011100000111;
		Coeff[574] <= 15'b000011100001010;
		Coeff[575] <= 15'b000011100001110;
		Coeff[576] <= 15'b000011100010001;
		Coeff[577] <= 15'b000011100010100;
		Coeff[578] <= 15'b000011100010111;
		Coeff[579] <= 15'b000011100011010;
		Coeff[580] <= 15'b000011100011101;
		Coeff[581] <= 15'b000011100100000;
		Coeff[582] <= 15'b000011100100011;
		Coeff[583] <= 15'b000011100100111;
		Coeff[584] <= 15'b000011100101010;
		Coeff[585] <= 15'b000011100101101;
		Coeff[586] <= 15'b000011100110000;
		Coeff[587] <= 15'b000011100110011;
		Coeff[588] <= 15'b000011100110110;
		Coeff[589] <= 15'b000011100111001;
		Coeff[590] <= 15'b000011100111101;
		Coeff[591] <= 15'b000011101000000;
		Coeff[592] <= 15'b000011101000011;
		Coeff[593] <= 15'b000011101000110;
		Coeff[594] <= 15'b000011101001001;
		Coeff[595] <= 15'b000011101001100;
		Coeff[596] <= 15'b000011101001111;
		Coeff[597] <= 15'b000011101010011;
		Coeff[598] <= 15'b000011101010110;
		Coeff[599] <= 15'b000011101011001;
		Coeff[600] <= 15'b000011101011100;
		Coeff[601] <= 15'b000011101011111;
		Coeff[602] <= 15'b000011101100010;
		Coeff[603] <= 15'b000011101100101;
		Coeff[604] <= 15'b000011101101000;
		Coeff[605] <= 15'b000011101101100;
		Coeff[606] <= 15'b000011101101111;
		Coeff[607] <= 15'b000011101110010;
		Coeff[608] <= 15'b000011101110101;
		Coeff[609] <= 15'b000011101111000;
		Coeff[610] <= 15'b000011101111011;
		Coeff[611] <= 15'b000011101111110;
		Coeff[612] <= 15'b000011110000010;
		Coeff[613] <= 15'b000011110000101;
		Coeff[614] <= 15'b000011110001000;
		Coeff[615] <= 15'b000011110001011;
		Coeff[616] <= 15'b000011110001110;
		Coeff[617] <= 15'b000011110010001;
		Coeff[618] <= 15'b000011110010100;
		Coeff[619] <= 15'b000011110011000;
		Coeff[620] <= 15'b000011110011011;
		Coeff[621] <= 15'b000011110011110;
		Coeff[622] <= 15'b000011110100001;
		Coeff[623] <= 15'b000011110100100;
		Coeff[624] <= 15'b000011110100111;
		Coeff[625] <= 15'b000011110101010;
		Coeff[626] <= 15'b000011110101101;
		Coeff[627] <= 15'b000011110110001;
		Coeff[628] <= 15'b000011110110100;
		Coeff[629] <= 15'b000011110110111;
		Coeff[630] <= 15'b000011110111010;
		Coeff[631] <= 15'b000011110111101;
		Coeff[632] <= 15'b000011111000000;
		Coeff[633] <= 15'b000011111000011;
		Coeff[634] <= 15'b000011111000111;
		Coeff[635] <= 15'b000011111001010;
		Coeff[636] <= 15'b000011111001101;
		Coeff[637] <= 15'b000011111010000;
		Coeff[638] <= 15'b000011111010011;
		Coeff[639] <= 15'b000011111010110;
		Coeff[640] <= 15'b000011111011001;
		Coeff[641] <= 15'b000011111011100;
		Coeff[642] <= 15'b000011111100000;
		Coeff[643] <= 15'b000011111100011;
		Coeff[644] <= 15'b000011111100110;
		Coeff[645] <= 15'b000011111101001;
		Coeff[646] <= 15'b000011111101100;
		Coeff[647] <= 15'b000011111101111;
		Coeff[648] <= 15'b000011111110010;
		Coeff[649] <= 15'b000011111110110;
		Coeff[650] <= 15'b000011111111001;
		Coeff[651] <= 15'b000011111111100;
		Coeff[652] <= 15'b000011111111111;
		Coeff[653] <= 15'b000100000000010;
		Coeff[654] <= 15'b000100000000101;
		Coeff[655] <= 15'b000100000001000;
		Coeff[656] <= 15'b000100000001100;
		Coeff[657] <= 15'b000100000001111;
		Coeff[658] <= 15'b000100000010010;
		Coeff[659] <= 15'b000100000010101;
		Coeff[660] <= 15'b000100000011000;
		Coeff[661] <= 15'b000100000011011;
		Coeff[662] <= 15'b000100000011110;
		Coeff[663] <= 15'b000100000100001;
		Coeff[664] <= 15'b000100000100101;
		Coeff[665] <= 15'b000100000101000;
		Coeff[666] <= 15'b000100000101011;
		Coeff[667] <= 15'b000100000101110;
		Coeff[668] <= 15'b000100000110001;
		Coeff[669] <= 15'b000100000110100;
		Coeff[670] <= 15'b000100000110111;
		Coeff[671] <= 15'b000100000111011;
		Coeff[672] <= 15'b000100000111110;
		Coeff[673] <= 15'b000100001000001;
		Coeff[674] <= 15'b000100001000100;
		Coeff[675] <= 15'b000100001000111;
		Coeff[676] <= 15'b000100001001010;
		Coeff[677] <= 15'b000100001001101;
		Coeff[678] <= 15'b000100001010001;
		Coeff[679] <= 15'b000100001010100;
		Coeff[680] <= 15'b000100001010111;
		Coeff[681] <= 15'b000100001011010;
		Coeff[682] <= 15'b000100001011101;
		Coeff[683] <= 15'b000100001100000;
		Coeff[684] <= 15'b000100001100011;
		Coeff[685] <= 15'b000100001100110;
		Coeff[686] <= 15'b000100001101010;
		Coeff[687] <= 15'b000100001101101;
		Coeff[688] <= 15'b000100001110000;
		Coeff[689] <= 15'b000100001110011;
		Coeff[690] <= 15'b000100001110110;
		Coeff[691] <= 15'b000100001111001;
		Coeff[692] <= 15'b000100001111100;
		Coeff[693] <= 15'b000100010000000;
		Coeff[694] <= 15'b000100010000011;
		Coeff[695] <= 15'b000100010000110;
		Coeff[696] <= 15'b000100010001001;
		Coeff[697] <= 15'b000100010001100;
		Coeff[698] <= 15'b000100010001111;
		Coeff[699] <= 15'b000100010010010;
		Coeff[700] <= 15'b000100010010101;
		Coeff[701] <= 15'b000100010011001;
		Coeff[702] <= 15'b000100010011100;
		Coeff[703] <= 15'b000100010011111;
		Coeff[704] <= 15'b000100010100010;
		Coeff[705] <= 15'b000100010100101;
		Coeff[706] <= 15'b000100010101000;
		Coeff[707] <= 15'b000100010101011;
		Coeff[708] <= 15'b000100010101111;
		Coeff[709] <= 15'b000100010110010;
		Coeff[710] <= 15'b000100010110101;
		Coeff[711] <= 15'b000100010111000;
		Coeff[712] <= 15'b000100010111011;
		Coeff[713] <= 15'b000100010111110;
		Coeff[714] <= 15'b000100011000001;
		Coeff[715] <= 15'b000100011000100;
		Coeff[716] <= 15'b000100011001000;
		Coeff[717] <= 15'b000100011001011;
		Coeff[718] <= 15'b000100011001110;
		Coeff[719] <= 15'b000100011010001;
		Coeff[720] <= 15'b000100011010100;
		Coeff[721] <= 15'b000100011010111;
		Coeff[722] <= 15'b000100011011010;
		Coeff[723] <= 15'b000100011011110;
		Coeff[724] <= 15'b000100011100001;
		Coeff[725] <= 15'b000100011100100;
		Coeff[726] <= 15'b000100011100111;
		Coeff[727] <= 15'b000100011101010;
		Coeff[728] <= 15'b000100011101101;
		Coeff[729] <= 15'b000100011110000;
		Coeff[730] <= 15'b000100011110011;
		Coeff[731] <= 15'b000100011110111;
		Coeff[732] <= 15'b000100011111010;
		Coeff[733] <= 15'b000100011111101;
		Coeff[734] <= 15'b000100100000000;
		Coeff[735] <= 15'b000100100000011;
		Coeff[736] <= 15'b000100100000110;
		Coeff[737] <= 15'b000100100001001;
		Coeff[738] <= 15'b000100100001101;
		Coeff[739] <= 15'b000100100010000;
		Coeff[740] <= 15'b000100100010011;
		Coeff[741] <= 15'b000100100010110;
		Coeff[742] <= 15'b000100100011001;
		Coeff[743] <= 15'b000100100011100;
		Coeff[744] <= 15'b000100100011111;
		Coeff[745] <= 15'b000100100100010;
		Coeff[746] <= 15'b000100100100110;
		Coeff[747] <= 15'b000100100101001;
		Coeff[748] <= 15'b000100100101100;
		Coeff[749] <= 15'b000100100101111;
		Coeff[750] <= 15'b000100100110010;
		Coeff[751] <= 15'b000100100110101;
		Coeff[752] <= 15'b000100100111000;
		Coeff[753] <= 15'b000100100111100;
		Coeff[754] <= 15'b000100100111111;
		Coeff[755] <= 15'b000100101000010;
		Coeff[756] <= 15'b000100101000101;
		Coeff[757] <= 15'b000100101001000;
		Coeff[758] <= 15'b000100101001011;
		Coeff[759] <= 15'b000100101001110;
		Coeff[760] <= 15'b000100101010001;
		Coeff[761] <= 15'b000100101010101;
		Coeff[762] <= 15'b000100101011000;
		Coeff[763] <= 15'b000100101011011;
		Coeff[764] <= 15'b000100101011110;
		Coeff[765] <= 15'b000100101100001;
		Coeff[766] <= 15'b000100101100100;
		Coeff[767] <= 15'b000100101100111;
		Coeff[768] <= 15'b000100101101011;
		Coeff[769] <= 15'b000100101101110;
		Coeff[770] <= 15'b000100101110001;
		Coeff[771] <= 15'b000100101110100;
		Coeff[772] <= 15'b000100101110111;
		Coeff[773] <= 15'b000100101111010;
		Coeff[774] <= 15'b000100101111101;
		Coeff[775] <= 15'b000100110000000;
		Coeff[776] <= 15'b000100110000100;
		Coeff[777] <= 15'b000100110000111;
		Coeff[778] <= 15'b000100110001010;
		Coeff[779] <= 15'b000100110001101;
		Coeff[780] <= 15'b000100110010000;
		Coeff[781] <= 15'b000100110010011;
		Coeff[782] <= 15'b000100110010110;
		Coeff[783] <= 15'b000100110011010;
		Coeff[784] <= 15'b000100110011101;
		Coeff[785] <= 15'b000100110100000;
		Coeff[786] <= 15'b000100110100011;
		Coeff[787] <= 15'b000100110100110;
		Coeff[788] <= 15'b000100110101001;
		Coeff[789] <= 15'b000100110101100;
		Coeff[790] <= 15'b000100110101111;
		Coeff[791] <= 15'b000100110110011;
		Coeff[792] <= 15'b000100110110110;
		Coeff[793] <= 15'b000100110111001;
		Coeff[794] <= 15'b000100110111100;
		Coeff[795] <= 15'b000100110111111;
		Coeff[796] <= 15'b000100111000010;
		Coeff[797] <= 15'b000100111000101;
		Coeff[798] <= 15'b000100111001001;
		Coeff[799] <= 15'b000100111001100;
		Coeff[800] <= 15'b000100111001111;
		Coeff[801] <= 15'b000100111010010;
		Coeff[802] <= 15'b000100111010101;
		Coeff[803] <= 15'b000100111011000;
		Coeff[804] <= 15'b000100111011011;
		Coeff[805] <= 15'b000100111011110;
		Coeff[806] <= 15'b000100111100010;
		Coeff[807] <= 15'b000100111100101;
		Coeff[808] <= 15'b000100111101000;
		Coeff[809] <= 15'b000100111101011;
		Coeff[810] <= 15'b000100111101110;
		Coeff[811] <= 15'b000100111110001;
		Coeff[812] <= 15'b000100111110100;
		Coeff[813] <= 15'b000100111111000;
		Coeff[814] <= 15'b000100111111011;
		Coeff[815] <= 15'b000100111111110;
		Coeff[816] <= 15'b000101000000001;
		Coeff[817] <= 15'b000101000000100;
		Coeff[818] <= 15'b000101000000111;
		Coeff[819] <= 15'b000101000001010;
		Coeff[820] <= 15'b000101000001101;
		Coeff[821] <= 15'b000101000010001;
		Coeff[822] <= 15'b000101000010100;
		Coeff[823] <= 15'b000101000010111;
		Coeff[824] <= 15'b000101000011010;
		Coeff[825] <= 15'b000101000011101;
		Coeff[826] <= 15'b000101000100000;
		Coeff[827] <= 15'b000101000100011;
		Coeff[828] <= 15'b000101000100111;
		Coeff[829] <= 15'b000101000101010;
		Coeff[830] <= 15'b000101000101101;
		Coeff[831] <= 15'b000101000110000;
		Coeff[832] <= 15'b000101000110011;
		Coeff[833] <= 15'b000101000110110;
		Coeff[834] <= 15'b000101000111001;
		Coeff[835] <= 15'b000101000111100;
		Coeff[836] <= 15'b000101001000000;
		Coeff[837] <= 15'b000101001000011;
		Coeff[838] <= 15'b000101001000110;
		Coeff[839] <= 15'b000101001001001;
		Coeff[840] <= 15'b000101001001100;
		Coeff[841] <= 15'b000101001001111;
		Coeff[842] <= 15'b000101001010010;
		Coeff[843] <= 15'b000101001010101;
		Coeff[844] <= 15'b000101001011001;
		Coeff[845] <= 15'b000101001011100;
		Coeff[846] <= 15'b000101001011111;
		Coeff[847] <= 15'b000101001100010;
		Coeff[848] <= 15'b000101001100101;
		Coeff[849] <= 15'b000101001101000;
		Coeff[850] <= 15'b000101001101011;
		Coeff[851] <= 15'b000101001101111;
		Coeff[852] <= 15'b000101001110010;
		Coeff[853] <= 15'b000101001110101;
		Coeff[854] <= 15'b000101001111000;
		Coeff[855] <= 15'b000101001111011;
		Coeff[856] <= 15'b000101001111110;
		Coeff[857] <= 15'b000101010000001;
		Coeff[858] <= 15'b000101010000100;
		Coeff[859] <= 15'b000101010001000;
		Coeff[860] <= 15'b000101010001011;
		Coeff[861] <= 15'b000101010001110;
		Coeff[862] <= 15'b000101010010001;
		Coeff[863] <= 15'b000101010010100;
		Coeff[864] <= 15'b000101010010111;
		Coeff[865] <= 15'b000101010011010;
		Coeff[866] <= 15'b000101010011101;
		Coeff[867] <= 15'b000101010100001;
		Coeff[868] <= 15'b000101010100100;
		Coeff[869] <= 15'b000101010100111;
		Coeff[870] <= 15'b000101010101010;
		Coeff[871] <= 15'b000101010101101;
		Coeff[872] <= 15'b000101010110000;
		Coeff[873] <= 15'b000101010110011;
		Coeff[874] <= 15'b000101010110111;
		Coeff[875] <= 15'b000101010111010;
		Coeff[876] <= 15'b000101010111101;
		Coeff[877] <= 15'b000101011000000;
		Coeff[878] <= 15'b000101011000011;
		Coeff[879] <= 15'b000101011000110;
		Coeff[880] <= 15'b000101011001001;
		Coeff[881] <= 15'b000101011001100;
		Coeff[882] <= 15'b000101011010000;
		Coeff[883] <= 15'b000101011010011;
		Coeff[884] <= 15'b000101011010110;
		Coeff[885] <= 15'b000101011011001;
		Coeff[886] <= 15'b000101011011100;
		Coeff[887] <= 15'b000101011011111;
		Coeff[888] <= 15'b000101011100010;
		Coeff[889] <= 15'b000101011100101;
		Coeff[890] <= 15'b000101011101001;
		Coeff[891] <= 15'b000101011101100;
		Coeff[892] <= 15'b000101011101111;
		Coeff[893] <= 15'b000101011110010;
		Coeff[894] <= 15'b000101011110101;
		Coeff[895] <= 15'b000101011111000;
		Coeff[896] <= 15'b000101011111011;
		Coeff[897] <= 15'b000101011111111;
		Coeff[898] <= 15'b000101100000010;
		Coeff[899] <= 15'b000101100000101;
		Coeff[900] <= 15'b000101100001000;
		Coeff[901] <= 15'b000101100001011;
		Coeff[902] <= 15'b000101100001110;
		Coeff[903] <= 15'b000101100010001;
		Coeff[904] <= 15'b000101100010100;
		Coeff[905] <= 15'b000101100011000;
		Coeff[906] <= 15'b000101100011011;
		Coeff[907] <= 15'b000101100011110;
		Coeff[908] <= 15'b000101100100001;
		Coeff[909] <= 15'b000101100100100;
		Coeff[910] <= 15'b000101100100111;
		Coeff[911] <= 15'b000101100101010;
		Coeff[912] <= 15'b000101100101101;
		Coeff[913] <= 15'b000101100110001;
		Coeff[914] <= 15'b000101100110100;
		Coeff[915] <= 15'b000101100110111;
		Coeff[916] <= 15'b000101100111010;
		Coeff[917] <= 15'b000101100111101;
		Coeff[918] <= 15'b000101101000000;
		Coeff[919] <= 15'b000101101000011;
		Coeff[920] <= 15'b000101101000111;
		Coeff[921] <= 15'b000101101001010;
		Coeff[922] <= 15'b000101101001101;
		Coeff[923] <= 15'b000101101010000;
		Coeff[924] <= 15'b000101101010011;
		Coeff[925] <= 15'b000101101010110;
		Coeff[926] <= 15'b000101101011001;
		Coeff[927] <= 15'b000101101011100;
		Coeff[928] <= 15'b000101101100000;
		Coeff[929] <= 15'b000101101100011;
		Coeff[930] <= 15'b000101101100110;
		Coeff[931] <= 15'b000101101101001;
		Coeff[932] <= 15'b000101101101100;
		Coeff[933] <= 15'b000101101101111;
		Coeff[934] <= 15'b000101101110010;
		Coeff[935] <= 15'b000101101110101;
		Coeff[936] <= 15'b000101101111001;
		Coeff[937] <= 15'b000101101111100;
		Coeff[938] <= 15'b000101101111111;
		Coeff[939] <= 15'b000101110000010;
		Coeff[940] <= 15'b000101110000101;
		Coeff[941] <= 15'b000101110001000;
		Coeff[942] <= 15'b000101110001011;
		Coeff[943] <= 15'b000101110001110;
		Coeff[944] <= 15'b000101110010010;
		Coeff[945] <= 15'b000101110010101;
		Coeff[946] <= 15'b000101110011000;
		Coeff[947] <= 15'b000101110011011;
		Coeff[948] <= 15'b000101110011110;
		Coeff[949] <= 15'b000101110100001;
		Coeff[950] <= 15'b000101110100100;
		Coeff[951] <= 15'b000101110101000;
		Coeff[952] <= 15'b000101110101011;
		Coeff[953] <= 15'b000101110101110;
		Coeff[954] <= 15'b000101110110001;
		Coeff[955] <= 15'b000101110110100;
		Coeff[956] <= 15'b000101110110111;
		Coeff[957] <= 15'b000101110111010;
		Coeff[958] <= 15'b000101110111101;
		Coeff[959] <= 15'b000101111000001;
		Coeff[960] <= 15'b000101111000100;
		Coeff[961] <= 15'b000101111000111;
		Coeff[962] <= 15'b000101111001010;
		Coeff[963] <= 15'b000101111001101;
		Coeff[964] <= 15'b000101111010000;
		Coeff[965] <= 15'b000101111010011;
		Coeff[966] <= 15'b000101111010110;
		Coeff[967] <= 15'b000101111011010;
		Coeff[968] <= 15'b000101111011101;
		Coeff[969] <= 15'b000101111100000;
		Coeff[970] <= 15'b000101111100011;
		Coeff[971] <= 15'b000101111100110;
		Coeff[972] <= 15'b000101111101001;
		Coeff[973] <= 15'b000101111101100;
		Coeff[974] <= 15'b000101111101111;
		Coeff[975] <= 15'b000101111110011;
		Coeff[976] <= 15'b000101111110110;
		Coeff[977] <= 15'b000101111111001;
		Coeff[978] <= 15'b000101111111100;
		Coeff[979] <= 15'b000101111111111;
		Coeff[980] <= 15'b000110000000010;
		Coeff[981] <= 15'b000110000000101;
		Coeff[982] <= 15'b000110000001000;
		Coeff[983] <= 15'b000110000001100;
		Coeff[984] <= 15'b000110000001111;
		Coeff[985] <= 15'b000110000010010;
		Coeff[986] <= 15'b000110000010101;
		Coeff[987] <= 15'b000110000011000;
		Coeff[988] <= 15'b000110000011011;
		Coeff[989] <= 15'b000110000011110;
		Coeff[990] <= 15'b000110000100010;
		Coeff[991] <= 15'b000110000100101;
		Coeff[992] <= 15'b000110000101000;
		Coeff[993] <= 15'b000110000101011;
		Coeff[994] <= 15'b000110000101110;
		Coeff[995] <= 15'b000110000110001;
		Coeff[996] <= 15'b000110000110100;
		Coeff[997] <= 15'b000110000110111;
		Coeff[998] <= 15'b000110000111011;
		Coeff[999] <= 15'b000110000111110;
		Coeff[1000] <= 15'b000110001000001;
		Coeff[1001] <= 15'b000110001000100;
		Coeff[1002] <= 15'b000110001000111;
		Coeff[1003] <= 15'b000110001001010;
		Coeff[1004] <= 15'b000110001001101;
		Coeff[1005] <= 15'b000110001010000;
		Coeff[1006] <= 15'b000110001010100;
		Coeff[1007] <= 15'b000110001010111;
		Coeff[1008] <= 15'b000110001011010;
		Coeff[1009] <= 15'b000110001011101;
		Coeff[1010] <= 15'b000110001100000;
		Coeff[1011] <= 15'b000110001100011;
		Coeff[1012] <= 15'b000110001100110;
		Coeff[1013] <= 15'b000110001101001;
		Coeff[1014] <= 15'b000110001101101;
		Coeff[1015] <= 15'b000110001110000;
		Coeff[1016] <= 15'b000110001110011;
		Coeff[1017] <= 15'b000110001110110;
		Coeff[1018] <= 15'b000110001111001;
		Coeff[1019] <= 15'b000110001111100;
		Coeff[1020] <= 15'b000110001111111;
		Coeff[1021] <= 15'b000110010000010;
		Coeff[1022] <= 15'b000110010000110;
		Coeff[1023] <= 15'b000110010001001;
		Coeff[1024] <= 15'b000110010001100;
		Coeff[1025] <= 15'b000110010001111;
		Coeff[1026] <= 15'b000110010010010;
		Coeff[1027] <= 15'b000110010010101;
		Coeff[1028] <= 15'b000110010011000;
		Coeff[1029] <= 15'b000110010011011;
		Coeff[1030] <= 15'b000110010011111;
		Coeff[1031] <= 15'b000110010100010;
		Coeff[1032] <= 15'b000110010100101;
		Coeff[1033] <= 15'b000110010101000;
		Coeff[1034] <= 15'b000110010101011;
		Coeff[1035] <= 15'b000110010101110;
		Coeff[1036] <= 15'b000110010110001;
		Coeff[1037] <= 15'b000110010110100;
		Coeff[1038] <= 15'b000110010111000;
		Coeff[1039] <= 15'b000110010111011;
		Coeff[1040] <= 15'b000110010111110;
		Coeff[1041] <= 15'b000110011000001;
		Coeff[1042] <= 15'b000110011000100;
		Coeff[1043] <= 15'b000110011000111;
		Coeff[1044] <= 15'b000110011001010;
		Coeff[1045] <= 15'b000110011001101;
		Coeff[1046] <= 15'b000110011010001;
		Coeff[1047] <= 15'b000110011010100;
		Coeff[1048] <= 15'b000110011010111;
		Coeff[1049] <= 15'b000110011011010;
		Coeff[1050] <= 15'b000110011011101;
		Coeff[1051] <= 15'b000110011100000;
		Coeff[1052] <= 15'b000110011100011;
		Coeff[1053] <= 15'b000110011100110;
		Coeff[1054] <= 15'b000110011101010;
		Coeff[1055] <= 15'b000110011101101;
		Coeff[1056] <= 15'b000110011110000;
		Coeff[1057] <= 15'b000110011110011;
		Coeff[1058] <= 15'b000110011110110;
		Coeff[1059] <= 15'b000110011111001;
		Coeff[1060] <= 15'b000110011111100;
		Coeff[1061] <= 15'b000110011111111;
		Coeff[1062] <= 15'b000110100000011;
		Coeff[1063] <= 15'b000110100000110;
		Coeff[1064] <= 15'b000110100001001;
		Coeff[1065] <= 15'b000110100001100;
		Coeff[1066] <= 15'b000110100001111;
		Coeff[1067] <= 15'b000110100010010;
		Coeff[1068] <= 15'b000110100010101;
		Coeff[1069] <= 15'b000110100011000;
		Coeff[1070] <= 15'b000110100011100;
		Coeff[1071] <= 15'b000110100011111;
		Coeff[1072] <= 15'b000110100100010;
		Coeff[1073] <= 15'b000110100100101;
		Coeff[1074] <= 15'b000110100101000;
		Coeff[1075] <= 15'b000110100101011;
		Coeff[1076] <= 15'b000110100101110;
		Coeff[1077] <= 15'b000110100110001;
		Coeff[1078] <= 15'b000110100110101;
		Coeff[1079] <= 15'b000110100111000;
		Coeff[1080] <= 15'b000110100111011;
		Coeff[1081] <= 15'b000110100111110;
		Coeff[1082] <= 15'b000110101000001;
		Coeff[1083] <= 15'b000110101000100;
		Coeff[1084] <= 15'b000110101000111;
		Coeff[1085] <= 15'b000110101001010;
		Coeff[1086] <= 15'b000110101001110;
		Coeff[1087] <= 15'b000110101010001;
		Coeff[1088] <= 15'b000110101010100;
		Coeff[1089] <= 15'b000110101010111;
		Coeff[1090] <= 15'b000110101011010;
		Coeff[1091] <= 15'b000110101011101;
		Coeff[1092] <= 15'b000110101100000;
		Coeff[1093] <= 15'b000110101100011;
		Coeff[1094] <= 15'b000110101100111;
		Coeff[1095] <= 15'b000110101101010;
		Coeff[1096] <= 15'b000110101101101;
		Coeff[1097] <= 15'b000110101110000;
		Coeff[1098] <= 15'b000110101110011;
		Coeff[1099] <= 15'b000110101110110;
		Coeff[1100] <= 15'b000110101111001;
		Coeff[1101] <= 15'b000110101111100;
		Coeff[1102] <= 15'b000110110000000;
		Coeff[1103] <= 15'b000110110000011;
		Coeff[1104] <= 15'b000110110000110;
		Coeff[1105] <= 15'b000110110001001;
		Coeff[1106] <= 15'b000110110001100;
		Coeff[1107] <= 15'b000110110001111;
		Coeff[1108] <= 15'b000110110010010;
		Coeff[1109] <= 15'b000110110010101;
		Coeff[1110] <= 15'b000110110011001;
		Coeff[1111] <= 15'b000110110011100;
		Coeff[1112] <= 15'b000110110011111;
		Coeff[1113] <= 15'b000110110100010;
		Coeff[1114] <= 15'b000110110100101;
		Coeff[1115] <= 15'b000110110101000;
		Coeff[1116] <= 15'b000110110101011;
		Coeff[1117] <= 15'b000110110101110;
		Coeff[1118] <= 15'b000110110110010;
		Coeff[1119] <= 15'b000110110110101;
		Coeff[1120] <= 15'b000110110111000;
		Coeff[1121] <= 15'b000110110111011;
		Coeff[1122] <= 15'b000110110111110;
		Coeff[1123] <= 15'b000110111000001;
		Coeff[1124] <= 15'b000110111000100;
		Coeff[1125] <= 15'b000110111000111;
		Coeff[1126] <= 15'b000110111001011;
		Coeff[1127] <= 15'b000110111001110;
		Coeff[1128] <= 15'b000110111010001;
		Coeff[1129] <= 15'b000110111010100;
		Coeff[1130] <= 15'b000110111010111;
		Coeff[1131] <= 15'b000110111011010;
		Coeff[1132] <= 15'b000110111011101;
		Coeff[1133] <= 15'b000110111100000;
		Coeff[1134] <= 15'b000110111100100;
		Coeff[1135] <= 15'b000110111100111;
		Coeff[1136] <= 15'b000110111101010;
		Coeff[1137] <= 15'b000110111101101;
		Coeff[1138] <= 15'b000110111110000;
		Coeff[1139] <= 15'b000110111110011;
		Coeff[1140] <= 15'b000110111110110;
		Coeff[1141] <= 15'b000110111111001;
		Coeff[1142] <= 15'b000110111111101;
		Coeff[1143] <= 15'b000111000000000;
		Coeff[1144] <= 15'b000111000000011;
		Coeff[1145] <= 15'b000111000000110;
		Coeff[1146] <= 15'b000111000001001;
		Coeff[1147] <= 15'b000111000001100;
		Coeff[1148] <= 15'b000111000001111;
		Coeff[1149] <= 15'b000111000010010;
		Coeff[1150] <= 15'b000111000010110;
		Coeff[1151] <= 15'b000111000011001;
		Coeff[1152] <= 15'b000111000011100;
		Coeff[1153] <= 15'b000111000011111;
		Coeff[1154] <= 15'b000111000100010;
		Coeff[1155] <= 15'b000111000100101;
		Coeff[1156] <= 15'b000111000101000;
		Coeff[1157] <= 15'b000111000101011;
		Coeff[1158] <= 15'b000111000101110;
		Coeff[1159] <= 15'b000111000110010;
		Coeff[1160] <= 15'b000111000110101;
		Coeff[1161] <= 15'b000111000111000;
		Coeff[1162] <= 15'b000111000111011;
		Coeff[1163] <= 15'b000111000111110;
		Coeff[1164] <= 15'b000111001000001;
		Coeff[1165] <= 15'b000111001000100;
		Coeff[1166] <= 15'b000111001000111;
		Coeff[1167] <= 15'b000111001001011;
		Coeff[1168] <= 15'b000111001001110;
		Coeff[1169] <= 15'b000111001010001;
		Coeff[1170] <= 15'b000111001010100;
		Coeff[1171] <= 15'b000111001010111;
		Coeff[1172] <= 15'b000111001011010;
		Coeff[1173] <= 15'b000111001011101;
		Coeff[1174] <= 15'b000111001100000;
		Coeff[1175] <= 15'b000111001100100;
		Coeff[1176] <= 15'b000111001100111;
		Coeff[1177] <= 15'b000111001101010;
		Coeff[1178] <= 15'b000111001101101;
		Coeff[1179] <= 15'b000111001110000;
		Coeff[1180] <= 15'b000111001110011;
		Coeff[1181] <= 15'b000111001110110;
		Coeff[1182] <= 15'b000111001111001;
		Coeff[1183] <= 15'b000111001111101;
		Coeff[1184] <= 15'b000111010000000;
		Coeff[1185] <= 15'b000111010000011;
		Coeff[1186] <= 15'b000111010000110;
		Coeff[1187] <= 15'b000111010001001;
		Coeff[1188] <= 15'b000111010001100;
		Coeff[1189] <= 15'b000111010001111;
		Coeff[1190] <= 15'b000111010010010;
		Coeff[1191] <= 15'b000111010010110;
		Coeff[1192] <= 15'b000111010011001;
		Coeff[1193] <= 15'b000111010011100;
		Coeff[1194] <= 15'b000111010011111;
		Coeff[1195] <= 15'b000111010100010;
		Coeff[1196] <= 15'b000111010100101;
		Coeff[1197] <= 15'b000111010101000;
		Coeff[1198] <= 15'b000111010101011;
		Coeff[1199] <= 15'b000111010101110;
		Coeff[1200] <= 15'b000111010110010;
		Coeff[1201] <= 15'b000111010110101;
		Coeff[1202] <= 15'b000111010111000;
		Coeff[1203] <= 15'b000111010111011;
		Coeff[1204] <= 15'b000111010111110;
		Coeff[1205] <= 15'b000111011000001;
		Coeff[1206] <= 15'b000111011000100;
		Coeff[1207] <= 15'b000111011000111;
		Coeff[1208] <= 15'b000111011001011;
		Coeff[1209] <= 15'b000111011001110;
		Coeff[1210] <= 15'b000111011010001;
		Coeff[1211] <= 15'b000111011010100;
		Coeff[1212] <= 15'b000111011010111;
		Coeff[1213] <= 15'b000111011011010;
		Coeff[1214] <= 15'b000111011011101;
		Coeff[1215] <= 15'b000111011100000;
		Coeff[1216] <= 15'b000111011100100;
		Coeff[1217] <= 15'b000111011100111;
		Coeff[1218] <= 15'b000111011101010;
		Coeff[1219] <= 15'b000111011101101;
		Coeff[1220] <= 15'b000111011110000;
		Coeff[1221] <= 15'b000111011110011;
		Coeff[1222] <= 15'b000111011110110;
		Coeff[1223] <= 15'b000111011111001;
		Coeff[1224] <= 15'b000111011111100;
		Coeff[1225] <= 15'b000111100000000;
		Coeff[1226] <= 15'b000111100000011;
		Coeff[1227] <= 15'b000111100000110;
		Coeff[1228] <= 15'b000111100001001;
		Coeff[1229] <= 15'b000111100001100;
		Coeff[1230] <= 15'b000111100001111;
		Coeff[1231] <= 15'b000111100010010;
		Coeff[1232] <= 15'b000111100010101;
		Coeff[1233] <= 15'b000111100011001;
		Coeff[1234] <= 15'b000111100011100;
		Coeff[1235] <= 15'b000111100011111;
		Coeff[1236] <= 15'b000111100100010;
		Coeff[1237] <= 15'b000111100100101;
		Coeff[1238] <= 15'b000111100101000;
		Coeff[1239] <= 15'b000111100101011;
		Coeff[1240] <= 15'b000111100101110;
		Coeff[1241] <= 15'b000111100110010;
		Coeff[1242] <= 15'b000111100110101;
		Coeff[1243] <= 15'b000111100111000;
		Coeff[1244] <= 15'b000111100111011;
		Coeff[1245] <= 15'b000111100111110;
		Coeff[1246] <= 15'b000111101000001;
		Coeff[1247] <= 15'b000111101000100;
		Coeff[1248] <= 15'b000111101000111;
		Coeff[1249] <= 15'b000111101001010;
		Coeff[1250] <= 15'b000111101001110;
		Coeff[1251] <= 15'b000111101010001;
		Coeff[1252] <= 15'b000111101010100;
		Coeff[1253] <= 15'b000111101010111;
		Coeff[1254] <= 15'b000111101011010;
		Coeff[1255] <= 15'b000111101011101;
		Coeff[1256] <= 15'b000111101100000;
		Coeff[1257] <= 15'b000111101100011;
		Coeff[1258] <= 15'b000111101100111;
		Coeff[1259] <= 15'b000111101101010;
		Coeff[1260] <= 15'b000111101101101;
		Coeff[1261] <= 15'b000111101110000;
		Coeff[1262] <= 15'b000111101110011;
		Coeff[1263] <= 15'b000111101110110;
		Coeff[1264] <= 15'b000111101111001;
		Coeff[1265] <= 15'b000111101111100;
		Coeff[1266] <= 15'b000111101111111;
		Coeff[1267] <= 15'b000111110000011;
		Coeff[1268] <= 15'b000111110000110;
		Coeff[1269] <= 15'b000111110001001;
		Coeff[1270] <= 15'b000111110001100;
		Coeff[1271] <= 15'b000111110001111;
		Coeff[1272] <= 15'b000111110010010;
		Coeff[1273] <= 15'b000111110010101;
		Coeff[1274] <= 15'b000111110011000;
		Coeff[1275] <= 15'b000111110011100;
		Coeff[1276] <= 15'b000111110011111;
		Coeff[1277] <= 15'b000111110100010;
		Coeff[1278] <= 15'b000111110100101;
		Coeff[1279] <= 15'b000111110101000;
		Coeff[1280] <= 15'b000111110101011;
		Coeff[1281] <= 15'b000111110101110;
		Coeff[1282] <= 15'b000111110110001;
		Coeff[1283] <= 15'b000111110110101;
		Coeff[1284] <= 15'b000111110111000;
		Coeff[1285] <= 15'b000111110111011;
		Coeff[1286] <= 15'b000111110111110;
		Coeff[1287] <= 15'b000111111000001;
		Coeff[1288] <= 15'b000111111000100;
		Coeff[1289] <= 15'b000111111000111;
		Coeff[1290] <= 15'b000111111001010;
		Coeff[1291] <= 15'b000111111001101;
		Coeff[1292] <= 15'b000111111010001;
		Coeff[1293] <= 15'b000111111010100;
		Coeff[1294] <= 15'b000111111010111;
		Coeff[1295] <= 15'b000111111011010;
		Coeff[1296] <= 15'b000111111011101;
		Coeff[1297] <= 15'b000111111100000;
		Coeff[1298] <= 15'b000111111100011;
		Coeff[1299] <= 15'b000111111100110;
		Coeff[1300] <= 15'b000111111101010;
		Coeff[1301] <= 15'b000111111101101;
		Coeff[1302] <= 15'b000111111110000;
		Coeff[1303] <= 15'b000111111110011;
		Coeff[1304] <= 15'b000111111110110;
		Coeff[1305] <= 15'b000111111111001;
		Coeff[1306] <= 15'b000111111111100;
		Coeff[1307] <= 15'b000111111111111;
		Coeff[1308] <= 15'b001000000000010;
		Coeff[1309] <= 15'b001000000000110;
		Coeff[1310] <= 15'b001000000001001;
		Coeff[1311] <= 15'b001000000001100;
		Coeff[1312] <= 15'b001000000001111;
		Coeff[1313] <= 15'b001000000010010;
		Coeff[1314] <= 15'b001000000010101;
		Coeff[1315] <= 15'b001000000011000;
		Coeff[1316] <= 15'b001000000011011;
		Coeff[1317] <= 15'b001000000011110;
		Coeff[1318] <= 15'b001000000100010;
		Coeff[1319] <= 15'b001000000100101;
		Coeff[1320] <= 15'b001000000101000;
		Coeff[1321] <= 15'b001000000101011;
		Coeff[1322] <= 15'b001000000101110;
		Coeff[1323] <= 15'b001000000110001;
		Coeff[1324] <= 15'b001000000110100;
		Coeff[1325] <= 15'b001000000110111;
		Coeff[1326] <= 15'b001000000111011;
		Coeff[1327] <= 15'b001000000111110;
		Coeff[1328] <= 15'b001000001000001;
		Coeff[1329] <= 15'b001000001000100;
		Coeff[1330] <= 15'b001000001000111;
		Coeff[1331] <= 15'b001000001001010;
		Coeff[1332] <= 15'b001000001001101;
		Coeff[1333] <= 15'b001000001010000;
		Coeff[1334] <= 15'b001000001010011;
		Coeff[1335] <= 15'b001000001010111;
		Coeff[1336] <= 15'b001000001011010;
		Coeff[1337] <= 15'b001000001011101;
		Coeff[1338] <= 15'b001000001100000;
		Coeff[1339] <= 15'b001000001100011;
		Coeff[1340] <= 15'b001000001100110;
		Coeff[1341] <= 15'b001000001101001;
		Coeff[1342] <= 15'b001000001101100;
		Coeff[1343] <= 15'b001000001110000;
		Coeff[1344] <= 15'b001000001110011;
		Coeff[1345] <= 15'b001000001110110;
		Coeff[1346] <= 15'b001000001111001;
		Coeff[1347] <= 15'b001000001111100;
		Coeff[1348] <= 15'b001000001111111;
		Coeff[1349] <= 15'b001000010000010;
		Coeff[1350] <= 15'b001000010000101;
		Coeff[1351] <= 15'b001000010001000;
		Coeff[1352] <= 15'b001000010001100;
		Coeff[1353] <= 15'b001000010001111;
		Coeff[1354] <= 15'b001000010010010;
		Coeff[1355] <= 15'b001000010010101;
		Coeff[1356] <= 15'b001000010011000;
		Coeff[1357] <= 15'b001000010011011;
		Coeff[1358] <= 15'b001000010011110;
		Coeff[1359] <= 15'b001000010100001;
		Coeff[1360] <= 15'b001000010100100;
		Coeff[1361] <= 15'b001000010101000;
		Coeff[1362] <= 15'b001000010101011;
		Coeff[1363] <= 15'b001000010101110;
		Coeff[1364] <= 15'b001000010110001;
		Coeff[1365] <= 15'b001000010110100;
		Coeff[1366] <= 15'b001000010110111;
		Coeff[1367] <= 15'b001000010111010;
		Coeff[1368] <= 15'b001000010111101;
		Coeff[1369] <= 15'b001000011000001;
		Coeff[1370] <= 15'b001000011000100;
		Coeff[1371] <= 15'b001000011000111;
		Coeff[1372] <= 15'b001000011001010;
		Coeff[1373] <= 15'b001000011001101;
		Coeff[1374] <= 15'b001000011010000;
		Coeff[1375] <= 15'b001000011010011;
		Coeff[1376] <= 15'b001000011010110;
		Coeff[1377] <= 15'b001000011011001;
		Coeff[1378] <= 15'b001000011011101;
		Coeff[1379] <= 15'b001000011100000;
		Coeff[1380] <= 15'b001000011100011;
		Coeff[1381] <= 15'b001000011100110;
		Coeff[1382] <= 15'b001000011101001;
		Coeff[1383] <= 15'b001000011101100;
		Coeff[1384] <= 15'b001000011101111;
		Coeff[1385] <= 15'b001000011110010;
		Coeff[1386] <= 15'b001000011110101;
		Coeff[1387] <= 15'b001000011111001;
		Coeff[1388] <= 15'b001000011111100;
		Coeff[1389] <= 15'b001000011111111;
		Coeff[1390] <= 15'b001000100000010;
		Coeff[1391] <= 15'b001000100000101;
		Coeff[1392] <= 15'b001000100001000;
		Coeff[1393] <= 15'b001000100001011;
		Coeff[1394] <= 15'b001000100001110;
		Coeff[1395] <= 15'b001000100010001;
		Coeff[1396] <= 15'b001000100010101;
		Coeff[1397] <= 15'b001000100011000;
		Coeff[1398] <= 15'b001000100011011;
		Coeff[1399] <= 15'b001000100011110;
		Coeff[1400] <= 15'b001000100100001;
		Coeff[1401] <= 15'b001000100100100;
		Coeff[1402] <= 15'b001000100100111;
		Coeff[1403] <= 15'b001000100101010;
		Coeff[1404] <= 15'b001000100101101;
		Coeff[1405] <= 15'b001000100110001;
		Coeff[1406] <= 15'b001000100110100;
		Coeff[1407] <= 15'b001000100110111;
		Coeff[1408] <= 15'b001000100111010;
		Coeff[1409] <= 15'b001000100111101;
		Coeff[1410] <= 15'b001000101000000;
		Coeff[1411] <= 15'b001000101000011;
		Coeff[1412] <= 15'b001000101000110;
		Coeff[1413] <= 15'b001000101001010;
		Coeff[1414] <= 15'b001000101001101;
		Coeff[1415] <= 15'b001000101010000;
		Coeff[1416] <= 15'b001000101010011;
		Coeff[1417] <= 15'b001000101010110;
		Coeff[1418] <= 15'b001000101011001;
		Coeff[1419] <= 15'b001000101011100;
		Coeff[1420] <= 15'b001000101011111;
		Coeff[1421] <= 15'b001000101100010;
		Coeff[1422] <= 15'b001000101100110;
		Coeff[1423] <= 15'b001000101101001;
		Coeff[1424] <= 15'b001000101101100;
		Coeff[1425] <= 15'b001000101101111;
		Coeff[1426] <= 15'b001000101110010;
		Coeff[1427] <= 15'b001000101110101;
		Coeff[1428] <= 15'b001000101111000;
		Coeff[1429] <= 15'b001000101111011;
		Coeff[1430] <= 15'b001000101111110;
		Coeff[1431] <= 15'b001000110000010;
		Coeff[1432] <= 15'b001000110000101;
		Coeff[1433] <= 15'b001000110001000;
		Coeff[1434] <= 15'b001000110001011;
		Coeff[1435] <= 15'b001000110001110;
		Coeff[1436] <= 15'b001000110010001;
		Coeff[1437] <= 15'b001000110010100;
		Coeff[1438] <= 15'b001000110010111;
		Coeff[1439] <= 15'b001000110011010;
		Coeff[1440] <= 15'b001000110011110;
		Coeff[1441] <= 15'b001000110100001;
		Coeff[1442] <= 15'b001000110100100;
		Coeff[1443] <= 15'b001000110100111;
		Coeff[1444] <= 15'b001000110101010;
		Coeff[1445] <= 15'b001000110101101;
		Coeff[1446] <= 15'b001000110110000;
		Coeff[1447] <= 15'b001000110110011;
		Coeff[1448] <= 15'b001000110110110;
		Coeff[1449] <= 15'b001000110111010;
		Coeff[1450] <= 15'b001000110111101;
		Coeff[1451] <= 15'b001000111000000;
		Coeff[1452] <= 15'b001000111000011;
		Coeff[1453] <= 15'b001000111000110;
		Coeff[1454] <= 15'b001000111001001;
		Coeff[1455] <= 15'b001000111001100;
		Coeff[1456] <= 15'b001000111001111;
		Coeff[1457] <= 15'b001000111010010;
		Coeff[1458] <= 15'b001000111010110;
		Coeff[1459] <= 15'b001000111011001;
		Coeff[1460] <= 15'b001000111011100;
		Coeff[1461] <= 15'b001000111011111;
		Coeff[1462] <= 15'b001000111100010;
		Coeff[1463] <= 15'b001000111100101;
		Coeff[1464] <= 15'b001000111101000;
		Coeff[1465] <= 15'b001000111101011;
		Coeff[1466] <= 15'b001000111101110;
		Coeff[1467] <= 15'b001000111110010;
		Coeff[1468] <= 15'b001000111110101;
		Coeff[1469] <= 15'b001000111111000;
		Coeff[1470] <= 15'b001000111111011;
		Coeff[1471] <= 15'b001000111111110;
		Coeff[1472] <= 15'b001001000000001;
		Coeff[1473] <= 15'b001001000000100;
		Coeff[1474] <= 15'b001001000000111;
		Coeff[1475] <= 15'b001001000001010;
		Coeff[1476] <= 15'b001001000001110;
		Coeff[1477] <= 15'b001001000010001;
		Coeff[1478] <= 15'b001001000010100;
		Coeff[1479] <= 15'b001001000010111;
		Coeff[1480] <= 15'b001001000011010;
		Coeff[1481] <= 15'b001001000011101;
		Coeff[1482] <= 15'b001001000100000;
		Coeff[1483] <= 15'b001001000100011;
		Coeff[1484] <= 15'b001001000100110;
		Coeff[1485] <= 15'b001001000101010;
		Coeff[1486] <= 15'b001001000101101;
		Coeff[1487] <= 15'b001001000110000;
		Coeff[1488] <= 15'b001001000110011;
		Coeff[1489] <= 15'b001001000110110;
		Coeff[1490] <= 15'b001001000111001;
		Coeff[1491] <= 15'b001001000111100;
		Coeff[1492] <= 15'b001001000111111;
		Coeff[1493] <= 15'b001001001000010;
		Coeff[1494] <= 15'b001001001000110;
		Coeff[1495] <= 15'b001001001001001;
		Coeff[1496] <= 15'b001001001001100;
		Coeff[1497] <= 15'b001001001001111;
		Coeff[1498] <= 15'b001001001010010;
		Coeff[1499] <= 15'b001001001010101;
		Coeff[1500] <= 15'b001001001011000;
		Coeff[1501] <= 15'b001001001011011;
		Coeff[1502] <= 15'b001001001011110;
		Coeff[1503] <= 15'b001001001100001;
		Coeff[1504] <= 15'b001001001100101;
		Coeff[1505] <= 15'b001001001101000;
		Coeff[1506] <= 15'b001001001101011;
		Coeff[1507] <= 15'b001001001101110;
		Coeff[1508] <= 15'b001001001110001;
		Coeff[1509] <= 15'b001001001110100;
		Coeff[1510] <= 15'b001001001110111;
		Coeff[1511] <= 15'b001001001111010;
		Coeff[1512] <= 15'b001001001111101;
		Coeff[1513] <= 15'b001001010000001;
		Coeff[1514] <= 15'b001001010000100;
		Coeff[1515] <= 15'b001001010000111;
		Coeff[1516] <= 15'b001001010001010;
		Coeff[1517] <= 15'b001001010001101;
		Coeff[1518] <= 15'b001001010010000;
		Coeff[1519] <= 15'b001001010010011;
		Coeff[1520] <= 15'b001001010010110;
		Coeff[1521] <= 15'b001001010011001;
		Coeff[1522] <= 15'b001001010011101;
		Coeff[1523] <= 15'b001001010100000;
		Coeff[1524] <= 15'b001001010100011;
		Coeff[1525] <= 15'b001001010100110;
		Coeff[1526] <= 15'b001001010101001;
		Coeff[1527] <= 15'b001001010101100;
		Coeff[1528] <= 15'b001001010101111;
		Coeff[1529] <= 15'b001001010110010;
		Coeff[1530] <= 15'b001001010110101;
		Coeff[1531] <= 15'b001001010111001;
		Coeff[1532] <= 15'b001001010111100;
		Coeff[1533] <= 15'b001001010111111;
		Coeff[1534] <= 15'b001001011000010;
		Coeff[1535] <= 15'b001001011000101;
		Coeff[1536] <= 15'b001001011001000;
		Coeff[1537] <= 15'b001001011001011;
		Coeff[1538] <= 15'b001001011001110;
		Coeff[1539] <= 15'b001001011010001;
		Coeff[1540] <= 15'b001001011010100;
		Coeff[1541] <= 15'b001001011011000;
		Coeff[1542] <= 15'b001001011011011;
		Coeff[1543] <= 15'b001001011011110;
		Coeff[1544] <= 15'b001001011100001;
		Coeff[1545] <= 15'b001001011100100;
		Coeff[1546] <= 15'b001001011100111;
		Coeff[1547] <= 15'b001001011101010;
		Coeff[1548] <= 15'b001001011101101;
		Coeff[1549] <= 15'b001001011110000;
		Coeff[1550] <= 15'b001001011110100;
		Coeff[1551] <= 15'b001001011110111;
		Coeff[1552] <= 15'b001001011111010;
		Coeff[1553] <= 15'b001001011111101;
		Coeff[1554] <= 15'b001001100000000;
		Coeff[1555] <= 15'b001001100000011;
		Coeff[1556] <= 15'b001001100000110;
		Coeff[1557] <= 15'b001001100001001;
		Coeff[1558] <= 15'b001001100001100;
		Coeff[1559] <= 15'b001001100010000;
		Coeff[1560] <= 15'b001001100010011;
		Coeff[1561] <= 15'b001001100010110;
		Coeff[1562] <= 15'b001001100011001;
		Coeff[1563] <= 15'b001001100011100;
		Coeff[1564] <= 15'b001001100011111;
		Coeff[1565] <= 15'b001001100100010;
		Coeff[1566] <= 15'b001001100100101;
		Coeff[1567] <= 15'b001001100101000;
		Coeff[1568] <= 15'b001001100101011;
		Coeff[1569] <= 15'b001001100101111;
		Coeff[1570] <= 15'b001001100110010;
		Coeff[1571] <= 15'b001001100110101;
		Coeff[1572] <= 15'b001001100111000;
		Coeff[1573] <= 15'b001001100111011;
		Coeff[1574] <= 15'b001001100111110;
		Coeff[1575] <= 15'b001001101000001;
		Coeff[1576] <= 15'b001001101000100;
		Coeff[1577] <= 15'b001001101000111;
		Coeff[1578] <= 15'b001001101001011;
		Coeff[1579] <= 15'b001001101001110;
		Coeff[1580] <= 15'b001001101010001;
		Coeff[1581] <= 15'b001001101010100;
		Coeff[1582] <= 15'b001001101010111;
		Coeff[1583] <= 15'b001001101011010;
		Coeff[1584] <= 15'b001001101011101;
		Coeff[1585] <= 15'b001001101100000;
		Coeff[1586] <= 15'b001001101100011;
		Coeff[1587] <= 15'b001001101100110;
		Coeff[1588] <= 15'b001001101101010;
		Coeff[1589] <= 15'b001001101101101;
		Coeff[1590] <= 15'b001001101110000;
		Coeff[1591] <= 15'b001001101110011;
		Coeff[1592] <= 15'b001001101110110;
		Coeff[1593] <= 15'b001001101111001;
		Coeff[1594] <= 15'b001001101111100;
		Coeff[1595] <= 15'b001001101111111;
		Coeff[1596] <= 15'b001001110000010;
		Coeff[1597] <= 15'b001001110000110;
		Coeff[1598] <= 15'b001001110001001;
		Coeff[1599] <= 15'b001001110001100;
		Coeff[1600] <= 15'b001001110001111;
		Coeff[1601] <= 15'b001001110010010;
		Coeff[1602] <= 15'b001001110010101;
		Coeff[1603] <= 15'b001001110011000;
		Coeff[1604] <= 15'b001001110011011;
		Coeff[1605] <= 15'b001001110011110;
		Coeff[1606] <= 15'b001001110100001;
		Coeff[1607] <= 15'b001001110100101;
		Coeff[1608] <= 15'b001001110101000;
		Coeff[1609] <= 15'b001001110101011;
		Coeff[1610] <= 15'b001001110101110;
		Coeff[1611] <= 15'b001001110110001;
		Coeff[1612] <= 15'b001001110110100;
		Coeff[1613] <= 15'b001001110110111;
		Coeff[1614] <= 15'b001001110111010;
		Coeff[1615] <= 15'b001001110111101;
		Coeff[1616] <= 15'b001001111000001;
		Coeff[1617] <= 15'b001001111000100;
		Coeff[1618] <= 15'b001001111000111;
		Coeff[1619] <= 15'b001001111001010;
		Coeff[1620] <= 15'b001001111001101;
		Coeff[1621] <= 15'b001001111010000;
		Coeff[1622] <= 15'b001001111010011;
		Coeff[1623] <= 15'b001001111010110;
		Coeff[1624] <= 15'b001001111011001;
		Coeff[1625] <= 15'b001001111011100;
		Coeff[1626] <= 15'b001001111100000;
		Coeff[1627] <= 15'b001001111100011;
		Coeff[1628] <= 15'b001001111100110;
		Coeff[1629] <= 15'b001001111101001;
		Coeff[1630] <= 15'b001001111101100;
		Coeff[1631] <= 15'b001001111101111;
		Coeff[1632] <= 15'b001001111110010;
		Coeff[1633] <= 15'b001001111110101;
		Coeff[1634] <= 15'b001001111111000;
		Coeff[1635] <= 15'b001001111111011;
		Coeff[1636] <= 15'b001001111111111;
		Coeff[1637] <= 15'b001010000000010;
		Coeff[1638] <= 15'b001010000000101;
		Coeff[1639] <= 15'b001010000001000;
		Coeff[1640] <= 15'b001010000001011;
		Coeff[1641] <= 15'b001010000001110;
		Coeff[1642] <= 15'b001010000010001;
		Coeff[1643] <= 15'b001010000010100;
		Coeff[1644] <= 15'b001010000010111;
		Coeff[1645] <= 15'b001010000011011;
		Coeff[1646] <= 15'b001010000011110;
		Coeff[1647] <= 15'b001010000100001;
		Coeff[1648] <= 15'b001010000100100;
		Coeff[1649] <= 15'b001010000100111;
		Coeff[1650] <= 15'b001010000101010;
		Coeff[1651] <= 15'b001010000101101;
		Coeff[1652] <= 15'b001010000110000;
		Coeff[1653] <= 15'b001010000110011;
		Coeff[1654] <= 15'b001010000110110;
		Coeff[1655] <= 15'b001010000111010;
		Coeff[1656] <= 15'b001010000111101;
		Coeff[1657] <= 15'b001010001000000;
		Coeff[1658] <= 15'b001010001000011;
		Coeff[1659] <= 15'b001010001000110;
		Coeff[1660] <= 15'b001010001001001;
		Coeff[1661] <= 15'b001010001001100;
		Coeff[1662] <= 15'b001010001001111;
		Coeff[1663] <= 15'b001010001010010;
		Coeff[1664] <= 15'b001010001010101;
		Coeff[1665] <= 15'b001010001011001;
		Coeff[1666] <= 15'b001010001011100;
		Coeff[1667] <= 15'b001010001011111;
		Coeff[1668] <= 15'b001010001100010;
		Coeff[1669] <= 15'b001010001100101;
		Coeff[1670] <= 15'b001010001101000;
		Coeff[1671] <= 15'b001010001101011;
		Coeff[1672] <= 15'b001010001101110;
		Coeff[1673] <= 15'b001010001110001;
		Coeff[1674] <= 15'b001010001110100;
		Coeff[1675] <= 15'b001010001111000;
		Coeff[1676] <= 15'b001010001111011;
		Coeff[1677] <= 15'b001010001111110;
		Coeff[1678] <= 15'b001010010000001;
		Coeff[1679] <= 15'b001010010000100;
		Coeff[1680] <= 15'b001010010000111;
		Coeff[1681] <= 15'b001010010001010;
		Coeff[1682] <= 15'b001010010001101;
		Coeff[1683] <= 15'b001010010010000;
		Coeff[1684] <= 15'b001010010010011;
		Coeff[1685] <= 15'b001010010010111;
		Coeff[1686] <= 15'b001010010011010;
		Coeff[1687] <= 15'b001010010011101;
		Coeff[1688] <= 15'b001010010100000;
		Coeff[1689] <= 15'b001010010100011;
		Coeff[1690] <= 15'b001010010100110;
		Coeff[1691] <= 15'b001010010101001;
		Coeff[1692] <= 15'b001010010101100;
		Coeff[1693] <= 15'b001010010101111;
		Coeff[1694] <= 15'b001010010110010;
		Coeff[1695] <= 15'b001010010110110;
		Coeff[1696] <= 15'b001010010111001;
		Coeff[1697] <= 15'b001010010111100;
		Coeff[1698] <= 15'b001010010111111;
		Coeff[1699] <= 15'b001010011000010;
		Coeff[1700] <= 15'b001010011000101;
		Coeff[1701] <= 15'b001010011001000;
		Coeff[1702] <= 15'b001010011001011;
		Coeff[1703] <= 15'b001010011001110;
		Coeff[1704] <= 15'b001010011010001;
		Coeff[1705] <= 15'b001010011010101;
		Coeff[1706] <= 15'b001010011011000;
		Coeff[1707] <= 15'b001010011011011;
		Coeff[1708] <= 15'b001010011011110;
		Coeff[1709] <= 15'b001010011100001;
		Coeff[1710] <= 15'b001010011100100;
		Coeff[1711] <= 15'b001010011100111;
		Coeff[1712] <= 15'b001010011101010;
		Coeff[1713] <= 15'b001010011101101;
		Coeff[1714] <= 15'b001010011110000;
		Coeff[1715] <= 15'b001010011110100;
		Coeff[1716] <= 15'b001010011110111;
		Coeff[1717] <= 15'b001010011111010;
		Coeff[1718] <= 15'b001010011111101;
		Coeff[1719] <= 15'b001010100000000;
		Coeff[1720] <= 15'b001010100000011;
		Coeff[1721] <= 15'b001010100000110;
		Coeff[1722] <= 15'b001010100001001;
		Coeff[1723] <= 15'b001010100001100;
		Coeff[1724] <= 15'b001010100001111;
		Coeff[1725] <= 15'b001010100010011;
		Coeff[1726] <= 15'b001010100010110;
		Coeff[1727] <= 15'b001010100011001;
		Coeff[1728] <= 15'b001010100011100;
		Coeff[1729] <= 15'b001010100011111;
		Coeff[1730] <= 15'b001010100100010;
		Coeff[1731] <= 15'b001010100100101;
		Coeff[1732] <= 15'b001010100101000;
		Coeff[1733] <= 15'b001010100101011;
		Coeff[1734] <= 15'b001010100101110;
		Coeff[1735] <= 15'b001010100110010;
		Coeff[1736] <= 15'b001010100110101;
		Coeff[1737] <= 15'b001010100111000;
		Coeff[1738] <= 15'b001010100111011;
		Coeff[1739] <= 15'b001010100111110;
		Coeff[1740] <= 15'b001010101000001;
		Coeff[1741] <= 15'b001010101000100;
		Coeff[1742] <= 15'b001010101000111;
		Coeff[1743] <= 15'b001010101001010;
		Coeff[1744] <= 15'b001010101001101;
		Coeff[1745] <= 15'b001010101010001;
		Coeff[1746] <= 15'b001010101010100;
		Coeff[1747] <= 15'b001010101010111;
		Coeff[1748] <= 15'b001010101011010;
		Coeff[1749] <= 15'b001010101011101;
		Coeff[1750] <= 15'b001010101100000;
		Coeff[1751] <= 15'b001010101100011;
		Coeff[1752] <= 15'b001010101100110;
		Coeff[1753] <= 15'b001010101101001;
		Coeff[1754] <= 15'b001010101101100;
		Coeff[1755] <= 15'b001010101110000;
		Coeff[1756] <= 15'b001010101110011;
		Coeff[1757] <= 15'b001010101110110;
		Coeff[1758] <= 15'b001010101111001;
		Coeff[1759] <= 15'b001010101111100;
		Coeff[1760] <= 15'b001010101111111;
		Coeff[1761] <= 15'b001010110000010;
		Coeff[1762] <= 15'b001010110000101;
		Coeff[1763] <= 15'b001010110001000;
		Coeff[1764] <= 15'b001010110001011;
		Coeff[1765] <= 15'b001010110001110;
		Coeff[1766] <= 15'b001010110010010;
		Coeff[1767] <= 15'b001010110010101;
		Coeff[1768] <= 15'b001010110011000;
		Coeff[1769] <= 15'b001010110011011;
		Coeff[1770] <= 15'b001010110011110;
		Coeff[1771] <= 15'b001010110100001;
		Coeff[1772] <= 15'b001010110100100;
		Coeff[1773] <= 15'b001010110100111;
		Coeff[1774] <= 15'b001010110101010;
		Coeff[1775] <= 15'b001010110101101;
		Coeff[1776] <= 15'b001010110110001;
		Coeff[1777] <= 15'b001010110110100;
		Coeff[1778] <= 15'b001010110110111;
		Coeff[1779] <= 15'b001010110111010;
		Coeff[1780] <= 15'b001010110111101;
		Coeff[1781] <= 15'b001010111000000;
		Coeff[1782] <= 15'b001010111000011;
		Coeff[1783] <= 15'b001010111000110;
		Coeff[1784] <= 15'b001010111001001;
		Coeff[1785] <= 15'b001010111001100;
		Coeff[1786] <= 15'b001010111010000;
		Coeff[1787] <= 15'b001010111010011;
		Coeff[1788] <= 15'b001010111010110;
		Coeff[1789] <= 15'b001010111011001;
		Coeff[1790] <= 15'b001010111011100;
		Coeff[1791] <= 15'b001010111011111;
		Coeff[1792] <= 15'b001010111100010;
		Coeff[1793] <= 15'b001010111100101;
		Coeff[1794] <= 15'b001010111101000;
		Coeff[1795] <= 15'b001010111101011;
		Coeff[1796] <= 15'b001010111101110;
		Coeff[1797] <= 15'b001010111110010;
		Coeff[1798] <= 15'b001010111110101;
		Coeff[1799] <= 15'b001010111111000;
		Coeff[1800] <= 15'b001010111111011;
		Coeff[1801] <= 15'b001010111111110;
		Coeff[1802] <= 15'b001011000000001;
		Coeff[1803] <= 15'b001011000000100;
		Coeff[1804] <= 15'b001011000000111;
		Coeff[1805] <= 15'b001011000001010;
		Coeff[1806] <= 15'b001011000001101;
		Coeff[1807] <= 15'b001011000010001;
		Coeff[1808] <= 15'b001011000010100;
		Coeff[1809] <= 15'b001011000010111;
		Coeff[1810] <= 15'b001011000011010;
		Coeff[1811] <= 15'b001011000011101;
		Coeff[1812] <= 15'b001011000100000;
		Coeff[1813] <= 15'b001011000100011;
		Coeff[1814] <= 15'b001011000100110;
		Coeff[1815] <= 15'b001011000101001;
		Coeff[1816] <= 15'b001011000101100;
		Coeff[1817] <= 15'b001011000101111;
		Coeff[1818] <= 15'b001011000110011;
		Coeff[1819] <= 15'b001011000110110;
		Coeff[1820] <= 15'b001011000111001;
		Coeff[1821] <= 15'b001011000111100;
		Coeff[1822] <= 15'b001011000111111;
		Coeff[1823] <= 15'b001011001000010;
		Coeff[1824] <= 15'b001011001000101;
		Coeff[1825] <= 15'b001011001001000;
		Coeff[1826] <= 15'b001011001001011;
		Coeff[1827] <= 15'b001011001001110;
		Coeff[1828] <= 15'b001011001010001;
		Coeff[1829] <= 15'b001011001010101;
		Coeff[1830] <= 15'b001011001011000;
		Coeff[1831] <= 15'b001011001011011;
		Coeff[1832] <= 15'b001011001011110;
		Coeff[1833] <= 15'b001011001100001;
		Coeff[1834] <= 15'b001011001100100;
		Coeff[1835] <= 15'b001011001100111;
		Coeff[1836] <= 15'b001011001101010;
		Coeff[1837] <= 15'b001011001101101;
		Coeff[1838] <= 15'b001011001110000;
		Coeff[1839] <= 15'b001011001110100;
		Coeff[1840] <= 15'b001011001110111;
		Coeff[1841] <= 15'b001011001111010;
		Coeff[1842] <= 15'b001011001111101;
		Coeff[1843] <= 15'b001011010000000;
		Coeff[1844] <= 15'b001011010000011;
		Coeff[1845] <= 15'b001011010000110;
		Coeff[1846] <= 15'b001011010001001;
		Coeff[1847] <= 15'b001011010001100;
		Coeff[1848] <= 15'b001011010001111;
		Coeff[1849] <= 15'b001011010010010;
		Coeff[1850] <= 15'b001011010010110;
		Coeff[1851] <= 15'b001011010011001;
		Coeff[1852] <= 15'b001011010011100;
		Coeff[1853] <= 15'b001011010011111;
		Coeff[1854] <= 15'b001011010100010;
		Coeff[1855] <= 15'b001011010100101;
		Coeff[1856] <= 15'b001011010101000;
		Coeff[1857] <= 15'b001011010101011;
		Coeff[1858] <= 15'b001011010101110;
		Coeff[1859] <= 15'b001011010110001;
		Coeff[1860] <= 15'b001011010110100;
		Coeff[1861] <= 15'b001011010111000;
		Coeff[1862] <= 15'b001011010111011;
		Coeff[1863] <= 15'b001011010111110;
		Coeff[1864] <= 15'b001011011000001;
		Coeff[1865] <= 15'b001011011000100;
		Coeff[1866] <= 15'b001011011000111;
		Coeff[1867] <= 15'b001011011001010;
		Coeff[1868] <= 15'b001011011001101;
		Coeff[1869] <= 15'b001011011010000;
		Coeff[1870] <= 15'b001011011010011;
		Coeff[1871] <= 15'b001011011010110;
		Coeff[1872] <= 15'b001011011011010;
		Coeff[1873] <= 15'b001011011011101;
		Coeff[1874] <= 15'b001011011100000;
		Coeff[1875] <= 15'b001011011100011;
		Coeff[1876] <= 15'b001011011100110;
		Coeff[1877] <= 15'b001011011101001;
		Coeff[1878] <= 15'b001011011101100;
		Coeff[1879] <= 15'b001011011101111;
		Coeff[1880] <= 15'b001011011110010;
		Coeff[1881] <= 15'b001011011110101;
		Coeff[1882] <= 15'b001011011111000;
		Coeff[1883] <= 15'b001011011111100;
		Coeff[1884] <= 15'b001011011111111;
		Coeff[1885] <= 15'b001011100000010;
		Coeff[1886] <= 15'b001011100000101;
		Coeff[1887] <= 15'b001011100001000;
		Coeff[1888] <= 15'b001011100001011;
		Coeff[1889] <= 15'b001011100001110;
		Coeff[1890] <= 15'b001011100010001;
		Coeff[1891] <= 15'b001011100010100;
		Coeff[1892] <= 15'b001011100010111;
		Coeff[1893] <= 15'b001011100011010;
		Coeff[1894] <= 15'b001011100011110;
		Coeff[1895] <= 15'b001011100100001;
		Coeff[1896] <= 15'b001011100100100;
		Coeff[1897] <= 15'b001011100100111;
		Coeff[1898] <= 15'b001011100101010;
		Coeff[1899] <= 15'b001011100101101;
		Coeff[1900] <= 15'b001011100110000;
		Coeff[1901] <= 15'b001011100110011;
		Coeff[1902] <= 15'b001011100110110;
		Coeff[1903] <= 15'b001011100111001;
		Coeff[1904] <= 15'b001011100111100;
		Coeff[1905] <= 15'b001011101000000;
		Coeff[1906] <= 15'b001011101000011;
		Coeff[1907] <= 15'b001011101000110;
		Coeff[1908] <= 15'b001011101001001;
		Coeff[1909] <= 15'b001011101001100;
		Coeff[1910] <= 15'b001011101001111;
		Coeff[1911] <= 15'b001011101010010;
		Coeff[1912] <= 15'b001011101010101;
		Coeff[1913] <= 15'b001011101011000;
		Coeff[1914] <= 15'b001011101011011;
		Coeff[1915] <= 15'b001011101011110;
		Coeff[1916] <= 15'b001011101100001;
		Coeff[1917] <= 15'b001011101100101;
		Coeff[1918] <= 15'b001011101101000;
		Coeff[1919] <= 15'b001011101101011;
		Coeff[1920] <= 15'b001011101101110;
		Coeff[1921] <= 15'b001011101110001;
		Coeff[1922] <= 15'b001011101110100;
		Coeff[1923] <= 15'b001011101110111;
		Coeff[1924] <= 15'b001011101111010;
		Coeff[1925] <= 15'b001011101111101;
		Coeff[1926] <= 15'b001011110000000;
		Coeff[1927] <= 15'b001011110000011;
		Coeff[1928] <= 15'b001011110000111;
		Coeff[1929] <= 15'b001011110001010;
		Coeff[1930] <= 15'b001011110001101;
		Coeff[1931] <= 15'b001011110010000;
		Coeff[1932] <= 15'b001011110010011;
		Coeff[1933] <= 15'b001011110010110;
		Coeff[1934] <= 15'b001011110011001;
		Coeff[1935] <= 15'b001011110011100;
		Coeff[1936] <= 15'b001011110011111;
		Coeff[1937] <= 15'b001011110100010;
		Coeff[1938] <= 15'b001011110100101;
		Coeff[1939] <= 15'b001011110101001;
		Coeff[1940] <= 15'b001011110101100;
		Coeff[1941] <= 15'b001011110101111;
		Coeff[1942] <= 15'b001011110110010;
		Coeff[1943] <= 15'b001011110110101;
		Coeff[1944] <= 15'b001011110111000;
		Coeff[1945] <= 15'b001011110111011;
		Coeff[1946] <= 15'b001011110111110;
		Coeff[1947] <= 15'b001011111000001;
		Coeff[1948] <= 15'b001011111000100;
		Coeff[1949] <= 15'b001011111000111;
		Coeff[1950] <= 15'b001011111001010;
		Coeff[1951] <= 15'b001011111001110;
		Coeff[1952] <= 15'b001011111010001;
		Coeff[1953] <= 15'b001011111010100;
		Coeff[1954] <= 15'b001011111010111;
		Coeff[1955] <= 15'b001011111011010;
		Coeff[1956] <= 15'b001011111011101;
		Coeff[1957] <= 15'b001011111100000;
		Coeff[1958] <= 15'b001011111100011;
		Coeff[1959] <= 15'b001011111100110;
		Coeff[1960] <= 15'b001011111101001;
		Coeff[1961] <= 15'b001011111101100;
		Coeff[1962] <= 15'b001011111110000;
		Coeff[1963] <= 15'b001011111110011;
		Coeff[1964] <= 15'b001011111110110;
		Coeff[1965] <= 15'b001011111111001;
		Coeff[1966] <= 15'b001011111111100;
		Coeff[1967] <= 15'b001011111111111;
		Coeff[1968] <= 15'b001100000000010;
		Coeff[1969] <= 15'b001100000000101;
		Coeff[1970] <= 15'b001100000001000;
		Coeff[1971] <= 15'b001100000001011;
		Coeff[1972] <= 15'b001100000001110;
		Coeff[1973] <= 15'b001100000010001;
		Coeff[1974] <= 15'b001100000010101;
		Coeff[1975] <= 15'b001100000011000;
		Coeff[1976] <= 15'b001100000011011;
		Coeff[1977] <= 15'b001100000011110;
		Coeff[1978] <= 15'b001100000100001;
		Coeff[1979] <= 15'b001100000100100;
		Coeff[1980] <= 15'b001100000100111;
		Coeff[1981] <= 15'b001100000101010;
		Coeff[1982] <= 15'b001100000101101;
		Coeff[1983] <= 15'b001100000110000;
		Coeff[1984] <= 15'b001100000110011;
		Coeff[1985] <= 15'b001100000110110;
		Coeff[1986] <= 15'b001100000111010;
		Coeff[1987] <= 15'b001100000111101;
		Coeff[1988] <= 15'b001100001000000;
		Coeff[1989] <= 15'b001100001000011;
		Coeff[1990] <= 15'b001100001000110;
		Coeff[1991] <= 15'b001100001001001;
		Coeff[1992] <= 15'b001100001001100;
		Coeff[1993] <= 15'b001100001001111;
		Coeff[1994] <= 15'b001100001010010;
		Coeff[1995] <= 15'b001100001010101;
		Coeff[1996] <= 15'b001100001011000;
		Coeff[1997] <= 15'b001100001011100;
		Coeff[1998] <= 15'b001100001011111;
		Coeff[1999] <= 15'b001100001100010;
		Coeff[2000] <= 15'b001100001100101;
		Coeff[2001] <= 15'b001100001101000;
		Coeff[2002] <= 15'b001100001101011;
		Coeff[2003] <= 15'b001100001101110;
		Coeff[2004] <= 15'b001100001110001;
		Coeff[2005] <= 15'b001100001110100;
		Coeff[2006] <= 15'b001100001110111;
		Coeff[2007] <= 15'b001100001111010;
		Coeff[2008] <= 15'b001100001111101;
		Coeff[2009] <= 15'b001100010000001;
		Coeff[2010] <= 15'b001100010000100;
		Coeff[2011] <= 15'b001100010000111;
		Coeff[2012] <= 15'b001100010001010;
		Coeff[2013] <= 15'b001100010001101;
		Coeff[2014] <= 15'b001100010010000;
		Coeff[2015] <= 15'b001100010010011;
		Coeff[2016] <= 15'b001100010010110;
		Coeff[2017] <= 15'b001100010011001;
		Coeff[2018] <= 15'b001100010011100;
		Coeff[2019] <= 15'b001100010011111;
		Coeff[2020] <= 15'b001100010100010;
		Coeff[2021] <= 15'b001100010100110;
		Coeff[2022] <= 15'b001100010101001;
		Coeff[2023] <= 15'b001100010101100;
		Coeff[2024] <= 15'b001100010101111;
		Coeff[2025] <= 15'b001100010110010;
		Coeff[2026] <= 15'b001100010110101;
		Coeff[2027] <= 15'b001100010111000;
		Coeff[2028] <= 15'b001100010111011;
		Coeff[2029] <= 15'b001100010111110;
		Coeff[2030] <= 15'b001100011000001;
		Coeff[2031] <= 15'b001100011000100;
		Coeff[2032] <= 15'b001100011000111;
		Coeff[2033] <= 15'b001100011001010;
		Coeff[2034] <= 15'b001100011001110;
		Coeff[2035] <= 15'b001100011010001;
		Coeff[2036] <= 15'b001100011010100;
		Coeff[2037] <= 15'b001100011010111;
		Coeff[2038] <= 15'b001100011011010;
		Coeff[2039] <= 15'b001100011011101;
		Coeff[2040] <= 15'b001100011100000;
		Coeff[2041] <= 15'b001100011100011;
		Coeff[2042] <= 15'b001100011100110;
		Coeff[2043] <= 15'b001100011101001;
		Coeff[2044] <= 15'b001100011101100;
		Coeff[2045] <= 15'b001100011101111;
		Coeff[2046] <= 15'b001100011110011;
		Coeff[2047] <= 15'b001100011110110;
		Coeff[2048] <= 15'b001100011111001;
		Coeff[2049] <= 15'b001100011111100;
		Coeff[2050] <= 15'b001100011111111;
		Coeff[2051] <= 15'b001100100000010;
		Coeff[2052] <= 15'b001100100000101;
		Coeff[2053] <= 15'b001100100001000;
		Coeff[2054] <= 15'b001100100001011;
		Coeff[2055] <= 15'b001100100001110;
		Coeff[2056] <= 15'b001100100010001;
		Coeff[2057] <= 15'b001100100010100;
		Coeff[2058] <= 15'b001100100011000;
		Coeff[2059] <= 15'b001100100011011;
		Coeff[2060] <= 15'b001100100011110;
		Coeff[2061] <= 15'b001100100100001;
		Coeff[2062] <= 15'b001100100100100;
		Coeff[2063] <= 15'b001100100100111;
		Coeff[2064] <= 15'b001100100101010;
		Coeff[2065] <= 15'b001100100101101;
		Coeff[2066] <= 15'b001100100110000;
		Coeff[2067] <= 15'b001100100110011;
		Coeff[2068] <= 15'b001100100110110;
		Coeff[2069] <= 15'b001100100111001;
		Coeff[2070] <= 15'b001100100111100;
		Coeff[2071] <= 15'b001100101000000;
		Coeff[2072] <= 15'b001100101000011;
		Coeff[2073] <= 15'b001100101000110;
		Coeff[2074] <= 15'b001100101001001;
		Coeff[2075] <= 15'b001100101001100;
		Coeff[2076] <= 15'b001100101001111;
		Coeff[2077] <= 15'b001100101010010;
		Coeff[2078] <= 15'b001100101010101;
		Coeff[2079] <= 15'b001100101011000;
		Coeff[2080] <= 15'b001100101011011;
		Coeff[2081] <= 15'b001100101011110;
		Coeff[2082] <= 15'b001100101100001;
		Coeff[2083] <= 15'b001100101100101;
		Coeff[2084] <= 15'b001100101101000;
		Coeff[2085] <= 15'b001100101101011;
		Coeff[2086] <= 15'b001100101101110;
		Coeff[2087] <= 15'b001100101110001;
		Coeff[2088] <= 15'b001100101110100;
		Coeff[2089] <= 15'b001100101110111;
		Coeff[2090] <= 15'b001100101111010;
		Coeff[2091] <= 15'b001100101111101;
		Coeff[2092] <= 15'b001100110000000;
		Coeff[2093] <= 15'b001100110000011;
		Coeff[2094] <= 15'b001100110000110;
		Coeff[2095] <= 15'b001100110001001;
		Coeff[2096] <= 15'b001100110001101;
		Coeff[2097] <= 15'b001100110010000;
		Coeff[2098] <= 15'b001100110010011;
		Coeff[2099] <= 15'b001100110010110;
		Coeff[2100] <= 15'b001100110011001;
		Coeff[2101] <= 15'b001100110011100;
		Coeff[2102] <= 15'b001100110011111;
		Coeff[2103] <= 15'b001100110100010;
		Coeff[2104] <= 15'b001100110100101;
		Coeff[2105] <= 15'b001100110101000;
		Coeff[2106] <= 15'b001100110101011;
		Coeff[2107] <= 15'b001100110101110;
		Coeff[2108] <= 15'b001100110110001;
		Coeff[2109] <= 15'b001100110110101;
		Coeff[2110] <= 15'b001100110111000;
		Coeff[2111] <= 15'b001100110111011;
		Coeff[2112] <= 15'b001100110111110;
		Coeff[2113] <= 15'b001100111000001;
		Coeff[2114] <= 15'b001100111000100;
		Coeff[2115] <= 15'b001100111000111;
		Coeff[2116] <= 15'b001100111001010;
		Coeff[2117] <= 15'b001100111001101;
		Coeff[2118] <= 15'b001100111010000;
		Coeff[2119] <= 15'b001100111010011;
		Coeff[2120] <= 15'b001100111010110;
		Coeff[2121] <= 15'b001100111011001;
		Coeff[2122] <= 15'b001100111011101;
		Coeff[2123] <= 15'b001100111100000;
		Coeff[2124] <= 15'b001100111100011;
		Coeff[2125] <= 15'b001100111100110;
		Coeff[2126] <= 15'b001100111101001;
		Coeff[2127] <= 15'b001100111101100;
		Coeff[2128] <= 15'b001100111101111;
		Coeff[2129] <= 15'b001100111110010;
		Coeff[2130] <= 15'b001100111110101;
		Coeff[2131] <= 15'b001100111111000;
		Coeff[2132] <= 15'b001100111111011;
		Coeff[2133] <= 15'b001100111111110;
		Coeff[2134] <= 15'b001101000000001;
		Coeff[2135] <= 15'b001101000000101;
		Coeff[2136] <= 15'b001101000001000;
		Coeff[2137] <= 15'b001101000001011;
		Coeff[2138] <= 15'b001101000001110;
		Coeff[2139] <= 15'b001101000010001;
		Coeff[2140] <= 15'b001101000010100;
		Coeff[2141] <= 15'b001101000010111;
		Coeff[2142] <= 15'b001101000011010;
		Coeff[2143] <= 15'b001101000011101;
		Coeff[2144] <= 15'b001101000100000;
		Coeff[2145] <= 15'b001101000100011;
		Coeff[2146] <= 15'b001101000100110;
		Coeff[2147] <= 15'b001101000101001;
		Coeff[2148] <= 15'b001101000101101;
		Coeff[2149] <= 15'b001101000110000;
		Coeff[2150] <= 15'b001101000110011;
		Coeff[2151] <= 15'b001101000110110;
		Coeff[2152] <= 15'b001101000111001;
		Coeff[2153] <= 15'b001101000111100;
		Coeff[2154] <= 15'b001101000111111;
		Coeff[2155] <= 15'b001101001000010;
		Coeff[2156] <= 15'b001101001000101;
		Coeff[2157] <= 15'b001101001001000;
		Coeff[2158] <= 15'b001101001001011;
		Coeff[2159] <= 15'b001101001001110;
		Coeff[2160] <= 15'b001101001010001;
		Coeff[2161] <= 15'b001101001010101;
		Coeff[2162] <= 15'b001101001011000;
		Coeff[2163] <= 15'b001101001011011;
		Coeff[2164] <= 15'b001101001011110;
		Coeff[2165] <= 15'b001101001100001;
		Coeff[2166] <= 15'b001101001100100;
		Coeff[2167] <= 15'b001101001100111;
		Coeff[2168] <= 15'b001101001101010;
		Coeff[2169] <= 15'b001101001101101;
		Coeff[2170] <= 15'b001101001110000;
		Coeff[2171] <= 15'b001101001110011;
		Coeff[2172] <= 15'b001101001110110;
		Coeff[2173] <= 15'b001101001111001;
		Coeff[2174] <= 15'b001101001111100;
		Coeff[2175] <= 15'b001101010000000;
		Coeff[2176] <= 15'b001101010000011;
		Coeff[2177] <= 15'b001101010000110;
		Coeff[2178] <= 15'b001101010001001;
		Coeff[2179] <= 15'b001101010001100;
		Coeff[2180] <= 15'b001101010001111;
		Coeff[2181] <= 15'b001101010010010;
		Coeff[2182] <= 15'b001101010010101;
		Coeff[2183] <= 15'b001101010011000;
		Coeff[2184] <= 15'b001101010011011;
		Coeff[2185] <= 15'b001101010011110;
		Coeff[2186] <= 15'b001101010100001;
		Coeff[2187] <= 15'b001101010100100;
		Coeff[2188] <= 15'b001101010101000;
		Coeff[2189] <= 15'b001101010101011;
		Coeff[2190] <= 15'b001101010101110;
		Coeff[2191] <= 15'b001101010110001;
		Coeff[2192] <= 15'b001101010110100;
		Coeff[2193] <= 15'b001101010110111;
		Coeff[2194] <= 15'b001101010111010;
		Coeff[2195] <= 15'b001101010111101;
		Coeff[2196] <= 15'b001101011000000;
		Coeff[2197] <= 15'b001101011000011;
		Coeff[2198] <= 15'b001101011000110;
		Coeff[2199] <= 15'b001101011001001;
		Coeff[2200] <= 15'b001101011001100;
		Coeff[2201] <= 15'b001101011001111;
		Coeff[2202] <= 15'b001101011010011;
		Coeff[2203] <= 15'b001101011010110;
		Coeff[2204] <= 15'b001101011011001;
		Coeff[2205] <= 15'b001101011011100;
		Coeff[2206] <= 15'b001101011011111;
		Coeff[2207] <= 15'b001101011100010;
		Coeff[2208] <= 15'b001101011100101;
		Coeff[2209] <= 15'b001101011101000;
		Coeff[2210] <= 15'b001101011101011;
		Coeff[2211] <= 15'b001101011101110;
		Coeff[2212] <= 15'b001101011110001;
		Coeff[2213] <= 15'b001101011110100;
		Coeff[2214] <= 15'b001101011110111;
		Coeff[2215] <= 15'b001101011111010;
		Coeff[2216] <= 15'b001101011111110;
		Coeff[2217] <= 15'b001101100000001;
		Coeff[2218] <= 15'b001101100000100;
		Coeff[2219] <= 15'b001101100000111;
		Coeff[2220] <= 15'b001101100001010;
		Coeff[2221] <= 15'b001101100001101;
		Coeff[2222] <= 15'b001101100010000;
		Coeff[2223] <= 15'b001101100010011;
		Coeff[2224] <= 15'b001101100010110;
		Coeff[2225] <= 15'b001101100011001;
		Coeff[2226] <= 15'b001101100011100;
		Coeff[2227] <= 15'b001101100011111;
		Coeff[2228] <= 15'b001101100100010;
		Coeff[2229] <= 15'b001101100100101;
		Coeff[2230] <= 15'b001101100101001;
		Coeff[2231] <= 15'b001101100101100;
		Coeff[2232] <= 15'b001101100101111;
		Coeff[2233] <= 15'b001101100110010;
		Coeff[2234] <= 15'b001101100110101;
		Coeff[2235] <= 15'b001101100111000;
		Coeff[2236] <= 15'b001101100111011;
		Coeff[2237] <= 15'b001101100111110;
		Coeff[2238] <= 15'b001101101000001;
		Coeff[2239] <= 15'b001101101000100;
		Coeff[2240] <= 15'b001101101000111;
		Coeff[2241] <= 15'b001101101001010;
		Coeff[2242] <= 15'b001101101001101;
		Coeff[2243] <= 15'b001101101010000;
		Coeff[2244] <= 15'b001101101010011;
		Coeff[2245] <= 15'b001101101010111;
		Coeff[2246] <= 15'b001101101011010;
		Coeff[2247] <= 15'b001101101011101;
		Coeff[2248] <= 15'b001101101100000;
		Coeff[2249] <= 15'b001101101100011;
		Coeff[2250] <= 15'b001101101100110;
		Coeff[2251] <= 15'b001101101101001;
		Coeff[2252] <= 15'b001101101101100;
		Coeff[2253] <= 15'b001101101101111;
		Coeff[2254] <= 15'b001101101110010;
		Coeff[2255] <= 15'b001101101110101;
		Coeff[2256] <= 15'b001101101111000;
		Coeff[2257] <= 15'b001101101111011;
		Coeff[2258] <= 15'b001101101111110;
		Coeff[2259] <= 15'b001101110000010;
		Coeff[2260] <= 15'b001101110000101;
		Coeff[2261] <= 15'b001101110001000;
		Coeff[2262] <= 15'b001101110001011;
		Coeff[2263] <= 15'b001101110001110;
		Coeff[2264] <= 15'b001101110010001;
		Coeff[2265] <= 15'b001101110010100;
		Coeff[2266] <= 15'b001101110010111;
		Coeff[2267] <= 15'b001101110011010;
		Coeff[2268] <= 15'b001101110011101;
		Coeff[2269] <= 15'b001101110100000;
		Coeff[2270] <= 15'b001101110100011;
		Coeff[2271] <= 15'b001101110100110;
		Coeff[2272] <= 15'b001101110101001;
		Coeff[2273] <= 15'b001101110101100;
		Coeff[2274] <= 15'b001101110110000;
		Coeff[2275] <= 15'b001101110110011;
		Coeff[2276] <= 15'b001101110110110;
		Coeff[2277] <= 15'b001101110111001;
		Coeff[2278] <= 15'b001101110111100;
		Coeff[2279] <= 15'b001101110111111;
		Coeff[2280] <= 15'b001101111000010;
		Coeff[2281] <= 15'b001101111000101;
		Coeff[2282] <= 15'b001101111001000;
		Coeff[2283] <= 15'b001101111001011;
		Coeff[2284] <= 15'b001101111001110;
		Coeff[2285] <= 15'b001101111010001;
		Coeff[2286] <= 15'b001101111010100;
		Coeff[2287] <= 15'b001101111010111;
		Coeff[2288] <= 15'b001101111011010;
		Coeff[2289] <= 15'b001101111011110;
		Coeff[2290] <= 15'b001101111100001;
		Coeff[2291] <= 15'b001101111100100;
		Coeff[2292] <= 15'b001101111100111;
		Coeff[2293] <= 15'b001101111101010;
		Coeff[2294] <= 15'b001101111101101;
		Coeff[2295] <= 15'b001101111110000;
		Coeff[2296] <= 15'b001101111110011;
		Coeff[2297] <= 15'b001101111110110;
		Coeff[2298] <= 15'b001101111111001;
		Coeff[2299] <= 15'b001101111111100;
		Coeff[2300] <= 15'b001101111111111;
		Coeff[2301] <= 15'b001110000000010;
		Coeff[2302] <= 15'b001110000000101;
		Coeff[2303] <= 15'b001110000001000;
		Coeff[2304] <= 15'b001110000001100;
		Coeff[2305] <= 15'b001110000001111;
		Coeff[2306] <= 15'b001110000010010;
		Coeff[2307] <= 15'b001110000010101;
		Coeff[2308] <= 15'b001110000011000;
		Coeff[2309] <= 15'b001110000011011;
		Coeff[2310] <= 15'b001110000011110;
		Coeff[2311] <= 15'b001110000100001;
		Coeff[2312] <= 15'b001110000100100;
		Coeff[2313] <= 15'b001110000100111;
		Coeff[2314] <= 15'b001110000101010;
		Coeff[2315] <= 15'b001110000101101;
		Coeff[2316] <= 15'b001110000110000;
		Coeff[2317] <= 15'b001110000110011;
		Coeff[2318] <= 15'b001110000110110;
		Coeff[2319] <= 15'b001110000111001;
		Coeff[2320] <= 15'b001110000111101;
		Coeff[2321] <= 15'b001110001000000;
		Coeff[2322] <= 15'b001110001000011;
		Coeff[2323] <= 15'b001110001000110;
		Coeff[2324] <= 15'b001110001001001;
		Coeff[2325] <= 15'b001110001001100;
		Coeff[2326] <= 15'b001110001001111;
		Coeff[2327] <= 15'b001110001010010;
		Coeff[2328] <= 15'b001110001010101;
		Coeff[2329] <= 15'b001110001011000;
		Coeff[2330] <= 15'b001110001011011;
		Coeff[2331] <= 15'b001110001011110;
		Coeff[2332] <= 15'b001110001100001;
		Coeff[2333] <= 15'b001110001100100;
		Coeff[2334] <= 15'b001110001100111;
		Coeff[2335] <= 15'b001110001101011;
		Coeff[2336] <= 15'b001110001101110;
		Coeff[2337] <= 15'b001110001110001;
		Coeff[2338] <= 15'b001110001110100;
		Coeff[2339] <= 15'b001110001110111;
		Coeff[2340] <= 15'b001110001111010;
		Coeff[2341] <= 15'b001110001111101;
		Coeff[2342] <= 15'b001110010000000;
		Coeff[2343] <= 15'b001110010000011;
		Coeff[2344] <= 15'b001110010000110;
		Coeff[2345] <= 15'b001110010001001;
		Coeff[2346] <= 15'b001110010001100;
		Coeff[2347] <= 15'b001110010001111;
		Coeff[2348] <= 15'b001110010010010;
		Coeff[2349] <= 15'b001110010010101;
		Coeff[2350] <= 15'b001110010011000;
		Coeff[2351] <= 15'b001110010011100;
		Coeff[2352] <= 15'b001110010011111;
		Coeff[2353] <= 15'b001110010100010;
		Coeff[2354] <= 15'b001110010100101;
		Coeff[2355] <= 15'b001110010101000;
		Coeff[2356] <= 15'b001110010101011;
		Coeff[2357] <= 15'b001110010101110;
		Coeff[2358] <= 15'b001110010110001;
		Coeff[2359] <= 15'b001110010110100;
		Coeff[2360] <= 15'b001110010110111;
		Coeff[2361] <= 15'b001110010111010;
		Coeff[2362] <= 15'b001110010111101;
		Coeff[2363] <= 15'b001110011000000;
		Coeff[2364] <= 15'b001110011000011;
		Coeff[2365] <= 15'b001110011000110;
		Coeff[2366] <= 15'b001110011001001;
		Coeff[2367] <= 15'b001110011001100;
		Coeff[2368] <= 15'b001110011010000;
		Coeff[2369] <= 15'b001110011010011;
		Coeff[2370] <= 15'b001110011010110;
		Coeff[2371] <= 15'b001110011011001;
		Coeff[2372] <= 15'b001110011011100;
		Coeff[2373] <= 15'b001110011011111;
		Coeff[2374] <= 15'b001110011100010;
		Coeff[2375] <= 15'b001110011100101;
		Coeff[2376] <= 15'b001110011101000;
		Coeff[2377] <= 15'b001110011101011;
		Coeff[2378] <= 15'b001110011101110;
		Coeff[2379] <= 15'b001110011110001;
		Coeff[2380] <= 15'b001110011110100;
		Coeff[2381] <= 15'b001110011110111;
		Coeff[2382] <= 15'b001110011111010;
		Coeff[2383] <= 15'b001110011111101;
		Coeff[2384] <= 15'b001110100000001;
		Coeff[2385] <= 15'b001110100000100;
		Coeff[2386] <= 15'b001110100000111;
		Coeff[2387] <= 15'b001110100001010;
		Coeff[2388] <= 15'b001110100001101;
		Coeff[2389] <= 15'b001110100010000;
		Coeff[2390] <= 15'b001110100010011;
		Coeff[2391] <= 15'b001110100010110;
		Coeff[2392] <= 15'b001110100011001;
		Coeff[2393] <= 15'b001110100011100;
		Coeff[2394] <= 15'b001110100011111;
		Coeff[2395] <= 15'b001110100100010;
		Coeff[2396] <= 15'b001110100100101;
		Coeff[2397] <= 15'b001110100101000;
		Coeff[2398] <= 15'b001110100101011;
		Coeff[2399] <= 15'b001110100101110;
		Coeff[2400] <= 15'b001110100110001;
		Coeff[2401] <= 15'b001110100110101;
		Coeff[2402] <= 15'b001110100111000;
		Coeff[2403] <= 15'b001110100111011;
		Coeff[2404] <= 15'b001110100111110;
		Coeff[2405] <= 15'b001110101000001;
		Coeff[2406] <= 15'b001110101000100;
		Coeff[2407] <= 15'b001110101000111;
		Coeff[2408] <= 15'b001110101001010;
		Coeff[2409] <= 15'b001110101001101;
		Coeff[2410] <= 15'b001110101010000;
		Coeff[2411] <= 15'b001110101010011;
		Coeff[2412] <= 15'b001110101010110;
		Coeff[2413] <= 15'b001110101011001;
		Coeff[2414] <= 15'b001110101011100;
		Coeff[2415] <= 15'b001110101011111;
		Coeff[2416] <= 15'b001110101100010;
		Coeff[2417] <= 15'b001110101100101;
		Coeff[2418] <= 15'b001110101101001;
		Coeff[2419] <= 15'b001110101101100;
		Coeff[2420] <= 15'b001110101101111;
		Coeff[2421] <= 15'b001110101110010;
		Coeff[2422] <= 15'b001110101110101;
		Coeff[2423] <= 15'b001110101111000;
		Coeff[2424] <= 15'b001110101111011;
		Coeff[2425] <= 15'b001110101111110;
		Coeff[2426] <= 15'b001110110000001;
		Coeff[2427] <= 15'b001110110000100;
		Coeff[2428] <= 15'b001110110000111;
		Coeff[2429] <= 15'b001110110001010;
		Coeff[2430] <= 15'b001110110001101;
		Coeff[2431] <= 15'b001110110010000;
		Coeff[2432] <= 15'b001110110010011;
		Coeff[2433] <= 15'b001110110010110;
		Coeff[2434] <= 15'b001110110011001;
		Coeff[2435] <= 15'b001110110011100;
		Coeff[2436] <= 15'b001110110100000;
		Coeff[2437] <= 15'b001110110100011;
		Coeff[2438] <= 15'b001110110100110;
		Coeff[2439] <= 15'b001110110101001;
		Coeff[2440] <= 15'b001110110101100;
		Coeff[2441] <= 15'b001110110101111;
		Coeff[2442] <= 15'b001110110110010;
		Coeff[2443] <= 15'b001110110110101;
		Coeff[2444] <= 15'b001110110111000;
		Coeff[2445] <= 15'b001110110111011;
		Coeff[2446] <= 15'b001110110111110;
		Coeff[2447] <= 15'b001110111000001;
		Coeff[2448] <= 15'b001110111000100;
		Coeff[2449] <= 15'b001110111000111;
		Coeff[2450] <= 15'b001110111001010;
		Coeff[2451] <= 15'b001110111001101;
		Coeff[2452] <= 15'b001110111010000;
		Coeff[2453] <= 15'b001110111010011;
		Coeff[2454] <= 15'b001110111010111;
		Coeff[2455] <= 15'b001110111011010;
		Coeff[2456] <= 15'b001110111011101;
		Coeff[2457] <= 15'b001110111100000;
		Coeff[2458] <= 15'b001110111100011;
		Coeff[2459] <= 15'b001110111100110;
		Coeff[2460] <= 15'b001110111101001;
		Coeff[2461] <= 15'b001110111101100;
		Coeff[2462] <= 15'b001110111101111;
		Coeff[2463] <= 15'b001110111110010;
		Coeff[2464] <= 15'b001110111110101;
		Coeff[2465] <= 15'b001110111111000;
		Coeff[2466] <= 15'b001110111111011;
		Coeff[2467] <= 15'b001110111111110;
		Coeff[2468] <= 15'b001111000000001;
		Coeff[2469] <= 15'b001111000000100;
		Coeff[2470] <= 15'b001111000000111;
		Coeff[2471] <= 15'b001111000001010;
		Coeff[2472] <= 15'b001111000001110;
		Coeff[2473] <= 15'b001111000010001;
		Coeff[2474] <= 15'b001111000010100;
		Coeff[2475] <= 15'b001111000010111;
		Coeff[2476] <= 15'b001111000011010;
		Coeff[2477] <= 15'b001111000011101;
		Coeff[2478] <= 15'b001111000100000;
		Coeff[2479] <= 15'b001111000100011;
		Coeff[2480] <= 15'b001111000100110;
		Coeff[2481] <= 15'b001111000101001;
		Coeff[2482] <= 15'b001111000101100;
		Coeff[2483] <= 15'b001111000101111;
		Coeff[2484] <= 15'b001111000110010;
		Coeff[2485] <= 15'b001111000110101;
		Coeff[2486] <= 15'b001111000111000;
		Coeff[2487] <= 15'b001111000111011;
		Coeff[2488] <= 15'b001111000111110;
		Coeff[2489] <= 15'b001111001000001;
		Coeff[2490] <= 15'b001111001000100;
		Coeff[2491] <= 15'b001111001001000;
		Coeff[2492] <= 15'b001111001001011;
		Coeff[2493] <= 15'b001111001001110;
		Coeff[2494] <= 15'b001111001010001;
		Coeff[2495] <= 15'b001111001010100;
		Coeff[2496] <= 15'b001111001010111;
		Coeff[2497] <= 15'b001111001011010;
		Coeff[2498] <= 15'b001111001011101;
		Coeff[2499] <= 15'b001111001100000;
		Coeff[2500] <= 15'b001111001100011;
		Coeff[2501] <= 15'b001111001100110;
		Coeff[2502] <= 15'b001111001101001;
		Coeff[2503] <= 15'b001111001101100;
		Coeff[2504] <= 15'b001111001101111;
		Coeff[2505] <= 15'b001111001110010;
		Coeff[2506] <= 15'b001111001110101;
		Coeff[2507] <= 15'b001111001111000;
		Coeff[2508] <= 15'b001111001111011;
		Coeff[2509] <= 15'b001111001111110;
		Coeff[2510] <= 15'b001111010000010;
		Coeff[2511] <= 15'b001111010000101;
		Coeff[2512] <= 15'b001111010001000;
		Coeff[2513] <= 15'b001111010001011;
		Coeff[2514] <= 15'b001111010001110;
		Coeff[2515] <= 15'b001111010010001;
		Coeff[2516] <= 15'b001111010010100;
		Coeff[2517] <= 15'b001111010010111;
		Coeff[2518] <= 15'b001111010011010;
		Coeff[2519] <= 15'b001111010011101;
		Coeff[2520] <= 15'b001111010100000;
		Coeff[2521] <= 15'b001111010100011;
		Coeff[2522] <= 15'b001111010100110;
		Coeff[2523] <= 15'b001111010101001;
		Coeff[2524] <= 15'b001111010101100;
		Coeff[2525] <= 15'b001111010101111;
		Coeff[2526] <= 15'b001111010110010;
		Coeff[2527] <= 15'b001111010110101;
		Coeff[2528] <= 15'b001111010111000;
		Coeff[2529] <= 15'b001111010111011;
		Coeff[2530] <= 15'b001111010111111;
		Coeff[2531] <= 15'b001111011000010;
		Coeff[2532] <= 15'b001111011000101;
		Coeff[2533] <= 15'b001111011001000;
		Coeff[2534] <= 15'b001111011001011;
		Coeff[2535] <= 15'b001111011001110;
		Coeff[2536] <= 15'b001111011010001;
		Coeff[2537] <= 15'b001111011010100;
		Coeff[2538] <= 15'b001111011010111;
		Coeff[2539] <= 15'b001111011011010;
		Coeff[2540] <= 15'b001111011011101;
		Coeff[2541] <= 15'b001111011100000;
		Coeff[2542] <= 15'b001111011100011;
		Coeff[2543] <= 15'b001111011100110;
		Coeff[2544] <= 15'b001111011101001;
		Coeff[2545] <= 15'b001111011101100;
		Coeff[2546] <= 15'b001111011101111;
		Coeff[2547] <= 15'b001111011110010;
		Coeff[2548] <= 15'b001111011110101;
		Coeff[2549] <= 15'b001111011111000;
		Coeff[2550] <= 15'b001111011111011;
		Coeff[2551] <= 15'b001111011111111;
		Coeff[2552] <= 15'b001111100000010;
		Coeff[2553] <= 15'b001111100000101;
		Coeff[2554] <= 15'b001111100001000;
		Coeff[2555] <= 15'b001111100001011;
		Coeff[2556] <= 15'b001111100001110;
		Coeff[2557] <= 15'b001111100010001;
		Coeff[2558] <= 15'b001111100010100;
		Coeff[2559] <= 15'b001111100010111;
		Coeff[2560] <= 15'b001111100011010;
		Coeff[2561] <= 15'b001111100011101;
		Coeff[2562] <= 15'b001111100100000;
		Coeff[2563] <= 15'b001111100100011;
		Coeff[2564] <= 15'b001111100100110;
		Coeff[2565] <= 15'b001111100101001;
		Coeff[2566] <= 15'b001111100101100;
		Coeff[2567] <= 15'b001111100101111;
		Coeff[2568] <= 15'b001111100110010;
		Coeff[2569] <= 15'b001111100110101;
		Coeff[2570] <= 15'b001111100111000;
		Coeff[2571] <= 15'b001111100111011;
		Coeff[2572] <= 15'b001111100111111;
		Coeff[2573] <= 15'b001111101000010;
		Coeff[2574] <= 15'b001111101000101;
		Coeff[2575] <= 15'b001111101001000;
		Coeff[2576] <= 15'b001111101001011;
		Coeff[2577] <= 15'b001111101001110;
		Coeff[2578] <= 15'b001111101010001;
		Coeff[2579] <= 15'b001111101010100;
		Coeff[2580] <= 15'b001111101010111;
		Coeff[2581] <= 15'b001111101011010;
		Coeff[2582] <= 15'b001111101011101;
		Coeff[2583] <= 15'b001111101100000;
		Coeff[2584] <= 15'b001111101100011;
		Coeff[2585] <= 15'b001111101100110;
		Coeff[2586] <= 15'b001111101101001;
		Coeff[2587] <= 15'b001111101101100;
		Coeff[2588] <= 15'b001111101101111;
		Coeff[2589] <= 15'b001111101110010;
		Coeff[2590] <= 15'b001111101110101;
		Coeff[2591] <= 15'b001111101111000;
		Coeff[2592] <= 15'b001111101111011;
		Coeff[2593] <= 15'b001111101111111;
		Coeff[2594] <= 15'b001111110000010;
		Coeff[2595] <= 15'b001111110000101;
		Coeff[2596] <= 15'b001111110001000;
		Coeff[2597] <= 15'b001111110001011;
		Coeff[2598] <= 15'b001111110001110;
		Coeff[2599] <= 15'b001111110010001;
		Coeff[2600] <= 15'b001111110010100;
		Coeff[2601] <= 15'b001111110010111;
		Coeff[2602] <= 15'b001111110011010;
		Coeff[2603] <= 15'b001111110011101;
		Coeff[2604] <= 15'b001111110100000;
		Coeff[2605] <= 15'b001111110100011;
		Coeff[2606] <= 15'b001111110100110;
		Coeff[2607] <= 15'b001111110101001;
		Coeff[2608] <= 15'b001111110101100;
		Coeff[2609] <= 15'b001111110101111;
		Coeff[2610] <= 15'b001111110110010;
		Coeff[2611] <= 15'b001111110110101;
		Coeff[2612] <= 15'b001111110111000;
		Coeff[2613] <= 15'b001111110111011;
		Coeff[2614] <= 15'b001111110111110;
		Coeff[2615] <= 15'b001111111000001;
		Coeff[2616] <= 15'b001111111000101;
		Coeff[2617] <= 15'b001111111001000;
		Coeff[2618] <= 15'b001111111001011;
		Coeff[2619] <= 15'b001111111001110;
		Coeff[2620] <= 15'b001111111010001;
		Coeff[2621] <= 15'b001111111010100;
		Coeff[2622] <= 15'b001111111010111;
		Coeff[2623] <= 15'b001111111011010;
		Coeff[2624] <= 15'b001111111011101;
		Coeff[2625] <= 15'b001111111100000;
		Coeff[2626] <= 15'b001111111100011;
		Coeff[2627] <= 15'b001111111100110;
		Coeff[2628] <= 15'b001111111101001;
		Coeff[2629] <= 15'b001111111101100;
		Coeff[2630] <= 15'b001111111101111;
		Coeff[2631] <= 15'b001111111110010;
		Coeff[2632] <= 15'b001111111110101;
		Coeff[2633] <= 15'b001111111111000;
		Coeff[2634] <= 15'b001111111111011;
		Coeff[2635] <= 15'b001111111111110;
		Coeff[2636] <= 15'b010000000000001;
		Coeff[2637] <= 15'b010000000000100;
		Coeff[2638] <= 15'b010000000000111;
		Coeff[2639] <= 15'b010000000001010;
		Coeff[2640] <= 15'b010000000001110;
		Coeff[2641] <= 15'b010000000010001;
		Coeff[2642] <= 15'b010000000010100;
		Coeff[2643] <= 15'b010000000010111;
		Coeff[2644] <= 15'b010000000011010;
		Coeff[2645] <= 15'b010000000011101;
		Coeff[2646] <= 15'b010000000100000;
		Coeff[2647] <= 15'b010000000100011;
		Coeff[2648] <= 15'b010000000100110;
		Coeff[2649] <= 15'b010000000101001;
		Coeff[2650] <= 15'b010000000101100;
		Coeff[2651] <= 15'b010000000101111;
		Coeff[2652] <= 15'b010000000110010;
		Coeff[2653] <= 15'b010000000110101;
		Coeff[2654] <= 15'b010000000111000;
		Coeff[2655] <= 15'b010000000111011;
		Coeff[2656] <= 15'b010000000111110;
		Coeff[2657] <= 15'b010000001000001;
		Coeff[2658] <= 15'b010000001000100;
		Coeff[2659] <= 15'b010000001000111;
		Coeff[2660] <= 15'b010000001001010;
		Coeff[2661] <= 15'b010000001001101;
		Coeff[2662] <= 15'b010000001010000;
		Coeff[2663] <= 15'b010000001010011;
		Coeff[2664] <= 15'b010000001010111;
		Coeff[2665] <= 15'b010000001011010;
		Coeff[2666] <= 15'b010000001011101;
		Coeff[2667] <= 15'b010000001100000;
		Coeff[2668] <= 15'b010000001100011;
		Coeff[2669] <= 15'b010000001100110;
		Coeff[2670] <= 15'b010000001101001;
		Coeff[2671] <= 15'b010000001101100;
		Coeff[2672] <= 15'b010000001101111;
		Coeff[2673] <= 15'b010000001110010;
		Coeff[2674] <= 15'b010000001110101;
		Coeff[2675] <= 15'b010000001111000;
		Coeff[2676] <= 15'b010000001111011;
		Coeff[2677] <= 15'b010000001111110;
		Coeff[2678] <= 15'b010000010000001;
		Coeff[2679] <= 15'b010000010000100;
		Coeff[2680] <= 15'b010000010000111;
		Coeff[2681] <= 15'b010000010001010;
		Coeff[2682] <= 15'b010000010001101;
		Coeff[2683] <= 15'b010000010010000;
		Coeff[2684] <= 15'b010000010010011;
		Coeff[2685] <= 15'b010000010010110;
		Coeff[2686] <= 15'b010000010011001;
		Coeff[2687] <= 15'b010000010011100;
		Coeff[2688] <= 15'b010000010011111;
		Coeff[2689] <= 15'b010000010100010;
		Coeff[2690] <= 15'b010000010100110;
		Coeff[2691] <= 15'b010000010101001;
		Coeff[2692] <= 15'b010000010101100;
		Coeff[2693] <= 15'b010000010101111;
		Coeff[2694] <= 15'b010000010110010;
		Coeff[2695] <= 15'b010000010110101;
		Coeff[2696] <= 15'b010000010111000;
		Coeff[2697] <= 15'b010000010111011;
		Coeff[2698] <= 15'b010000010111110;
		Coeff[2699] <= 15'b010000011000001;
		Coeff[2700] <= 15'b010000011000100;
		Coeff[2701] <= 15'b010000011000111;
		Coeff[2702] <= 15'b010000011001010;
		Coeff[2703] <= 15'b010000011001101;
		Coeff[2704] <= 15'b010000011010000;
		Coeff[2705] <= 15'b010000011010011;
		Coeff[2706] <= 15'b010000011010110;
		Coeff[2707] <= 15'b010000011011001;
		Coeff[2708] <= 15'b010000011011100;
		Coeff[2709] <= 15'b010000011011111;
		Coeff[2710] <= 15'b010000011100010;
		Coeff[2711] <= 15'b010000011100101;
		Coeff[2712] <= 15'b010000011101000;
		Coeff[2713] <= 15'b010000011101011;
		Coeff[2714] <= 15'b010000011101110;
		Coeff[2715] <= 15'b010000011110001;
		Coeff[2716] <= 15'b010000011110100;
		Coeff[2717] <= 15'b010000011111000;
		Coeff[2718] <= 15'b010000011111011;
		Coeff[2719] <= 15'b010000011111110;
		Coeff[2720] <= 15'b010000100000001;
		Coeff[2721] <= 15'b010000100000100;
		Coeff[2722] <= 15'b010000100000111;
		Coeff[2723] <= 15'b010000100001010;
		Coeff[2724] <= 15'b010000100001101;
		Coeff[2725] <= 15'b010000100010000;
		Coeff[2726] <= 15'b010000100010011;
		Coeff[2727] <= 15'b010000100010110;
		Coeff[2728] <= 15'b010000100011001;
		Coeff[2729] <= 15'b010000100011100;
		Coeff[2730] <= 15'b010000100011111;
		Coeff[2731] <= 15'b010000100100010;
		Coeff[2732] <= 15'b010000100100101;
		Coeff[2733] <= 15'b010000100101000;
		Coeff[2734] <= 15'b010000100101011;
		Coeff[2735] <= 15'b010000100101110;
		Coeff[2736] <= 15'b010000100110001;
		Coeff[2737] <= 15'b010000100110100;
		Coeff[2738] <= 15'b010000100110111;
		Coeff[2739] <= 15'b010000100111010;
		Coeff[2740] <= 15'b010000100111101;
		Coeff[2741] <= 15'b010000101000000;
		Coeff[2742] <= 15'b010000101000011;
		Coeff[2743] <= 15'b010000101000110;
		Coeff[2744] <= 15'b010000101001001;
		Coeff[2745] <= 15'b010000101001100;
		Coeff[2746] <= 15'b010000101010000;
		Coeff[2747] <= 15'b010000101010011;
		Coeff[2748] <= 15'b010000101010110;
		Coeff[2749] <= 15'b010000101011001;
		Coeff[2750] <= 15'b010000101011100;
		Coeff[2751] <= 15'b010000101011111;
		Coeff[2752] <= 15'b010000101100010;
		Coeff[2753] <= 15'b010000101100101;
		Coeff[2754] <= 15'b010000101101000;
		Coeff[2755] <= 15'b010000101101011;
		Coeff[2756] <= 15'b010000101101110;
		Coeff[2757] <= 15'b010000101110001;
		Coeff[2758] <= 15'b010000101110100;
		Coeff[2759] <= 15'b010000101110111;
		Coeff[2760] <= 15'b010000101111010;
		Coeff[2761] <= 15'b010000101111101;
		Coeff[2762] <= 15'b010000110000000;
		Coeff[2763] <= 15'b010000110000011;
		Coeff[2764] <= 15'b010000110000110;
		Coeff[2765] <= 15'b010000110001001;
		Coeff[2766] <= 15'b010000110001100;
		Coeff[2767] <= 15'b010000110001111;
		Coeff[2768] <= 15'b010000110010010;
		Coeff[2769] <= 15'b010000110010101;
		Coeff[2770] <= 15'b010000110011000;
		Coeff[2771] <= 15'b010000110011011;
		Coeff[2772] <= 15'b010000110011110;
		Coeff[2773] <= 15'b010000110100001;
		Coeff[2774] <= 15'b010000110100100;
		Coeff[2775] <= 15'b010000110100111;
		Coeff[2776] <= 15'b010000110101010;
		Coeff[2777] <= 15'b010000110101101;
		Coeff[2778] <= 15'b010000110110001;
		Coeff[2779] <= 15'b010000110110100;
		Coeff[2780] <= 15'b010000110110111;
		Coeff[2781] <= 15'b010000110111010;
		Coeff[2782] <= 15'b010000110111101;
		Coeff[2783] <= 15'b010000111000000;
		Coeff[2784] <= 15'b010000111000011;
		Coeff[2785] <= 15'b010000111000110;
		Coeff[2786] <= 15'b010000111001001;
		Coeff[2787] <= 15'b010000111001100;
		Coeff[2788] <= 15'b010000111001111;
		Coeff[2789] <= 15'b010000111010010;
		Coeff[2790] <= 15'b010000111010101;
		Coeff[2791] <= 15'b010000111011000;
		Coeff[2792] <= 15'b010000111011011;
		Coeff[2793] <= 15'b010000111011110;
		Coeff[2794] <= 15'b010000111100001;
		Coeff[2795] <= 15'b010000111100100;
		Coeff[2796] <= 15'b010000111100111;
		Coeff[2797] <= 15'b010000111101010;
		Coeff[2798] <= 15'b010000111101101;
		Coeff[2799] <= 15'b010000111110000;
		Coeff[2800] <= 15'b010000111110011;
		Coeff[2801] <= 15'b010000111110110;
		Coeff[2802] <= 15'b010000111111001;
		Coeff[2803] <= 15'b010000111111100;
		Coeff[2804] <= 15'b010000111111111;
		Coeff[2805] <= 15'b010001000000010;
		Coeff[2806] <= 15'b010001000000101;
		Coeff[2807] <= 15'b010001000001000;
		Coeff[2808] <= 15'b010001000001011;
		Coeff[2809] <= 15'b010001000001110;
		Coeff[2810] <= 15'b010001000010001;
		Coeff[2811] <= 15'b010001000010101;
		Coeff[2812] <= 15'b010001000011000;
		Coeff[2813] <= 15'b010001000011011;
		Coeff[2814] <= 15'b010001000011110;
		Coeff[2815] <= 15'b010001000100001;
		Coeff[2816] <= 15'b010001000100100;
		Coeff[2817] <= 15'b010001000100111;
		Coeff[2818] <= 15'b010001000101010;
		Coeff[2819] <= 15'b010001000101101;
		Coeff[2820] <= 15'b010001000110000;
		Coeff[2821] <= 15'b010001000110011;
		Coeff[2822] <= 15'b010001000110110;
		Coeff[2823] <= 15'b010001000111001;
		Coeff[2824] <= 15'b010001000111100;
		Coeff[2825] <= 15'b010001000111111;
		Coeff[2826] <= 15'b010001001000010;
		Coeff[2827] <= 15'b010001001000101;
		Coeff[2828] <= 15'b010001001001000;
		Coeff[2829] <= 15'b010001001001011;
		Coeff[2830] <= 15'b010001001001110;
		Coeff[2831] <= 15'b010001001010001;
		Coeff[2832] <= 15'b010001001010100;
		Coeff[2833] <= 15'b010001001010111;
		Coeff[2834] <= 15'b010001001011010;
		Coeff[2835] <= 15'b010001001011101;
		Coeff[2836] <= 15'b010001001100000;
		Coeff[2837] <= 15'b010001001100011;
		Coeff[2838] <= 15'b010001001100110;
		Coeff[2839] <= 15'b010001001101001;
		Coeff[2840] <= 15'b010001001101100;
		Coeff[2841] <= 15'b010001001101111;
		Coeff[2842] <= 15'b010001001110010;
		Coeff[2843] <= 15'b010001001110101;
		Coeff[2844] <= 15'b010001001111000;
		Coeff[2845] <= 15'b010001001111011;
		Coeff[2846] <= 15'b010001001111110;
		Coeff[2847] <= 15'b010001010000001;
		Coeff[2848] <= 15'b010001010000100;
		Coeff[2849] <= 15'b010001010001000;
		Coeff[2850] <= 15'b010001010001011;
		Coeff[2851] <= 15'b010001010001110;
		Coeff[2852] <= 15'b010001010010001;
		Coeff[2853] <= 15'b010001010010100;
		Coeff[2854] <= 15'b010001010010111;
		Coeff[2855] <= 15'b010001010011010;
		Coeff[2856] <= 15'b010001010011101;
		Coeff[2857] <= 15'b010001010100000;
		Coeff[2858] <= 15'b010001010100011;
		Coeff[2859] <= 15'b010001010100110;
		Coeff[2860] <= 15'b010001010101001;
		Coeff[2861] <= 15'b010001010101100;
		Coeff[2862] <= 15'b010001010101111;
		Coeff[2863] <= 15'b010001010110010;
		Coeff[2864] <= 15'b010001010110101;
		Coeff[2865] <= 15'b010001010111000;
		Coeff[2866] <= 15'b010001010111011;
		Coeff[2867] <= 15'b010001010111110;
		Coeff[2868] <= 15'b010001011000001;
		Coeff[2869] <= 15'b010001011000100;
		Coeff[2870] <= 15'b010001011000111;
		Coeff[2871] <= 15'b010001011001010;
		Coeff[2872] <= 15'b010001011001101;
		Coeff[2873] <= 15'b010001011010000;
		Coeff[2874] <= 15'b010001011010011;
		Coeff[2875] <= 15'b010001011010110;
		Coeff[2876] <= 15'b010001011011001;
		Coeff[2877] <= 15'b010001011011100;
		Coeff[2878] <= 15'b010001011011111;
		Coeff[2879] <= 15'b010001011100010;
		Coeff[2880] <= 15'b010001011100101;
		Coeff[2881] <= 15'b010001011101000;
		Coeff[2882] <= 15'b010001011101011;
		Coeff[2883] <= 15'b010001011101110;
		Coeff[2884] <= 15'b010001011110001;
		Coeff[2885] <= 15'b010001011110100;
		Coeff[2886] <= 15'b010001011110111;
		Coeff[2887] <= 15'b010001011111010;
		Coeff[2888] <= 15'b010001011111101;
		Coeff[2889] <= 15'b010001100000000;
		Coeff[2890] <= 15'b010001100000011;
		Coeff[2891] <= 15'b010001100000111;
		Coeff[2892] <= 15'b010001100001010;
		Coeff[2893] <= 15'b010001100001101;
		Coeff[2894] <= 15'b010001100010000;
		Coeff[2895] <= 15'b010001100010011;
		Coeff[2896] <= 15'b010001100010110;
		Coeff[2897] <= 15'b010001100011001;
		Coeff[2898] <= 15'b010001100011100;
		Coeff[2899] <= 15'b010001100011111;
		Coeff[2900] <= 15'b010001100100010;
		Coeff[2901] <= 15'b010001100100101;
		Coeff[2902] <= 15'b010001100101000;
		Coeff[2903] <= 15'b010001100101011;
		Coeff[2904] <= 15'b010001100101110;
		Coeff[2905] <= 15'b010001100110001;
		Coeff[2906] <= 15'b010001100110100;
		Coeff[2907] <= 15'b010001100110111;
		Coeff[2908] <= 15'b010001100111010;
		Coeff[2909] <= 15'b010001100111101;
		Coeff[2910] <= 15'b010001101000000;
		Coeff[2911] <= 15'b010001101000011;
		Coeff[2912] <= 15'b010001101000110;
		Coeff[2913] <= 15'b010001101001001;
		Coeff[2914] <= 15'b010001101001100;
		Coeff[2915] <= 15'b010001101001111;
		Coeff[2916] <= 15'b010001101010010;
		Coeff[2917] <= 15'b010001101010101;
		Coeff[2918] <= 15'b010001101011000;
		Coeff[2919] <= 15'b010001101011011;
		Coeff[2920] <= 15'b010001101011110;
		Coeff[2921] <= 15'b010001101100001;
		Coeff[2922] <= 15'b010001101100100;
		Coeff[2923] <= 15'b010001101100111;
		Coeff[2924] <= 15'b010001101101010;
		Coeff[2925] <= 15'b010001101101101;
		Coeff[2926] <= 15'b010001101110000;
		Coeff[2927] <= 15'b010001101110011;
		Coeff[2928] <= 15'b010001101110110;
		Coeff[2929] <= 15'b010001101111001;
		Coeff[2930] <= 15'b010001101111100;
		Coeff[2931] <= 15'b010001101111111;
		Coeff[2932] <= 15'b010001110000010;
		Coeff[2933] <= 15'b010001110000101;
		Coeff[2934] <= 15'b010001110001000;
		Coeff[2935] <= 15'b010001110001011;
		Coeff[2936] <= 15'b010001110001110;
		Coeff[2937] <= 15'b010001110010001;
		Coeff[2938] <= 15'b010001110010100;
		Coeff[2939] <= 15'b010001110010111;
		Coeff[2940] <= 15'b010001110011010;
		Coeff[2941] <= 15'b010001110011101;
		Coeff[2942] <= 15'b010001110100000;
		Coeff[2943] <= 15'b010001110100100;
		Coeff[2944] <= 15'b010001110100111;
		Coeff[2945] <= 15'b010001110101010;
		Coeff[2946] <= 15'b010001110101101;
		Coeff[2947] <= 15'b010001110110000;
		Coeff[2948] <= 15'b010001110110011;
		Coeff[2949] <= 15'b010001110110110;
		Coeff[2950] <= 15'b010001110111001;
		Coeff[2951] <= 15'b010001110111100;
		Coeff[2952] <= 15'b010001110111111;
		Coeff[2953] <= 15'b010001111000010;
		Coeff[2954] <= 15'b010001111000101;
		Coeff[2955] <= 15'b010001111001000;
		Coeff[2956] <= 15'b010001111001011;
		Coeff[2957] <= 15'b010001111001110;
		Coeff[2958] <= 15'b010001111010001;
		Coeff[2959] <= 15'b010001111010100;
		Coeff[2960] <= 15'b010001111010111;
		Coeff[2961] <= 15'b010001111011010;
		Coeff[2962] <= 15'b010001111011101;
		Coeff[2963] <= 15'b010001111100000;
		Coeff[2964] <= 15'b010001111100011;
		Coeff[2965] <= 15'b010001111100110;
		Coeff[2966] <= 15'b010001111101001;
		Coeff[2967] <= 15'b010001111101100;
		Coeff[2968] <= 15'b010001111101111;
		Coeff[2969] <= 15'b010001111110010;
		Coeff[2970] <= 15'b010001111110101;
		Coeff[2971] <= 15'b010001111111000;
		Coeff[2972] <= 15'b010001111111011;
		Coeff[2973] <= 15'b010001111111110;
		Coeff[2974] <= 15'b010010000000001;
		Coeff[2975] <= 15'b010010000000100;
		Coeff[2976] <= 15'b010010000000111;
		Coeff[2977] <= 15'b010010000001010;
		Coeff[2978] <= 15'b010010000001101;
		Coeff[2979] <= 15'b010010000010000;
		Coeff[2980] <= 15'b010010000010011;
		Coeff[2981] <= 15'b010010000010110;
		Coeff[2982] <= 15'b010010000011001;
		Coeff[2983] <= 15'b010010000011100;
		Coeff[2984] <= 15'b010010000011111;
		Coeff[2985] <= 15'b010010000100010;
		Coeff[2986] <= 15'b010010000100101;
		Coeff[2987] <= 15'b010010000101000;
		Coeff[2988] <= 15'b010010000101011;
		Coeff[2989] <= 15'b010010000101110;
		Coeff[2990] <= 15'b010010000110001;
		Coeff[2991] <= 15'b010010000110100;
		Coeff[2992] <= 15'b010010000110111;
		Coeff[2993] <= 15'b010010000111010;
		Coeff[2994] <= 15'b010010000111101;
		Coeff[2995] <= 15'b010010001000000;
		Coeff[2996] <= 15'b010010001000011;
		Coeff[2997] <= 15'b010010001000110;
		Coeff[2998] <= 15'b010010001001001;
		Coeff[2999] <= 15'b010010001001100;
		Coeff[3000] <= 15'b010010001001111;
		Coeff[3001] <= 15'b010010001010010;
		Coeff[3002] <= 15'b010010001010101;
		Coeff[3003] <= 15'b010010001011000;
		Coeff[3004] <= 15'b010010001011011;
		Coeff[3005] <= 15'b010010001011110;
		Coeff[3006] <= 15'b010010001100001;
		Coeff[3007] <= 15'b010010001100100;
		Coeff[3008] <= 15'b010010001100111;
		Coeff[3009] <= 15'b010010001101010;
		Coeff[3010] <= 15'b010010001101101;
		Coeff[3011] <= 15'b010010001110001;
		Coeff[3012] <= 15'b010010001110100;
		Coeff[3013] <= 15'b010010001110111;
		Coeff[3014] <= 15'b010010001111010;
		Coeff[3015] <= 15'b010010001111101;
		Coeff[3016] <= 15'b010010010000000;
		Coeff[3017] <= 15'b010010010000011;
		Coeff[3018] <= 15'b010010010000110;
		Coeff[3019] <= 15'b010010010001001;
		Coeff[3020] <= 15'b010010010001100;
		Coeff[3021] <= 15'b010010010001111;
		Coeff[3022] <= 15'b010010010010010;
		Coeff[3023] <= 15'b010010010010101;
		Coeff[3024] <= 15'b010010010011000;
		Coeff[3025] <= 15'b010010010011011;
		Coeff[3026] <= 15'b010010010011110;
		Coeff[3027] <= 15'b010010010100001;
		Coeff[3028] <= 15'b010010010100100;
		Coeff[3029] <= 15'b010010010100111;
		Coeff[3030] <= 15'b010010010101010;
		Coeff[3031] <= 15'b010010010101101;
		Coeff[3032] <= 15'b010010010110000;
		Coeff[3033] <= 15'b010010010110011;
		Coeff[3034] <= 15'b010010010110110;
		Coeff[3035] <= 15'b010010010111001;
		Coeff[3036] <= 15'b010010010111100;
		Coeff[3037] <= 15'b010010010111111;
		Coeff[3038] <= 15'b010010011000010;
		Coeff[3039] <= 15'b010010011000101;
		Coeff[3040] <= 15'b010010011001000;
		Coeff[3041] <= 15'b010010011001011;
		Coeff[3042] <= 15'b010010011001110;
		Coeff[3043] <= 15'b010010011010001;
		Coeff[3044] <= 15'b010010011010100;
		Coeff[3045] <= 15'b010010011010111;
		Coeff[3046] <= 15'b010010011011010;
		Coeff[3047] <= 15'b010010011011101;
		Coeff[3048] <= 15'b010010011100000;
		Coeff[3049] <= 15'b010010011100011;
		Coeff[3050] <= 15'b010010011100110;
		Coeff[3051] <= 15'b010010011101001;
		Coeff[3052] <= 15'b010010011101100;
		Coeff[3053] <= 15'b010010011101111;
		Coeff[3054] <= 15'b010010011110010;
		Coeff[3055] <= 15'b010010011110101;
		Coeff[3056] <= 15'b010010011111000;
		Coeff[3057] <= 15'b010010011111011;
		Coeff[3058] <= 15'b010010011111110;
		Coeff[3059] <= 15'b010010100000001;
		Coeff[3060] <= 15'b010010100000100;
		Coeff[3061] <= 15'b010010100000111;
		Coeff[3062] <= 15'b010010100001010;
		Coeff[3063] <= 15'b010010100001101;
		Coeff[3064] <= 15'b010010100010000;
		Coeff[3065] <= 15'b010010100010011;
		Coeff[3066] <= 15'b010010100010110;
		Coeff[3067] <= 15'b010010100011001;
		Coeff[3068] <= 15'b010010100011100;
		Coeff[3069] <= 15'b010010100011111;
		Coeff[3070] <= 15'b010010100100010;
		Coeff[3071] <= 15'b010010100100101;
		Coeff[3072] <= 15'b010010100101000;
		Coeff[3073] <= 15'b010010100101011;
		Coeff[3074] <= 15'b010010100101110;
		Coeff[3075] <= 15'b010010100110001;
		Coeff[3076] <= 15'b010010100110100;
		Coeff[3077] <= 15'b010010100110111;
		Coeff[3078] <= 15'b010010100111010;
		Coeff[3079] <= 15'b010010100111101;
		Coeff[3080] <= 15'b010010101000000;
		Coeff[3081] <= 15'b010010101000011;
		Coeff[3082] <= 15'b010010101000110;
		Coeff[3083] <= 15'b010010101001001;
		Coeff[3084] <= 15'b010010101001100;
		Coeff[3085] <= 15'b010010101001111;
		Coeff[3086] <= 15'b010010101010010;
		Coeff[3087] <= 15'b010010101010101;
		Coeff[3088] <= 15'b010010101011000;
		Coeff[3089] <= 15'b010010101011011;
		Coeff[3090] <= 15'b010010101011110;
		Coeff[3091] <= 15'b010010101100001;
		Coeff[3092] <= 15'b010010101100100;
		Coeff[3093] <= 15'b010010101100111;
		Coeff[3094] <= 15'b010010101101010;
		Coeff[3095] <= 15'b010010101101101;
		Coeff[3096] <= 15'b010010101110000;
		Coeff[3097] <= 15'b010010101110011;
		Coeff[3098] <= 15'b010010101110110;
		Coeff[3099] <= 15'b010010101111001;
		Coeff[3100] <= 15'b010010101111100;
		Coeff[3101] <= 15'b010010101111111;
		Coeff[3102] <= 15'b010010110000010;
		Coeff[3103] <= 15'b010010110000101;
		Coeff[3104] <= 15'b010010110001000;
		Coeff[3105] <= 15'b010010110001011;
		Coeff[3106] <= 15'b010010110001110;
		Coeff[3107] <= 15'b010010110010001;
		Coeff[3108] <= 15'b010010110010100;
		Coeff[3109] <= 15'b010010110010111;
		Coeff[3110] <= 15'b010010110011010;
		Coeff[3111] <= 15'b010010110011101;
		Coeff[3112] <= 15'b010010110100000;
		Coeff[3113] <= 15'b010010110100011;
		Coeff[3114] <= 15'b010010110100110;
		Coeff[3115] <= 15'b010010110101001;
		Coeff[3116] <= 15'b010010110101100;
		Coeff[3117] <= 15'b010010110101111;
		Coeff[3118] <= 15'b010010110110010;
		Coeff[3119] <= 15'b010010110110101;
		Coeff[3120] <= 15'b010010110111000;
		Coeff[3121] <= 15'b010010110111011;
		Coeff[3122] <= 15'b010010110111110;
		Coeff[3123] <= 15'b010010111000001;
		Coeff[3124] <= 15'b010010111000100;
		Coeff[3125] <= 15'b010010111000111;
		Coeff[3126] <= 15'b010010111001010;
		Coeff[3127] <= 15'b010010111001101;
		Coeff[3128] <= 15'b010010111010000;
		Coeff[3129] <= 15'b010010111010011;
		Coeff[3130] <= 15'b010010111010110;
		Coeff[3131] <= 15'b010010111011001;
		Coeff[3132] <= 15'b010010111011100;
		Coeff[3133] <= 15'b010010111011111;
		Coeff[3134] <= 15'b010010111100010;
		Coeff[3135] <= 15'b010010111100101;
		Coeff[3136] <= 15'b010010111101000;
		Coeff[3137] <= 15'b010010111101011;
		Coeff[3138] <= 15'b010010111101110;
		Coeff[3139] <= 15'b010010111110001;
		Coeff[3140] <= 15'b010010111110100;
		Coeff[3141] <= 15'b010010111110111;
		Coeff[3142] <= 15'b010010111111010;
		Coeff[3143] <= 15'b010010111111101;
		Coeff[3144] <= 15'b010011000000000;
		Coeff[3145] <= 15'b010011000000011;
		Coeff[3146] <= 15'b010011000000110;
		Coeff[3147] <= 15'b010011000001001;
		Coeff[3148] <= 15'b010011000001100;
		Coeff[3149] <= 15'b010011000001111;
		Coeff[3150] <= 15'b010011000010010;
		Coeff[3151] <= 15'b010011000010101;
		Coeff[3152] <= 15'b010011000011000;
		Coeff[3153] <= 15'b010011000011011;
		Coeff[3154] <= 15'b010011000011110;
		Coeff[3155] <= 15'b010011000100001;
		Coeff[3156] <= 15'b010011000100100;
		Coeff[3157] <= 15'b010011000100111;
		Coeff[3158] <= 15'b010011000101010;
		Coeff[3159] <= 15'b010011000101101;
		Coeff[3160] <= 15'b010011000110000;
		Coeff[3161] <= 15'b010011000110011;
		Coeff[3162] <= 15'b010011000110110;
		Coeff[3163] <= 15'b010011000111001;
		Coeff[3164] <= 15'b010011000111100;
		Coeff[3165] <= 15'b010011000111111;
		Coeff[3166] <= 15'b010011001000010;
		Coeff[3167] <= 15'b010011001000101;
		Coeff[3168] <= 15'b010011001001000;
		Coeff[3169] <= 15'b010011001001011;
		Coeff[3170] <= 15'b010011001001110;
		Coeff[3171] <= 15'b010011001010001;
		Coeff[3172] <= 15'b010011001010100;
		Coeff[3173] <= 15'b010011001010111;
		Coeff[3174] <= 15'b010011001011010;
		Coeff[3175] <= 15'b010011001011101;
		Coeff[3176] <= 15'b010011001100000;
		Coeff[3177] <= 15'b010011001100011;
		Coeff[3178] <= 15'b010011001100110;
		Coeff[3179] <= 15'b010011001101001;
		Coeff[3180] <= 15'b010011001101100;
		Coeff[3181] <= 15'b010011001101111;
		Coeff[3182] <= 15'b010011001110010;
		Coeff[3183] <= 15'b010011001110101;
		Coeff[3184] <= 15'b010011001111000;
		Coeff[3185] <= 15'b010011001111011;
		Coeff[3186] <= 15'b010011001111110;
		Coeff[3187] <= 15'b010011010000001;
		Coeff[3188] <= 15'b010011010000100;
		Coeff[3189] <= 15'b010011010000111;
		Coeff[3190] <= 15'b010011010001010;
		Coeff[3191] <= 15'b010011010001101;
		Coeff[3192] <= 15'b010011010010000;
		Coeff[3193] <= 15'b010011010010011;
		Coeff[3194] <= 15'b010011010010110;
		Coeff[3195] <= 15'b010011010011001;
		Coeff[3196] <= 15'b010011010011100;
		Coeff[3197] <= 15'b010011010011111;
		Coeff[3198] <= 15'b010011010100010;
		Coeff[3199] <= 15'b010011010100101;
		Coeff[3200] <= 15'b010011010101000;
		Coeff[3201] <= 15'b010011010101011;
		Coeff[3202] <= 15'b010011010101110;
		Coeff[3203] <= 15'b010011010110001;
		Coeff[3204] <= 15'b010011010110100;
		Coeff[3205] <= 15'b010011010110111;
		Coeff[3206] <= 15'b010011010111010;
		Coeff[3207] <= 15'b010011010111101;
		Coeff[3208] <= 15'b010011011000000;
		Coeff[3209] <= 15'b010011011000011;
		Coeff[3210] <= 15'b010011011000110;
		Coeff[3211] <= 15'b010011011001001;
		Coeff[3212] <= 15'b010011011001100;
		Coeff[3213] <= 15'b010011011001111;
		Coeff[3214] <= 15'b010011011010010;
		Coeff[3215] <= 15'b010011011010101;
		Coeff[3216] <= 15'b010011011011000;
		Coeff[3217] <= 15'b010011011011011;
		Coeff[3218] <= 15'b010011011011110;
		Coeff[3219] <= 15'b010011011100001;
		Coeff[3220] <= 15'b010011011100100;
		Coeff[3221] <= 15'b010011011100111;
		Coeff[3222] <= 15'b010011011101010;
		Coeff[3223] <= 15'b010011011101101;
		Coeff[3224] <= 15'b010011011110000;
		Coeff[3225] <= 15'b010011011110011;
		Coeff[3226] <= 15'b010011011110110;
		Coeff[3227] <= 15'b010011011111001;
		Coeff[3228] <= 15'b010011011111100;
		Coeff[3229] <= 15'b010011011111111;
		Coeff[3230] <= 15'b010011100000010;
		Coeff[3231] <= 15'b010011100000101;
		Coeff[3232] <= 15'b010011100001000;
		Coeff[3233] <= 15'b010011100001011;
		Coeff[3234] <= 15'b010011100001110;
		Coeff[3235] <= 15'b010011100010001;
		Coeff[3236] <= 15'b010011100010100;
		Coeff[3237] <= 15'b010011100010111;
		Coeff[3238] <= 15'b010011100011010;
		Coeff[3239] <= 15'b010011100011101;
		Coeff[3240] <= 15'b010011100100000;
		Coeff[3241] <= 15'b010011100100011;
		Coeff[3242] <= 15'b010011100100110;
		Coeff[3243] <= 15'b010011100101001;
		Coeff[3244] <= 15'b010011100101100;
		Coeff[3245] <= 15'b010011100101111;
		Coeff[3246] <= 15'b010011100110010;
		Coeff[3247] <= 15'b010011100110101;
		Coeff[3248] <= 15'b010011100111000;
		Coeff[3249] <= 15'b010011100111011;
		Coeff[3250] <= 15'b010011100111110;
		Coeff[3251] <= 15'b010011101000001;
		Coeff[3252] <= 15'b010011101000100;
		Coeff[3253] <= 15'b010011101000111;
		Coeff[3254] <= 15'b010011101001010;
		Coeff[3255] <= 15'b010011101001101;
		Coeff[3256] <= 15'b010011101010000;
		Coeff[3257] <= 15'b010011101010011;
		Coeff[3258] <= 15'b010011101010110;
		Coeff[3259] <= 15'b010011101011001;
		Coeff[3260] <= 15'b010011101011100;
		Coeff[3261] <= 15'b010011101011111;
		Coeff[3262] <= 15'b010011101100010;
		Coeff[3263] <= 15'b010011101100101;
		Coeff[3264] <= 15'b010011101101000;
		Coeff[3265] <= 15'b010011101101011;
		Coeff[3266] <= 15'b010011101101110;
		Coeff[3267] <= 15'b010011101110001;
		Coeff[3268] <= 15'b010011101110100;
		Coeff[3269] <= 15'b010011101110111;
		Coeff[3270] <= 15'b010011101111010;
		Coeff[3271] <= 15'b010011101111101;
		Coeff[3272] <= 15'b010011110000000;
		Coeff[3273] <= 15'b010011110000011;
		Coeff[3274] <= 15'b010011110000110;
		Coeff[3275] <= 15'b010011110001000;
		Coeff[3276] <= 15'b010011110001011;
		Coeff[3277] <= 15'b010011110001110;
		Coeff[3278] <= 15'b010011110010001;
		Coeff[3279] <= 15'b010011110010100;
		Coeff[3280] <= 15'b010011110010111;
		Coeff[3281] <= 15'b010011110011010;
		Coeff[3282] <= 15'b010011110011101;
		Coeff[3283] <= 15'b010011110100000;
		Coeff[3284] <= 15'b010011110100011;
		Coeff[3285] <= 15'b010011110100110;
		Coeff[3286] <= 15'b010011110101001;
		Coeff[3287] <= 15'b010011110101100;
		Coeff[3288] <= 15'b010011110101111;
		Coeff[3289] <= 15'b010011110110010;
		Coeff[3290] <= 15'b010011110110101;
		Coeff[3291] <= 15'b010011110111000;
		Coeff[3292] <= 15'b010011110111011;
		Coeff[3293] <= 15'b010011110111110;
		Coeff[3294] <= 15'b010011111000001;
		Coeff[3295] <= 15'b010011111000100;
		Coeff[3296] <= 15'b010011111000111;
		Coeff[3297] <= 15'b010011111001010;
		Coeff[3298] <= 15'b010011111001101;
		Coeff[3299] <= 15'b010011111010000;
		Coeff[3300] <= 15'b010011111010011;
		Coeff[3301] <= 15'b010011111010110;
		Coeff[3302] <= 15'b010011111011001;
		Coeff[3303] <= 15'b010011111011100;
		Coeff[3304] <= 15'b010011111011111;
		Coeff[3305] <= 15'b010011111100010;
		Coeff[3306] <= 15'b010011111100101;
		Coeff[3307] <= 15'b010011111101000;
		Coeff[3308] <= 15'b010011111101011;
		Coeff[3309] <= 15'b010011111101110;
		Coeff[3310] <= 15'b010011111110001;
		Coeff[3311] <= 15'b010011111110100;
		Coeff[3312] <= 15'b010011111110111;
		Coeff[3313] <= 15'b010011111111010;
		Coeff[3314] <= 15'b010011111111101;
		Coeff[3315] <= 15'b010100000000000;
		Coeff[3316] <= 15'b010100000000011;
		Coeff[3317] <= 15'b010100000000110;
		Coeff[3318] <= 15'b010100000001001;
		Coeff[3319] <= 15'b010100000001100;
		Coeff[3320] <= 15'b010100000001111;
		Coeff[3321] <= 15'b010100000010010;
		Coeff[3322] <= 15'b010100000010101;
		Coeff[3323] <= 15'b010100000011000;
		Coeff[3324] <= 15'b010100000011011;
		Coeff[3325] <= 15'b010100000011110;
		Coeff[3326] <= 15'b010100000100001;
		Coeff[3327] <= 15'b010100000100100;
		Coeff[3328] <= 15'b010100000100111;
		Coeff[3329] <= 15'b010100000101010;
		Coeff[3330] <= 15'b010100000101101;
		Coeff[3331] <= 15'b010100000110000;
		Coeff[3332] <= 15'b010100000110011;
		Coeff[3333] <= 15'b010100000110110;
		Coeff[3334] <= 15'b010100000111001;
		Coeff[3335] <= 15'b010100000111100;
		Coeff[3336] <= 15'b010100000111111;
		Coeff[3337] <= 15'b010100001000010;
		Coeff[3338] <= 15'b010100001000101;
		Coeff[3339] <= 15'b010100001001000;
		Coeff[3340] <= 15'b010100001001011;
		Coeff[3341] <= 15'b010100001001101;
		Coeff[3342] <= 15'b010100001010000;
		Coeff[3343] <= 15'b010100001010011;
		Coeff[3344] <= 15'b010100001010110;
		Coeff[3345] <= 15'b010100001011001;
		Coeff[3346] <= 15'b010100001011100;
		Coeff[3347] <= 15'b010100001011111;
		Coeff[3348] <= 15'b010100001100010;
		Coeff[3349] <= 15'b010100001100101;
		Coeff[3350] <= 15'b010100001101000;
		Coeff[3351] <= 15'b010100001101011;
		Coeff[3352] <= 15'b010100001101110;
		Coeff[3353] <= 15'b010100001110001;
		Coeff[3354] <= 15'b010100001110100;
		Coeff[3355] <= 15'b010100001110111;
		Coeff[3356] <= 15'b010100001111010;
		Coeff[3357] <= 15'b010100001111101;
		Coeff[3358] <= 15'b010100010000000;
		Coeff[3359] <= 15'b010100010000011;
		Coeff[3360] <= 15'b010100010000110;
		Coeff[3361] <= 15'b010100010001001;
		Coeff[3362] <= 15'b010100010001100;
		Coeff[3363] <= 15'b010100010001111;
		Coeff[3364] <= 15'b010100010010010;
		Coeff[3365] <= 15'b010100010010101;
		Coeff[3366] <= 15'b010100010011000;
		Coeff[3367] <= 15'b010100010011011;
		Coeff[3368] <= 15'b010100010011110;
		Coeff[3369] <= 15'b010100010100001;
		Coeff[3370] <= 15'b010100010100100;
		Coeff[3371] <= 15'b010100010100111;
		Coeff[3372] <= 15'b010100010101010;
		Coeff[3373] <= 15'b010100010101101;
		Coeff[3374] <= 15'b010100010110000;
		Coeff[3375] <= 15'b010100010110011;
		Coeff[3376] <= 15'b010100010110110;
		Coeff[3377] <= 15'b010100010111001;
		Coeff[3378] <= 15'b010100010111100;
		Coeff[3379] <= 15'b010100010111111;
		Coeff[3380] <= 15'b010100011000010;
		Coeff[3381] <= 15'b010100011000101;
		Coeff[3382] <= 15'b010100011001000;
		Coeff[3383] <= 15'b010100011001011;
		Coeff[3384] <= 15'b010100011001110;
		Coeff[3385] <= 15'b010100011010001;
		Coeff[3386] <= 15'b010100011010100;
		Coeff[3387] <= 15'b010100011010111;
		Coeff[3388] <= 15'b010100011011010;
		Coeff[3389] <= 15'b010100011011101;
		Coeff[3390] <= 15'b010100011011111;
		Coeff[3391] <= 15'b010100011100010;
		Coeff[3392] <= 15'b010100011100101;
		Coeff[3393] <= 15'b010100011101000;
		Coeff[3394] <= 15'b010100011101011;
		Coeff[3395] <= 15'b010100011101110;
		Coeff[3396] <= 15'b010100011110001;
		Coeff[3397] <= 15'b010100011110100;
		Coeff[3398] <= 15'b010100011110111;
		Coeff[3399] <= 15'b010100011111010;
		Coeff[3400] <= 15'b010100011111101;
		Coeff[3401] <= 15'b010100100000000;
		Coeff[3402] <= 15'b010100100000011;
		Coeff[3403] <= 15'b010100100000110;
		Coeff[3404] <= 15'b010100100001001;
		Coeff[3405] <= 15'b010100100001100;
		Coeff[3406] <= 15'b010100100001111;
		Coeff[3407] <= 15'b010100100010010;
		Coeff[3408] <= 15'b010100100010101;
		Coeff[3409] <= 15'b010100100011000;
		Coeff[3410] <= 15'b010100100011011;
		Coeff[3411] <= 15'b010100100011110;
		Coeff[3412] <= 15'b010100100100001;
		Coeff[3413] <= 15'b010100100100100;
		Coeff[3414] <= 15'b010100100100111;
		Coeff[3415] <= 15'b010100100101010;
		Coeff[3416] <= 15'b010100100101101;
		Coeff[3417] <= 15'b010100100110000;
		Coeff[3418] <= 15'b010100100110011;
		Coeff[3419] <= 15'b010100100110110;
		Coeff[3420] <= 15'b010100100111001;
		Coeff[3421] <= 15'b010100100111100;
		Coeff[3422] <= 15'b010100100111111;
		Coeff[3423] <= 15'b010100101000010;
		Coeff[3424] <= 15'b010100101000101;
		Coeff[3425] <= 15'b010100101001000;
		Coeff[3426] <= 15'b010100101001011;
		Coeff[3427] <= 15'b010100101001110;
		Coeff[3428] <= 15'b010100101010001;
		Coeff[3429] <= 15'b010100101010100;
		Coeff[3430] <= 15'b010100101010110;
		Coeff[3431] <= 15'b010100101011001;
		Coeff[3432] <= 15'b010100101011100;
		Coeff[3433] <= 15'b010100101011111;
		Coeff[3434] <= 15'b010100101100010;
		Coeff[3435] <= 15'b010100101100101;
		Coeff[3436] <= 15'b010100101101000;
		Coeff[3437] <= 15'b010100101101011;
		Coeff[3438] <= 15'b010100101101110;
		Coeff[3439] <= 15'b010100101110001;
		Coeff[3440] <= 15'b010100101110100;
		Coeff[3441] <= 15'b010100101110111;
		Coeff[3442] <= 15'b010100101111010;
		Coeff[3443] <= 15'b010100101111101;
		Coeff[3444] <= 15'b010100110000000;
		Coeff[3445] <= 15'b010100110000011;
		Coeff[3446] <= 15'b010100110000110;
		Coeff[3447] <= 15'b010100110001001;
		Coeff[3448] <= 15'b010100110001100;
		Coeff[3449] <= 15'b010100110001111;
		Coeff[3450] <= 15'b010100110010010;
		Coeff[3451] <= 15'b010100110010101;
		Coeff[3452] <= 15'b010100110011000;
		Coeff[3453] <= 15'b010100110011011;
		Coeff[3454] <= 15'b010100110011110;
		Coeff[3455] <= 15'b010100110100001;
		Coeff[3456] <= 15'b010100110100100;
		Coeff[3457] <= 15'b010100110100111;
		Coeff[3458] <= 15'b010100110101010;
		Coeff[3459] <= 15'b010100110101101;
		Coeff[3460] <= 15'b010100110110000;
		Coeff[3461] <= 15'b010100110110011;
		Coeff[3462] <= 15'b010100110110110;
		Coeff[3463] <= 15'b010100110111001;
		Coeff[3464] <= 15'b010100110111100;
		Coeff[3465] <= 15'b010100110111111;
		Coeff[3466] <= 15'b010100111000001;
		Coeff[3467] <= 15'b010100111000100;
		Coeff[3468] <= 15'b010100111000111;
		Coeff[3469] <= 15'b010100111001010;
		Coeff[3470] <= 15'b010100111001101;
		Coeff[3471] <= 15'b010100111010000;
		Coeff[3472] <= 15'b010100111010011;
		Coeff[3473] <= 15'b010100111010110;
		Coeff[3474] <= 15'b010100111011001;
		Coeff[3475] <= 15'b010100111011100;
		Coeff[3476] <= 15'b010100111011111;
		Coeff[3477] <= 15'b010100111100010;
		Coeff[3478] <= 15'b010100111100101;
		Coeff[3479] <= 15'b010100111101000;
		Coeff[3480] <= 15'b010100111101011;
		Coeff[3481] <= 15'b010100111101110;
		Coeff[3482] <= 15'b010100111110001;
		Coeff[3483] <= 15'b010100111110100;
		Coeff[3484] <= 15'b010100111110111;
		Coeff[3485] <= 15'b010100111111010;
		Coeff[3486] <= 15'b010100111111101;
		Coeff[3487] <= 15'b010101000000000;
		Coeff[3488] <= 15'b010101000000011;
		Coeff[3489] <= 15'b010101000000110;
		Coeff[3490] <= 15'b010101000001001;
		Coeff[3491] <= 15'b010101000001100;
		Coeff[3492] <= 15'b010101000001111;
		Coeff[3493] <= 15'b010101000010010;
		Coeff[3494] <= 15'b010101000010101;
		Coeff[3495] <= 15'b010101000011000;
		Coeff[3496] <= 15'b010101000011011;
		Coeff[3497] <= 15'b010101000011101;
		Coeff[3498] <= 15'b010101000100000;
		Coeff[3499] <= 15'b010101000100011;
		Coeff[3500] <= 15'b010101000100110;
		Coeff[3501] <= 15'b010101000101001;
		Coeff[3502] <= 15'b010101000101100;
		Coeff[3503] <= 15'b010101000101111;
		Coeff[3504] <= 15'b010101000110010;
		Coeff[3505] <= 15'b010101000110101;
		Coeff[3506] <= 15'b010101000111000;
		Coeff[3507] <= 15'b010101000111011;
		Coeff[3508] <= 15'b010101000111110;
		Coeff[3509] <= 15'b010101001000001;
		Coeff[3510] <= 15'b010101001000100;
		Coeff[3511] <= 15'b010101001000111;
		Coeff[3512] <= 15'b010101001001010;
		Coeff[3513] <= 15'b010101001001101;
		Coeff[3514] <= 15'b010101001010000;
		Coeff[3515] <= 15'b010101001010011;
		Coeff[3516] <= 15'b010101001010110;
		Coeff[3517] <= 15'b010101001011001;
		Coeff[3518] <= 15'b010101001011100;
		Coeff[3519] <= 15'b010101001011111;
		Coeff[3520] <= 15'b010101001100010;
		Coeff[3521] <= 15'b010101001100101;
		Coeff[3522] <= 15'b010101001101000;
		Coeff[3523] <= 15'b010101001101011;
		Coeff[3524] <= 15'b010101001101110;
		Coeff[3525] <= 15'b010101001110001;
		Coeff[3526] <= 15'b010101001110011;
		Coeff[3527] <= 15'b010101001110110;
		Coeff[3528] <= 15'b010101001111001;
		Coeff[3529] <= 15'b010101001111100;
		Coeff[3530] <= 15'b010101001111111;
		Coeff[3531] <= 15'b010101010000010;
		Coeff[3532] <= 15'b010101010000101;
		Coeff[3533] <= 15'b010101010001000;
		Coeff[3534] <= 15'b010101010001011;
		Coeff[3535] <= 15'b010101010001110;
		Coeff[3536] <= 15'b010101010010001;
		Coeff[3537] <= 15'b010101010010100;
		Coeff[3538] <= 15'b010101010010111;
		Coeff[3539] <= 15'b010101010011010;
		Coeff[3540] <= 15'b010101010011101;
		Coeff[3541] <= 15'b010101010100000;
		Coeff[3542] <= 15'b010101010100011;
		Coeff[3543] <= 15'b010101010100110;
		Coeff[3544] <= 15'b010101010101001;
		Coeff[3545] <= 15'b010101010101100;
		Coeff[3546] <= 15'b010101010101111;
		Coeff[3547] <= 15'b010101010110010;
		Coeff[3548] <= 15'b010101010110101;
		Coeff[3549] <= 15'b010101010111000;
		Coeff[3550] <= 15'b010101010111011;
		Coeff[3551] <= 15'b010101010111110;
		Coeff[3552] <= 15'b010101011000001;
		Coeff[3553] <= 15'b010101011000011;
		Coeff[3554] <= 15'b010101011000110;
		Coeff[3555] <= 15'b010101011001001;
		Coeff[3556] <= 15'b010101011001100;
		Coeff[3557] <= 15'b010101011001111;
		Coeff[3558] <= 15'b010101011010010;
		Coeff[3559] <= 15'b010101011010101;
		Coeff[3560] <= 15'b010101011011000;
		Coeff[3561] <= 15'b010101011011011;
		Coeff[3562] <= 15'b010101011011110;
		Coeff[3563] <= 15'b010101011100001;
		Coeff[3564] <= 15'b010101011100100;
		Coeff[3565] <= 15'b010101011100111;
		Coeff[3566] <= 15'b010101011101010;
		Coeff[3567] <= 15'b010101011101101;
		Coeff[3568] <= 15'b010101011110000;
		Coeff[3569] <= 15'b010101011110011;
		Coeff[3570] <= 15'b010101011110110;
		Coeff[3571] <= 15'b010101011111001;
		Coeff[3572] <= 15'b010101011111100;
		Coeff[3573] <= 15'b010101011111111;
		Coeff[3574] <= 15'b010101100000010;
		Coeff[3575] <= 15'b010101100000101;
		Coeff[3576] <= 15'b010101100001000;
		Coeff[3577] <= 15'b010101100001010;
		Coeff[3578] <= 15'b010101100001101;
		Coeff[3579] <= 15'b010101100010000;
		Coeff[3580] <= 15'b010101100010011;
		Coeff[3581] <= 15'b010101100010110;
		Coeff[3582] <= 15'b010101100011001;
		Coeff[3583] <= 15'b010101100011100;
		Coeff[3584] <= 15'b010101100011111;
		Coeff[3585] <= 15'b010101100100010;
		Coeff[3586] <= 15'b010101100100101;
		Coeff[3587] <= 15'b010101100101000;
		Coeff[3588] <= 15'b010101100101011;
		Coeff[3589] <= 15'b010101100101110;
		Coeff[3590] <= 15'b010101100110001;
		Coeff[3591] <= 15'b010101100110100;
		Coeff[3592] <= 15'b010101100110111;
		Coeff[3593] <= 15'b010101100111010;
		Coeff[3594] <= 15'b010101100111101;
		Coeff[3595] <= 15'b010101101000000;
		Coeff[3596] <= 15'b010101101000011;
		Coeff[3597] <= 15'b010101101000110;
		Coeff[3598] <= 15'b010101101001001;
		Coeff[3599] <= 15'b010101101001100;
		Coeff[3600] <= 15'b010101101001111;
		Coeff[3601] <= 15'b010101101010001;
		Coeff[3602] <= 15'b010101101010100;
		Coeff[3603] <= 15'b010101101010111;
		Coeff[3604] <= 15'b010101101011010;
		Coeff[3605] <= 15'b010101101011101;
		Coeff[3606] <= 15'b010101101100000;
		Coeff[3607] <= 15'b010101101100011;
		Coeff[3608] <= 15'b010101101100110;
		Coeff[3609] <= 15'b010101101101001;
		Coeff[3610] <= 15'b010101101101100;
		Coeff[3611] <= 15'b010101101101111;
		Coeff[3612] <= 15'b010101101110010;
		Coeff[3613] <= 15'b010101101110101;
		Coeff[3614] <= 15'b010101101111000;
		Coeff[3615] <= 15'b010101101111011;
		Coeff[3616] <= 15'b010101101111110;
		Coeff[3617] <= 15'b010101110000001;
		Coeff[3618] <= 15'b010101110000100;
		Coeff[3619] <= 15'b010101110000111;
		Coeff[3620] <= 15'b010101110001010;
		Coeff[3621] <= 15'b010101110001101;
		Coeff[3622] <= 15'b010101110010000;
		Coeff[3623] <= 15'b010101110010010;
		Coeff[3624] <= 15'b010101110010101;
		Coeff[3625] <= 15'b010101110011000;
		Coeff[3626] <= 15'b010101110011011;
		Coeff[3627] <= 15'b010101110011110;
		Coeff[3628] <= 15'b010101110100001;
		Coeff[3629] <= 15'b010101110100100;
		Coeff[3630] <= 15'b010101110100111;
		Coeff[3631] <= 15'b010101110101010;
		Coeff[3632] <= 15'b010101110101101;
		Coeff[3633] <= 15'b010101110110000;
		Coeff[3634] <= 15'b010101110110011;
		Coeff[3635] <= 15'b010101110110110;
		Coeff[3636] <= 15'b010101110111001;
		Coeff[3637] <= 15'b010101110111100;
		Coeff[3638] <= 15'b010101110111111;
		Coeff[3639] <= 15'b010101111000010;
		Coeff[3640] <= 15'b010101111000101;
		Coeff[3641] <= 15'b010101111001000;
		Coeff[3642] <= 15'b010101111001011;
		Coeff[3643] <= 15'b010101111001110;
		Coeff[3644] <= 15'b010101111010000;
		Coeff[3645] <= 15'b010101111010011;
		Coeff[3646] <= 15'b010101111010110;
		Coeff[3647] <= 15'b010101111011001;
		Coeff[3648] <= 15'b010101111011100;
		Coeff[3649] <= 15'b010101111011111;
		Coeff[3650] <= 15'b010101111100010;
		Coeff[3651] <= 15'b010101111100101;
		Coeff[3652] <= 15'b010101111101000;
		Coeff[3653] <= 15'b010101111101011;
		Coeff[3654] <= 15'b010101111101110;
		Coeff[3655] <= 15'b010101111110001;
		Coeff[3656] <= 15'b010101111110100;
		Coeff[3657] <= 15'b010101111110111;
		Coeff[3658] <= 15'b010101111111010;
		Coeff[3659] <= 15'b010101111111101;
		Coeff[3660] <= 15'b010110000000000;
		Coeff[3661] <= 15'b010110000000011;
		Coeff[3662] <= 15'b010110000000110;
		Coeff[3663] <= 15'b010110000001001;
		Coeff[3664] <= 15'b010110000001100;
		Coeff[3665] <= 15'b010110000001110;
		Coeff[3666] <= 15'b010110000010001;
		Coeff[3667] <= 15'b010110000010100;
		Coeff[3668] <= 15'b010110000010111;
		Coeff[3669] <= 15'b010110000011010;
		Coeff[3670] <= 15'b010110000011101;
		Coeff[3671] <= 15'b010110000100000;
		Coeff[3672] <= 15'b010110000100011;
		Coeff[3673] <= 15'b010110000100110;
		Coeff[3674] <= 15'b010110000101001;
		Coeff[3675] <= 15'b010110000101100;
		Coeff[3676] <= 15'b010110000101111;
		Coeff[3677] <= 15'b010110000110010;
		Coeff[3678] <= 15'b010110000110101;
		Coeff[3679] <= 15'b010110000111000;
		Coeff[3680] <= 15'b010110000111011;
		Coeff[3681] <= 15'b010110000111110;
		Coeff[3682] <= 15'b010110001000001;
		Coeff[3683] <= 15'b010110001000100;
		Coeff[3684] <= 15'b010110001000110;
		Coeff[3685] <= 15'b010110001001001;
		Coeff[3686] <= 15'b010110001001100;
		Coeff[3687] <= 15'b010110001001111;
		Coeff[3688] <= 15'b010110001010010;
		Coeff[3689] <= 15'b010110001010101;
		Coeff[3690] <= 15'b010110001011000;
		Coeff[3691] <= 15'b010110001011011;
		Coeff[3692] <= 15'b010110001011110;
		Coeff[3693] <= 15'b010110001100001;
		Coeff[3694] <= 15'b010110001100100;
		Coeff[3695] <= 15'b010110001100111;
		Coeff[3696] <= 15'b010110001101010;
		Coeff[3697] <= 15'b010110001101101;
		Coeff[3698] <= 15'b010110001110000;
		Coeff[3699] <= 15'b010110001110011;
		Coeff[3700] <= 15'b010110001110110;
		Coeff[3701] <= 15'b010110001111001;
		Coeff[3702] <= 15'b010110001111100;
		Coeff[3703] <= 15'b010110001111110;
		Coeff[3704] <= 15'b010110010000001;
		Coeff[3705] <= 15'b010110010000100;
		Coeff[3706] <= 15'b010110010000111;
		Coeff[3707] <= 15'b010110010001010;
		Coeff[3708] <= 15'b010110010001101;
		Coeff[3709] <= 15'b010110010010000;
		Coeff[3710] <= 15'b010110010010011;
		Coeff[3711] <= 15'b010110010010110;
		Coeff[3712] <= 15'b010110010011001;
		Coeff[3713] <= 15'b010110010011100;
		Coeff[3714] <= 15'b010110010011111;
		Coeff[3715] <= 15'b010110010100010;
		Coeff[3716] <= 15'b010110010100101;
		Coeff[3717] <= 15'b010110010101000;
		Coeff[3718] <= 15'b010110010101011;
		Coeff[3719] <= 15'b010110010101110;
		Coeff[3720] <= 15'b010110010110001;
		Coeff[3721] <= 15'b010110010110011;
		Coeff[3722] <= 15'b010110010110110;
		Coeff[3723] <= 15'b010110010111001;
		Coeff[3724] <= 15'b010110010111100;
		Coeff[3725] <= 15'b010110010111111;
		Coeff[3726] <= 15'b010110011000010;
		Coeff[3727] <= 15'b010110011000101;
		Coeff[3728] <= 15'b010110011001000;
		Coeff[3729] <= 15'b010110011001011;
		Coeff[3730] <= 15'b010110011001110;
		Coeff[3731] <= 15'b010110011010001;
		Coeff[3732] <= 15'b010110011010100;
		Coeff[3733] <= 15'b010110011010111;
		Coeff[3734] <= 15'b010110011011010;
		Coeff[3735] <= 15'b010110011011101;
		Coeff[3736] <= 15'b010110011100000;
		Coeff[3737] <= 15'b010110011100011;
		Coeff[3738] <= 15'b010110011100110;
		Coeff[3739] <= 15'b010110011101000;
		Coeff[3740] <= 15'b010110011101011;
		Coeff[3741] <= 15'b010110011101110;
		Coeff[3742] <= 15'b010110011110001;
		Coeff[3743] <= 15'b010110011110100;
		Coeff[3744] <= 15'b010110011110111;
		Coeff[3745] <= 15'b010110011111010;
		Coeff[3746] <= 15'b010110011111101;
		Coeff[3747] <= 15'b010110100000000;
		Coeff[3748] <= 15'b010110100000011;
		Coeff[3749] <= 15'b010110100000110;
		Coeff[3750] <= 15'b010110100001001;
		Coeff[3751] <= 15'b010110100001100;
		Coeff[3752] <= 15'b010110100001111;
		Coeff[3753] <= 15'b010110100010010;
		Coeff[3754] <= 15'b010110100010101;
		Coeff[3755] <= 15'b010110100011000;
		Coeff[3756] <= 15'b010110100011010;
		Coeff[3757] <= 15'b010110100011101;
		Coeff[3758] <= 15'b010110100100000;
		Coeff[3759] <= 15'b010110100100011;
		Coeff[3760] <= 15'b010110100100110;
		Coeff[3761] <= 15'b010110100101001;
		Coeff[3762] <= 15'b010110100101100;
		Coeff[3763] <= 15'b010110100101111;
		Coeff[3764] <= 15'b010110100110010;
		Coeff[3765] <= 15'b010110100110101;
		Coeff[3766] <= 15'b010110100111000;
		Coeff[3767] <= 15'b010110100111011;
		Coeff[3768] <= 15'b010110100111110;
		Coeff[3769] <= 15'b010110101000001;
		Coeff[3770] <= 15'b010110101000100;
		Coeff[3771] <= 15'b010110101000111;
		Coeff[3772] <= 15'b010110101001001;
		Coeff[3773] <= 15'b010110101001100;
		Coeff[3774] <= 15'b010110101001111;
		Coeff[3775] <= 15'b010110101010010;
		Coeff[3776] <= 15'b010110101010101;
		Coeff[3777] <= 15'b010110101011000;
		Coeff[3778] <= 15'b010110101011011;
		Coeff[3779] <= 15'b010110101011110;
		Coeff[3780] <= 15'b010110101100001;
		Coeff[3781] <= 15'b010110101100100;
		Coeff[3782] <= 15'b010110101100111;
		Coeff[3783] <= 15'b010110101101010;
		Coeff[3784] <= 15'b010110101101101;
		Coeff[3785] <= 15'b010110101110000;
		Coeff[3786] <= 15'b010110101110011;
		Coeff[3787] <= 15'b010110101110110;
		Coeff[3788] <= 15'b010110101111000;
		Coeff[3789] <= 15'b010110101111011;
		Coeff[3790] <= 15'b010110101111110;
		Coeff[3791] <= 15'b010110110000001;
		Coeff[3792] <= 15'b010110110000100;
		Coeff[3793] <= 15'b010110110000111;
		Coeff[3794] <= 15'b010110110001010;
		Coeff[3795] <= 15'b010110110001101;
		Coeff[3796] <= 15'b010110110010000;
		Coeff[3797] <= 15'b010110110010011;
		Coeff[3798] <= 15'b010110110010110;
		Coeff[3799] <= 15'b010110110011001;
		Coeff[3800] <= 15'b010110110011100;
		Coeff[3801] <= 15'b010110110011111;
		Coeff[3802] <= 15'b010110110100010;
		Coeff[3803] <= 15'b010110110100101;
		Coeff[3804] <= 15'b010110110100111;
		Coeff[3805] <= 15'b010110110101010;
		Coeff[3806] <= 15'b010110110101101;
		Coeff[3807] <= 15'b010110110110000;
		Coeff[3808] <= 15'b010110110110011;
		Coeff[3809] <= 15'b010110110110110;
		Coeff[3810] <= 15'b010110110111001;
		Coeff[3811] <= 15'b010110110111100;
		Coeff[3812] <= 15'b010110110111111;
		Coeff[3813] <= 15'b010110111000010;
		Coeff[3814] <= 15'b010110111000101;
		Coeff[3815] <= 15'b010110111001000;
		Coeff[3816] <= 15'b010110111001011;
		Coeff[3817] <= 15'b010110111001110;
		Coeff[3818] <= 15'b010110111010001;
		Coeff[3819] <= 15'b010110111010011;
		Coeff[3820] <= 15'b010110111010110;
		Coeff[3821] <= 15'b010110111011001;
		Coeff[3822] <= 15'b010110111011100;
		Coeff[3823] <= 15'b010110111011111;
		Coeff[3824] <= 15'b010110111100010;
		Coeff[3825] <= 15'b010110111100101;
		Coeff[3826] <= 15'b010110111101000;
		Coeff[3827] <= 15'b010110111101011;
		Coeff[3828] <= 15'b010110111101110;
		Coeff[3829] <= 15'b010110111110001;
		Coeff[3830] <= 15'b010110111110100;
		Coeff[3831] <= 15'b010110111110111;
		Coeff[3832] <= 15'b010110111111010;
		Coeff[3833] <= 15'b010110111111101;
		Coeff[3834] <= 15'b010110111111111;
		Coeff[3835] <= 15'b010111000000010;
		Coeff[3836] <= 15'b010111000000101;
		Coeff[3837] <= 15'b010111000001000;
		Coeff[3838] <= 15'b010111000001011;
		Coeff[3839] <= 15'b010111000001110;
		Coeff[3840] <= 15'b010111000010001;
		Coeff[3841] <= 15'b010111000010100;
		Coeff[3842] <= 15'b010111000010111;
		Coeff[3843] <= 15'b010111000011010;
		Coeff[3844] <= 15'b010111000011101;
		Coeff[3845] <= 15'b010111000100000;
		Coeff[3846] <= 15'b010111000100011;
		Coeff[3847] <= 15'b010111000100110;
		Coeff[3848] <= 15'b010111000101000;
		Coeff[3849] <= 15'b010111000101011;
		Coeff[3850] <= 15'b010111000101110;
		Coeff[3851] <= 15'b010111000110001;
		Coeff[3852] <= 15'b010111000110100;
		Coeff[3853] <= 15'b010111000110111;
		Coeff[3854] <= 15'b010111000111010;
		Coeff[3855] <= 15'b010111000111101;
		Coeff[3856] <= 15'b010111001000000;
		Coeff[3857] <= 15'b010111001000011;
		Coeff[3858] <= 15'b010111001000110;
		Coeff[3859] <= 15'b010111001001001;
		Coeff[3860] <= 15'b010111001001100;
		Coeff[3861] <= 15'b010111001001111;
		Coeff[3862] <= 15'b010111001010001;
		Coeff[3863] <= 15'b010111001010100;
		Coeff[3864] <= 15'b010111001010111;
		Coeff[3865] <= 15'b010111001011010;
		Coeff[3866] <= 15'b010111001011101;
		Coeff[3867] <= 15'b010111001100000;
		Coeff[3868] <= 15'b010111001100011;
		Coeff[3869] <= 15'b010111001100110;
		Coeff[3870] <= 15'b010111001101001;
		Coeff[3871] <= 15'b010111001101100;
		Coeff[3872] <= 15'b010111001101111;
		Coeff[3873] <= 15'b010111001110010;
		Coeff[3874] <= 15'b010111001110101;
		Coeff[3875] <= 15'b010111001111000;
		Coeff[3876] <= 15'b010111001111010;
		Coeff[3877] <= 15'b010111001111101;
		Coeff[3878] <= 15'b010111010000000;
		Coeff[3879] <= 15'b010111010000011;
		Coeff[3880] <= 15'b010111010000110;
		Coeff[3881] <= 15'b010111010001001;
		Coeff[3882] <= 15'b010111010001100;
		Coeff[3883] <= 15'b010111010001111;
		Coeff[3884] <= 15'b010111010010010;
		Coeff[3885] <= 15'b010111010010101;
		Coeff[3886] <= 15'b010111010011000;
		Coeff[3887] <= 15'b010111010011011;
		Coeff[3888] <= 15'b010111010011110;
		Coeff[3889] <= 15'b010111010100001;
		Coeff[3890] <= 15'b010111010100011;
		Coeff[3891] <= 15'b010111010100110;
		Coeff[3892] <= 15'b010111010101001;
		Coeff[3893] <= 15'b010111010101100;
		Coeff[3894] <= 15'b010111010101111;
		Coeff[3895] <= 15'b010111010110010;
		Coeff[3896] <= 15'b010111010110101;
		Coeff[3897] <= 15'b010111010111000;
		Coeff[3898] <= 15'b010111010111011;
		Coeff[3899] <= 15'b010111010111110;
		Coeff[3900] <= 15'b010111011000001;
		Coeff[3901] <= 15'b010111011000100;
		Coeff[3902] <= 15'b010111011000111;
		Coeff[3903] <= 15'b010111011001001;
		Coeff[3904] <= 15'b010111011001100;
		Coeff[3905] <= 15'b010111011001111;
		Coeff[3906] <= 15'b010111011010010;
		Coeff[3907] <= 15'b010111011010101;
		Coeff[3908] <= 15'b010111011011000;
		Coeff[3909] <= 15'b010111011011011;
		Coeff[3910] <= 15'b010111011011110;
		Coeff[3911] <= 15'b010111011100001;
		Coeff[3912] <= 15'b010111011100100;
		Coeff[3913] <= 15'b010111011100111;
		Coeff[3914] <= 15'b010111011101010;
		Coeff[3915] <= 15'b010111011101101;
		Coeff[3916] <= 15'b010111011101111;
		Coeff[3917] <= 15'b010111011110010;
		Coeff[3918] <= 15'b010111011110101;
		Coeff[3919] <= 15'b010111011111000;
		Coeff[3920] <= 15'b010111011111011;
		Coeff[3921] <= 15'b010111011111110;
		Coeff[3922] <= 15'b010111100000001;
		Coeff[3923] <= 15'b010111100000100;
		Coeff[3924] <= 15'b010111100000111;
		Coeff[3925] <= 15'b010111100001010;
		Coeff[3926] <= 15'b010111100001101;
		Coeff[3927] <= 15'b010111100010000;
		Coeff[3928] <= 15'b010111100010011;
		Coeff[3929] <= 15'b010111100010101;
		Coeff[3930] <= 15'b010111100011000;
		Coeff[3931] <= 15'b010111100011011;
		Coeff[3932] <= 15'b010111100011110;
		Coeff[3933] <= 15'b010111100100001;
		Coeff[3934] <= 15'b010111100100100;
		Coeff[3935] <= 15'b010111100100111;
		Coeff[3936] <= 15'b010111100101010;
		Coeff[3937] <= 15'b010111100101101;
		Coeff[3938] <= 15'b010111100110000;
		Coeff[3939] <= 15'b010111100110011;
		Coeff[3940] <= 15'b010111100110110;
		Coeff[3941] <= 15'b010111100111001;
		Coeff[3942] <= 15'b010111100111011;
		Coeff[3943] <= 15'b010111100111110;
		Coeff[3944] <= 15'b010111101000001;
		Coeff[3945] <= 15'b010111101000100;
		Coeff[3946] <= 15'b010111101000111;
		Coeff[3947] <= 15'b010111101001010;
		Coeff[3948] <= 15'b010111101001101;
		Coeff[3949] <= 15'b010111101010000;
		Coeff[3950] <= 15'b010111101010011;
		Coeff[3951] <= 15'b010111101010110;
		Coeff[3952] <= 15'b010111101011001;
		Coeff[3953] <= 15'b010111101011100;
		Coeff[3954] <= 15'b010111101011110;
		Coeff[3955] <= 15'b010111101100001;
		Coeff[3956] <= 15'b010111101100100;
		Coeff[3957] <= 15'b010111101100111;
		Coeff[3958] <= 15'b010111101101010;
		Coeff[3959] <= 15'b010111101101101;
		Coeff[3960] <= 15'b010111101110000;
		Coeff[3961] <= 15'b010111101110011;
		Coeff[3962] <= 15'b010111101110110;
		Coeff[3963] <= 15'b010111101111001;
		Coeff[3964] <= 15'b010111101111100;
		Coeff[3965] <= 15'b010111101111111;
		Coeff[3966] <= 15'b010111110000001;
		Coeff[3967] <= 15'b010111110000100;
		Coeff[3968] <= 15'b010111110000111;
		Coeff[3969] <= 15'b010111110001010;
		Coeff[3970] <= 15'b010111110001101;
		Coeff[3971] <= 15'b010111110010000;
		Coeff[3972] <= 15'b010111110010011;
		Coeff[3973] <= 15'b010111110010110;
		Coeff[3974] <= 15'b010111110011001;
		Coeff[3975] <= 15'b010111110011100;
		Coeff[3976] <= 15'b010111110011111;
		Coeff[3977] <= 15'b010111110100010;
		Coeff[3978] <= 15'b010111110100100;
		Coeff[3979] <= 15'b010111110100111;
		Coeff[3980] <= 15'b010111110101010;
		Coeff[3981] <= 15'b010111110101101;
		Coeff[3982] <= 15'b010111110110000;
		Coeff[3983] <= 15'b010111110110011;
		Coeff[3984] <= 15'b010111110110110;
		Coeff[3985] <= 15'b010111110111001;
		Coeff[3986] <= 15'b010111110111100;
		Coeff[3987] <= 15'b010111110111111;
		Coeff[3988] <= 15'b010111111000010;
		Coeff[3989] <= 15'b010111111000101;
		Coeff[3990] <= 15'b010111111000111;
		Coeff[3991] <= 15'b010111111001010;
		Coeff[3992] <= 15'b010111111001101;
		Coeff[3993] <= 15'b010111111010000;
		Coeff[3994] <= 15'b010111111010011;
		Coeff[3995] <= 15'b010111111010110;
		Coeff[3996] <= 15'b010111111011001;
		Coeff[3997] <= 15'b010111111011100;
		Coeff[3998] <= 15'b010111111011111;
		Coeff[3999] <= 15'b010111111100010;
		Coeff[4000] <= 15'b010111111100101;
		Coeff[4001] <= 15'b010111111101000;
		Coeff[4002] <= 15'b010111111101010;
		Coeff[4003] <= 15'b010111111101101;
		Coeff[4004] <= 15'b010111111110000;
		Coeff[4005] <= 15'b010111111110011;
		Coeff[4006] <= 15'b010111111110110;
		Coeff[4007] <= 15'b010111111111001;
		Coeff[4008] <= 15'b010111111111100;
		Coeff[4009] <= 15'b010111111111111;
		Coeff[4010] <= 15'b011000000000010;
		Coeff[4011] <= 15'b011000000000101;
		Coeff[4012] <= 15'b011000000001000;
		Coeff[4013] <= 15'b011000000001010;
		Coeff[4014] <= 15'b011000000001101;
		Coeff[4015] <= 15'b011000000010000;
		Coeff[4016] <= 15'b011000000010011;
		Coeff[4017] <= 15'b011000000010110;
		Coeff[4018] <= 15'b011000000011001;
		Coeff[4019] <= 15'b011000000011100;
		Coeff[4020] <= 15'b011000000011111;
		Coeff[4021] <= 15'b011000000100010;
		Coeff[4022] <= 15'b011000000100101;
		Coeff[4023] <= 15'b011000000101000;
		Coeff[4024] <= 15'b011000000101010;
		Coeff[4025] <= 15'b011000000101101;
		Coeff[4026] <= 15'b011000000110000;
		Coeff[4027] <= 15'b011000000110011;
		Coeff[4028] <= 15'b011000000110110;
		Coeff[4029] <= 15'b011000000111001;
		Coeff[4030] <= 15'b011000000111100;
		Coeff[4031] <= 15'b011000000111111;
		Coeff[4032] <= 15'b011000001000010;
		Coeff[4033] <= 15'b011000001000101;
		Coeff[4034] <= 15'b011000001001000;
		Coeff[4035] <= 15'b011000001001011;
		Coeff[4036] <= 15'b011000001001101;
		Coeff[4037] <= 15'b011000001010000;
		Coeff[4038] <= 15'b011000001010011;
		Coeff[4039] <= 15'b011000001010110;
		Coeff[4040] <= 15'b011000001011001;
		Coeff[4041] <= 15'b011000001011100;
		Coeff[4042] <= 15'b011000001011111;
		Coeff[4043] <= 15'b011000001100010;
		Coeff[4044] <= 15'b011000001100101;
		Coeff[4045] <= 15'b011000001101000;
		Coeff[4046] <= 15'b011000001101011;
		Coeff[4047] <= 15'b011000001101101;
		Coeff[4048] <= 15'b011000001110000;
		Coeff[4049] <= 15'b011000001110011;
		Coeff[4050] <= 15'b011000001110110;
		Coeff[4051] <= 15'b011000001111001;
		Coeff[4052] <= 15'b011000001111100;
		Coeff[4053] <= 15'b011000001111111;
		Coeff[4054] <= 15'b011000010000010;
		Coeff[4055] <= 15'b011000010000101;
		Coeff[4056] <= 15'b011000010001000;
		Coeff[4057] <= 15'b011000010001010;
		Coeff[4058] <= 15'b011000010001101;
		Coeff[4059] <= 15'b011000010010000;
		Coeff[4060] <= 15'b011000010010011;
		Coeff[4061] <= 15'b011000010010110;
		Coeff[4062] <= 15'b011000010011001;
		Coeff[4063] <= 15'b011000010011100;
		Coeff[4064] <= 15'b011000010011111;
		Coeff[4065] <= 15'b011000010100010;
		Coeff[4066] <= 15'b011000010100101;
		Coeff[4067] <= 15'b011000010101000;
		Coeff[4068] <= 15'b011000010101010;
		Coeff[4069] <= 15'b011000010101101;
		Coeff[4070] <= 15'b011000010110000;
		Coeff[4071] <= 15'b011000010110011;
		Coeff[4072] <= 15'b011000010110110;
		Coeff[4073] <= 15'b011000010111001;
		Coeff[4074] <= 15'b011000010111100;
		Coeff[4075] <= 15'b011000010111111;
		Coeff[4076] <= 15'b011000011000010;
		Coeff[4077] <= 15'b011000011000101;
		Coeff[4078] <= 15'b011000011001000;
		Coeff[4079] <= 15'b011000011001010;
		Coeff[4080] <= 15'b011000011001101;
		Coeff[4081] <= 15'b011000011010000;
		Coeff[4082] <= 15'b011000011010011;
		Coeff[4083] <= 15'b011000011010110;
		Coeff[4084] <= 15'b011000011011001;
		Coeff[4085] <= 15'b011000011011100;
		Coeff[4086] <= 15'b011000011011111;
		Coeff[4087] <= 15'b011000011100010;
		Coeff[4088] <= 15'b011000011100101;
		Coeff[4089] <= 15'b011000011100111;
		Coeff[4090] <= 15'b011000011101010;
		Coeff[4091] <= 15'b011000011101101;
		Coeff[4092] <= 15'b011000011110000;
		Coeff[4093] <= 15'b011000011110011;
		Coeff[4094] <= 15'b011000011110110;
		Coeff[4095] <= 15'b011000011111001;
		Coeff[4096] <= 15'b011000011111100;
		Coeff[4097] <= 15'b011000011111111;
		Coeff[4098] <= 15'b011000100000010;
		Coeff[4099] <= 15'b011000100000100;
		Coeff[4100] <= 15'b011000100000111;
		Coeff[4101] <= 15'b011000100001010;
		Coeff[4102] <= 15'b011000100001101;
		Coeff[4103] <= 15'b011000100010000;
		Coeff[4104] <= 15'b011000100010011;
		Coeff[4105] <= 15'b011000100010110;
		Coeff[4106] <= 15'b011000100011001;
		Coeff[4107] <= 15'b011000100011100;
		Coeff[4108] <= 15'b011000100011111;
		Coeff[4109] <= 15'b011000100100001;
		Coeff[4110] <= 15'b011000100100100;
		Coeff[4111] <= 15'b011000100100111;
		Coeff[4112] <= 15'b011000100101010;
		Coeff[4113] <= 15'b011000100101101;
		Coeff[4114] <= 15'b011000100110000;
		Coeff[4115] <= 15'b011000100110011;
		Coeff[4116] <= 15'b011000100110110;
		Coeff[4117] <= 15'b011000100111001;
		Coeff[4118] <= 15'b011000100111100;
		Coeff[4119] <= 15'b011000100111110;
		Coeff[4120] <= 15'b011000101000001;
		Coeff[4121] <= 15'b011000101000100;
		Coeff[4122] <= 15'b011000101000111;
		Coeff[4123] <= 15'b011000101001010;
		Coeff[4124] <= 15'b011000101001101;
		Coeff[4125] <= 15'b011000101010000;
		Coeff[4126] <= 15'b011000101010011;
		Coeff[4127] <= 15'b011000101010110;
		Coeff[4128] <= 15'b011000101011001;
		Coeff[4129] <= 15'b011000101011011;
		Coeff[4130] <= 15'b011000101011110;
		Coeff[4131] <= 15'b011000101100001;
		Coeff[4132] <= 15'b011000101100100;
		Coeff[4133] <= 15'b011000101100111;
		Coeff[4134] <= 15'b011000101101010;
		Coeff[4135] <= 15'b011000101101101;
		Coeff[4136] <= 15'b011000101110000;
		Coeff[4137] <= 15'b011000101110011;
		Coeff[4138] <= 15'b011000101110110;
		Coeff[4139] <= 15'b011000101111000;
		Coeff[4140] <= 15'b011000101111011;
		Coeff[4141] <= 15'b011000101111110;
		Coeff[4142] <= 15'b011000110000001;
		Coeff[4143] <= 15'b011000110000100;
		Coeff[4144] <= 15'b011000110000111;
		Coeff[4145] <= 15'b011000110001010;
		Coeff[4146] <= 15'b011000110001101;
		Coeff[4147] <= 15'b011000110010000;
		Coeff[4148] <= 15'b011000110010011;
		Coeff[4149] <= 15'b011000110010101;
		Coeff[4150] <= 15'b011000110011000;
		Coeff[4151] <= 15'b011000110011011;
		Coeff[4152] <= 15'b011000110011110;
		Coeff[4153] <= 15'b011000110100001;
		Coeff[4154] <= 15'b011000110100100;
		Coeff[4155] <= 15'b011000110100111;
		Coeff[4156] <= 15'b011000110101010;
		Coeff[4157] <= 15'b011000110101101;
		Coeff[4158] <= 15'b011000110110000;
		Coeff[4159] <= 15'b011000110110010;
		Coeff[4160] <= 15'b011000110110101;
		Coeff[4161] <= 15'b011000110111000;
		Coeff[4162] <= 15'b011000110111011;
		Coeff[4163] <= 15'b011000110111110;
		Coeff[4164] <= 15'b011000111000001;
		Coeff[4165] <= 15'b011000111000100;
		Coeff[4166] <= 15'b011000111000111;
		Coeff[4167] <= 15'b011000111001010;
		Coeff[4168] <= 15'b011000111001100;
		Coeff[4169] <= 15'b011000111001111;
		Coeff[4170] <= 15'b011000111010010;
		Coeff[4171] <= 15'b011000111010101;
		Coeff[4172] <= 15'b011000111011000;
		Coeff[4173] <= 15'b011000111011011;
		Coeff[4174] <= 15'b011000111011110;
		Coeff[4175] <= 15'b011000111100001;
		Coeff[4176] <= 15'b011000111100100;
		Coeff[4177] <= 15'b011000111100110;
		Coeff[4178] <= 15'b011000111101001;
		Coeff[4179] <= 15'b011000111101100;
		Coeff[4180] <= 15'b011000111101111;
		Coeff[4181] <= 15'b011000111110010;
		Coeff[4182] <= 15'b011000111110101;
		Coeff[4183] <= 15'b011000111111000;
		Coeff[4184] <= 15'b011000111111011;
		Coeff[4185] <= 15'b011000111111110;
		Coeff[4186] <= 15'b011001000000001;
		Coeff[4187] <= 15'b011001000000011;
		Coeff[4188] <= 15'b011001000000110;
		Coeff[4189] <= 15'b011001000001001;
		Coeff[4190] <= 15'b011001000001100;
		Coeff[4191] <= 15'b011001000001111;
		Coeff[4192] <= 15'b011001000010010;
		Coeff[4193] <= 15'b011001000010101;
		Coeff[4194] <= 15'b011001000011000;
		Coeff[4195] <= 15'b011001000011011;
		Coeff[4196] <= 15'b011001000011101;
		Coeff[4197] <= 15'b011001000100000;
		Coeff[4198] <= 15'b011001000100011;
		Coeff[4199] <= 15'b011001000100110;
		Coeff[4200] <= 15'b011001000101001;
		Coeff[4201] <= 15'b011001000101100;
		Coeff[4202] <= 15'b011001000101111;
		Coeff[4203] <= 15'b011001000110010;
		Coeff[4204] <= 15'b011001000110101;
		Coeff[4205] <= 15'b011001000110111;
		Coeff[4206] <= 15'b011001000111010;
		Coeff[4207] <= 15'b011001000111101;
		Coeff[4208] <= 15'b011001001000000;
		Coeff[4209] <= 15'b011001001000011;
		Coeff[4210] <= 15'b011001001000110;
		Coeff[4211] <= 15'b011001001001001;
		Coeff[4212] <= 15'b011001001001100;
		Coeff[4213] <= 15'b011001001001111;
		Coeff[4214] <= 15'b011001001010001;
		Coeff[4215] <= 15'b011001001010100;
		Coeff[4216] <= 15'b011001001010111;
		Coeff[4217] <= 15'b011001001011010;
		Coeff[4218] <= 15'b011001001011101;
		Coeff[4219] <= 15'b011001001100000;
		Coeff[4220] <= 15'b011001001100011;
		Coeff[4221] <= 15'b011001001100110;
		Coeff[4222] <= 15'b011001001101001;
		Coeff[4223] <= 15'b011001001101011;
		Coeff[4224] <= 15'b011001001101110;
		Coeff[4225] <= 15'b011001001110001;
		Coeff[4226] <= 15'b011001001110100;
		Coeff[4227] <= 15'b011001001110111;
		Coeff[4228] <= 15'b011001001111010;
		Coeff[4229] <= 15'b011001001111101;
		Coeff[4230] <= 15'b011001010000000;
		Coeff[4231] <= 15'b011001010000011;
		Coeff[4232] <= 15'b011001010000101;
		Coeff[4233] <= 15'b011001010001000;
		Coeff[4234] <= 15'b011001010001011;
		Coeff[4235] <= 15'b011001010001110;
		Coeff[4236] <= 15'b011001010010001;
		Coeff[4237] <= 15'b011001010010100;
		Coeff[4238] <= 15'b011001010010111;
		Coeff[4239] <= 15'b011001010011010;
		Coeff[4240] <= 15'b011001010011101;
		Coeff[4241] <= 15'b011001010011111;
		Coeff[4242] <= 15'b011001010100010;
		Coeff[4243] <= 15'b011001010100101;
		Coeff[4244] <= 15'b011001010101000;
		Coeff[4245] <= 15'b011001010101011;
		Coeff[4246] <= 15'b011001010101110;
		Coeff[4247] <= 15'b011001010110001;
		Coeff[4248] <= 15'b011001010110100;
		Coeff[4249] <= 15'b011001010110110;
		Coeff[4250] <= 15'b011001010111001;
		Coeff[4251] <= 15'b011001010111100;
		Coeff[4252] <= 15'b011001010111111;
		Coeff[4253] <= 15'b011001011000010;
		Coeff[4254] <= 15'b011001011000101;
		Coeff[4255] <= 15'b011001011001000;
		Coeff[4256] <= 15'b011001011001011;
		Coeff[4257] <= 15'b011001011001110;
		Coeff[4258] <= 15'b011001011010000;
		Coeff[4259] <= 15'b011001011010011;
		Coeff[4260] <= 15'b011001011010110;
		Coeff[4261] <= 15'b011001011011001;
		Coeff[4262] <= 15'b011001011011100;
		Coeff[4263] <= 15'b011001011011111;
		Coeff[4264] <= 15'b011001011100010;
		Coeff[4265] <= 15'b011001011100101;
		Coeff[4266] <= 15'b011001011101000;
		Coeff[4267] <= 15'b011001011101010;
		Coeff[4268] <= 15'b011001011101101;
		Coeff[4269] <= 15'b011001011110000;
		Coeff[4270] <= 15'b011001011110011;
		Coeff[4271] <= 15'b011001011110110;
		Coeff[4272] <= 15'b011001011111001;
		Coeff[4273] <= 15'b011001011111100;
		Coeff[4274] <= 15'b011001011111111;
		Coeff[4275] <= 15'b011001100000001;
		Coeff[4276] <= 15'b011001100000100;
		Coeff[4277] <= 15'b011001100000111;
		Coeff[4278] <= 15'b011001100001010;
		Coeff[4279] <= 15'b011001100001101;
		Coeff[4280] <= 15'b011001100010000;
		Coeff[4281] <= 15'b011001100010011;
		Coeff[4282] <= 15'b011001100010110;
		Coeff[4283] <= 15'b011001100011000;
		Coeff[4284] <= 15'b011001100011011;
		Coeff[4285] <= 15'b011001100011110;
		Coeff[4286] <= 15'b011001100100001;
		Coeff[4287] <= 15'b011001100100100;
		Coeff[4288] <= 15'b011001100100111;
		Coeff[4289] <= 15'b011001100101010;
		Coeff[4290] <= 15'b011001100101101;
		Coeff[4291] <= 15'b011001100110000;
		Coeff[4292] <= 15'b011001100110010;
		Coeff[4293] <= 15'b011001100110101;
		Coeff[4294] <= 15'b011001100111000;
		Coeff[4295] <= 15'b011001100111011;
		Coeff[4296] <= 15'b011001100111110;
		Coeff[4297] <= 15'b011001101000001;
		Coeff[4298] <= 15'b011001101000100;
		Coeff[4299] <= 15'b011001101000111;
		Coeff[4300] <= 15'b011001101001001;
		Coeff[4301] <= 15'b011001101001100;
		Coeff[4302] <= 15'b011001101001111;
		Coeff[4303] <= 15'b011001101010010;
		Coeff[4304] <= 15'b011001101010101;
		Coeff[4305] <= 15'b011001101011000;
		Coeff[4306] <= 15'b011001101011011;
		Coeff[4307] <= 15'b011001101011110;
		Coeff[4308] <= 15'b011001101100000;
		Coeff[4309] <= 15'b011001101100011;
		Coeff[4310] <= 15'b011001101100110;
		Coeff[4311] <= 15'b011001101101001;
		Coeff[4312] <= 15'b011001101101100;
		Coeff[4313] <= 15'b011001101101111;
		Coeff[4314] <= 15'b011001101110010;
		Coeff[4315] <= 15'b011001101110101;
		Coeff[4316] <= 15'b011001101110111;
		Coeff[4317] <= 15'b011001101111010;
		Coeff[4318] <= 15'b011001101111101;
		Coeff[4319] <= 15'b011001110000000;
		Coeff[4320] <= 15'b011001110000011;
		Coeff[4321] <= 15'b011001110000110;
		Coeff[4322] <= 15'b011001110001001;
		Coeff[4323] <= 15'b011001110001100;
		Coeff[4324] <= 15'b011001110001110;
		Coeff[4325] <= 15'b011001110010001;
		Coeff[4326] <= 15'b011001110010100;
		Coeff[4327] <= 15'b011001110010111;
		Coeff[4328] <= 15'b011001110011010;
		Coeff[4329] <= 15'b011001110011101;
		Coeff[4330] <= 15'b011001110100000;
		Coeff[4331] <= 15'b011001110100011;
		Coeff[4332] <= 15'b011001110100101;
		Coeff[4333] <= 15'b011001110101000;
		Coeff[4334] <= 15'b011001110101011;
		Coeff[4335] <= 15'b011001110101110;
		Coeff[4336] <= 15'b011001110110001;
		Coeff[4337] <= 15'b011001110110100;
		Coeff[4338] <= 15'b011001110110111;
		Coeff[4339] <= 15'b011001110111010;
		Coeff[4340] <= 15'b011001110111100;
		Coeff[4341] <= 15'b011001110111111;
		Coeff[4342] <= 15'b011001111000010;
		Coeff[4343] <= 15'b011001111000101;
		Coeff[4344] <= 15'b011001111001000;
		Coeff[4345] <= 15'b011001111001011;
		Coeff[4346] <= 15'b011001111001110;
		Coeff[4347] <= 15'b011001111010001;
		Coeff[4348] <= 15'b011001111010011;
		Coeff[4349] <= 15'b011001111010110;
		Coeff[4350] <= 15'b011001111011001;
		Coeff[4351] <= 15'b011001111011100;
		Coeff[4352] <= 15'b011001111011111;
		Coeff[4353] <= 15'b011001111100010;
		Coeff[4354] <= 15'b011001111100101;
		Coeff[4355] <= 15'b011001111101000;
		Coeff[4356] <= 15'b011001111101010;
		Coeff[4357] <= 15'b011001111101101;
		Coeff[4358] <= 15'b011001111110000;
		Coeff[4359] <= 15'b011001111110011;
		Coeff[4360] <= 15'b011001111110110;
		Coeff[4361] <= 15'b011001111111001;
		Coeff[4362] <= 15'b011001111111100;
		Coeff[4363] <= 15'b011001111111111;
		Coeff[4364] <= 15'b011010000000001;
		Coeff[4365] <= 15'b011010000000100;
		Coeff[4366] <= 15'b011010000000111;
		Coeff[4367] <= 15'b011010000001010;
		Coeff[4368] <= 15'b011010000001101;
		Coeff[4369] <= 15'b011010000010000;
		Coeff[4370] <= 15'b011010000010011;
		Coeff[4371] <= 15'b011010000010101;
		Coeff[4372] <= 15'b011010000011000;
		Coeff[4373] <= 15'b011010000011011;
		Coeff[4374] <= 15'b011010000011110;
		Coeff[4375] <= 15'b011010000100001;
		Coeff[4376] <= 15'b011010000100100;
		Coeff[4377] <= 15'b011010000100111;
		Coeff[4378] <= 15'b011010000101010;
		Coeff[4379] <= 15'b011010000101100;
		Coeff[4380] <= 15'b011010000101111;
		Coeff[4381] <= 15'b011010000110010;
		Coeff[4382] <= 15'b011010000110101;
		Coeff[4383] <= 15'b011010000111000;
		Coeff[4384] <= 15'b011010000111011;
		Coeff[4385] <= 15'b011010000111110;
		Coeff[4386] <= 15'b011010001000001;
		Coeff[4387] <= 15'b011010001000011;
		Coeff[4388] <= 15'b011010001000110;
		Coeff[4389] <= 15'b011010001001001;
		Coeff[4390] <= 15'b011010001001100;
		Coeff[4391] <= 15'b011010001001111;
		Coeff[4392] <= 15'b011010001010010;
		Coeff[4393] <= 15'b011010001010101;
		Coeff[4394] <= 15'b011010001010111;
		Coeff[4395] <= 15'b011010001011010;
		Coeff[4396] <= 15'b011010001011101;
		Coeff[4397] <= 15'b011010001100000;
		Coeff[4398] <= 15'b011010001100011;
		Coeff[4399] <= 15'b011010001100110;
		Coeff[4400] <= 15'b011010001101001;
		Coeff[4401] <= 15'b011010001101100;
		Coeff[4402] <= 15'b011010001101110;
		Coeff[4403] <= 15'b011010001110001;
		Coeff[4404] <= 15'b011010001110100;
		Coeff[4405] <= 15'b011010001110111;
		Coeff[4406] <= 15'b011010001111010;
		Coeff[4407] <= 15'b011010001111101;
		Coeff[4408] <= 15'b011010010000000;
		Coeff[4409] <= 15'b011010010000010;
		Coeff[4410] <= 15'b011010010000101;
		Coeff[4411] <= 15'b011010010001000;
		Coeff[4412] <= 15'b011010010001011;
		Coeff[4413] <= 15'b011010010001110;
		Coeff[4414] <= 15'b011010010010001;
		Coeff[4415] <= 15'b011010010010100;
		Coeff[4416] <= 15'b011010010010111;
		Coeff[4417] <= 15'b011010010011001;
		Coeff[4418] <= 15'b011010010011100;
		Coeff[4419] <= 15'b011010010011111;
		Coeff[4420] <= 15'b011010010100010;
		Coeff[4421] <= 15'b011010010100101;
		Coeff[4422] <= 15'b011010010101000;
		Coeff[4423] <= 15'b011010010101011;
		Coeff[4424] <= 15'b011010010101101;
		Coeff[4425] <= 15'b011010010110000;
		Coeff[4426] <= 15'b011010010110011;
		Coeff[4427] <= 15'b011010010110110;
		Coeff[4428] <= 15'b011010010111001;
		Coeff[4429] <= 15'b011010010111100;
		Coeff[4430] <= 15'b011010010111111;
		Coeff[4431] <= 15'b011010011000001;
		Coeff[4432] <= 15'b011010011000100;
		Coeff[4433] <= 15'b011010011000111;
		Coeff[4434] <= 15'b011010011001010;
		Coeff[4435] <= 15'b011010011001101;
		Coeff[4436] <= 15'b011010011010000;
		Coeff[4437] <= 15'b011010011010011;
		Coeff[4438] <= 15'b011010011010101;
		Coeff[4439] <= 15'b011010011011000;
		Coeff[4440] <= 15'b011010011011011;
		Coeff[4441] <= 15'b011010011011110;
		Coeff[4442] <= 15'b011010011100001;
		Coeff[4443] <= 15'b011010011100100;
		Coeff[4444] <= 15'b011010011100111;
		Coeff[4445] <= 15'b011010011101010;
		Coeff[4446] <= 15'b011010011101100;
		Coeff[4447] <= 15'b011010011101111;
		Coeff[4448] <= 15'b011010011110010;
		Coeff[4449] <= 15'b011010011110101;
		Coeff[4450] <= 15'b011010011111000;
		Coeff[4451] <= 15'b011010011111011;
		Coeff[4452] <= 15'b011010011111110;
		Coeff[4453] <= 15'b011010100000000;
		Coeff[4454] <= 15'b011010100000011;
		Coeff[4455] <= 15'b011010100000110;
		Coeff[4456] <= 15'b011010100001001;
		Coeff[4457] <= 15'b011010100001100;
		Coeff[4458] <= 15'b011010100001111;
		Coeff[4459] <= 15'b011010100010010;
		Coeff[4460] <= 15'b011010100010100;
		Coeff[4461] <= 15'b011010100010111;
		Coeff[4462] <= 15'b011010100011010;
		Coeff[4463] <= 15'b011010100011101;
		Coeff[4464] <= 15'b011010100100000;
		Coeff[4465] <= 15'b011010100100011;
		Coeff[4466] <= 15'b011010100100110;
		Coeff[4467] <= 15'b011010100101000;
		Coeff[4468] <= 15'b011010100101011;
		Coeff[4469] <= 15'b011010100101110;
		Coeff[4470] <= 15'b011010100110001;
		Coeff[4471] <= 15'b011010100110100;
		Coeff[4472] <= 15'b011010100110111;
		Coeff[4473] <= 15'b011010100111010;
		Coeff[4474] <= 15'b011010100111100;
		Coeff[4475] <= 15'b011010100111111;
		Coeff[4476] <= 15'b011010101000010;
		Coeff[4477] <= 15'b011010101000101;
		Coeff[4478] <= 15'b011010101001000;
		Coeff[4479] <= 15'b011010101001011;
		Coeff[4480] <= 15'b011010101001110;
		Coeff[4481] <= 15'b011010101010000;
		Coeff[4482] <= 15'b011010101010011;
		Coeff[4483] <= 15'b011010101010110;
		Coeff[4484] <= 15'b011010101011001;
		Coeff[4485] <= 15'b011010101011100;
		Coeff[4486] <= 15'b011010101011111;
		Coeff[4487] <= 15'b011010101100010;
		Coeff[4488] <= 15'b011010101100100;
		Coeff[4489] <= 15'b011010101100111;
		Coeff[4490] <= 15'b011010101101010;
		Coeff[4491] <= 15'b011010101101101;
		Coeff[4492] <= 15'b011010101110000;
		Coeff[4493] <= 15'b011010101110011;
		Coeff[4494] <= 15'b011010101110110;
		Coeff[4495] <= 15'b011010101111000;
		Coeff[4496] <= 15'b011010101111011;
		Coeff[4497] <= 15'b011010101111110;
		Coeff[4498] <= 15'b011010110000001;
		Coeff[4499] <= 15'b011010110000100;
		Coeff[4500] <= 15'b011010110000111;
		Coeff[4501] <= 15'b011010110001010;
		Coeff[4502] <= 15'b011010110001100;
		Coeff[4503] <= 15'b011010110001111;
		Coeff[4504] <= 15'b011010110010010;
		Coeff[4505] <= 15'b011010110010101;
		Coeff[4506] <= 15'b011010110011000;
		Coeff[4507] <= 15'b011010110011011;
		Coeff[4508] <= 15'b011010110011101;
		Coeff[4509] <= 15'b011010110100000;
		Coeff[4510] <= 15'b011010110100011;
		Coeff[4511] <= 15'b011010110100110;
		Coeff[4512] <= 15'b011010110101001;
		Coeff[4513] <= 15'b011010110101100;
		Coeff[4514] <= 15'b011010110101111;
		Coeff[4515] <= 15'b011010110110001;
		Coeff[4516] <= 15'b011010110110100;
		Coeff[4517] <= 15'b011010110110111;
		Coeff[4518] <= 15'b011010110111010;
		Coeff[4519] <= 15'b011010110111101;
		Coeff[4520] <= 15'b011010111000000;
		Coeff[4521] <= 15'b011010111000011;
		Coeff[4522] <= 15'b011010111000101;
		Coeff[4523] <= 15'b011010111001000;
		Coeff[4524] <= 15'b011010111001011;
		Coeff[4525] <= 15'b011010111001110;
		Coeff[4526] <= 15'b011010111010001;
		Coeff[4527] <= 15'b011010111010100;
		Coeff[4528] <= 15'b011010111010111;
		Coeff[4529] <= 15'b011010111011001;
		Coeff[4530] <= 15'b011010111011100;
		Coeff[4531] <= 15'b011010111011111;
		Coeff[4532] <= 15'b011010111100010;
		Coeff[4533] <= 15'b011010111100101;
		Coeff[4534] <= 15'b011010111101000;
		Coeff[4535] <= 15'b011010111101010;
		Coeff[4536] <= 15'b011010111101101;
		Coeff[4537] <= 15'b011010111110000;
		Coeff[4538] <= 15'b011010111110011;
		Coeff[4539] <= 15'b011010111110110;
		Coeff[4540] <= 15'b011010111111001;
		Coeff[4541] <= 15'b011010111111100;
		Coeff[4542] <= 15'b011010111111110;
		Coeff[4543] <= 15'b011011000000001;
		Coeff[4544] <= 15'b011011000000100;
		Coeff[4545] <= 15'b011011000000111;
		Coeff[4546] <= 15'b011011000001010;
		Coeff[4547] <= 15'b011011000001101;
		Coeff[4548] <= 15'b011011000001111;
		Coeff[4549] <= 15'b011011000010010;
		Coeff[4550] <= 15'b011011000010101;
		Coeff[4551] <= 15'b011011000011000;
		Coeff[4552] <= 15'b011011000011011;
		Coeff[4553] <= 15'b011011000011110;
		Coeff[4554] <= 15'b011011000100001;
		Coeff[4555] <= 15'b011011000100011;
		Coeff[4556] <= 15'b011011000100110;
		Coeff[4557] <= 15'b011011000101001;
		Coeff[4558] <= 15'b011011000101100;
		Coeff[4559] <= 15'b011011000101111;
		Coeff[4560] <= 15'b011011000110010;
		Coeff[4561] <= 15'b011011000110101;
		Coeff[4562] <= 15'b011011000110111;
		Coeff[4563] <= 15'b011011000111010;
		Coeff[4564] <= 15'b011011000111101;
		Coeff[4565] <= 15'b011011001000000;
		Coeff[4566] <= 15'b011011001000011;
		Coeff[4567] <= 15'b011011001000110;
		Coeff[4568] <= 15'b011011001001000;
		Coeff[4569] <= 15'b011011001001011;
		Coeff[4570] <= 15'b011011001001110;
		Coeff[4571] <= 15'b011011001010001;
		Coeff[4572] <= 15'b011011001010100;
		Coeff[4573] <= 15'b011011001010111;
		Coeff[4574] <= 15'b011011001011001;
		Coeff[4575] <= 15'b011011001011100;
		Coeff[4576] <= 15'b011011001011111;
		Coeff[4577] <= 15'b011011001100010;
		Coeff[4578] <= 15'b011011001100101;
		Coeff[4579] <= 15'b011011001101000;
		Coeff[4580] <= 15'b011011001101011;
		Coeff[4581] <= 15'b011011001101101;
		Coeff[4582] <= 15'b011011001110000;
		Coeff[4583] <= 15'b011011001110011;
		Coeff[4584] <= 15'b011011001110110;
		Coeff[4585] <= 15'b011011001111001;
		Coeff[4586] <= 15'b011011001111100;
		Coeff[4587] <= 15'b011011001111110;
		Coeff[4588] <= 15'b011011010000001;
		Coeff[4589] <= 15'b011011010000100;
		Coeff[4590] <= 15'b011011010000111;
		Coeff[4591] <= 15'b011011010001010;
		Coeff[4592] <= 15'b011011010001101;
		Coeff[4593] <= 15'b011011010010000;
		Coeff[4594] <= 15'b011011010010010;
		Coeff[4595] <= 15'b011011010010101;
		Coeff[4596] <= 15'b011011010011000;
		Coeff[4597] <= 15'b011011010011011;
		Coeff[4598] <= 15'b011011010011110;
		Coeff[4599] <= 15'b011011010100001;
		Coeff[4600] <= 15'b011011010100011;
		Coeff[4601] <= 15'b011011010100110;
		Coeff[4602] <= 15'b011011010101001;
		Coeff[4603] <= 15'b011011010101100;
		Coeff[4604] <= 15'b011011010101111;
		Coeff[4605] <= 15'b011011010110010;
		Coeff[4606] <= 15'b011011010110100;
		Coeff[4607] <= 15'b011011010110111;
		Coeff[4608] <= 15'b011011010111010;
		Coeff[4609] <= 15'b011011010111101;
		Coeff[4610] <= 15'b011011011000000;
		Coeff[4611] <= 15'b011011011000011;
		Coeff[4612] <= 15'b011011011000101;
		Coeff[4613] <= 15'b011011011001000;
		Coeff[4614] <= 15'b011011011001011;
		Coeff[4615] <= 15'b011011011001110;
		Coeff[4616] <= 15'b011011011010001;
		Coeff[4617] <= 15'b011011011010100;
		Coeff[4618] <= 15'b011011011010111;
		Coeff[4619] <= 15'b011011011011001;
		Coeff[4620] <= 15'b011011011011100;
		Coeff[4621] <= 15'b011011011011111;
		Coeff[4622] <= 15'b011011011100010;
		Coeff[4623] <= 15'b011011011100101;
		Coeff[4624] <= 15'b011011011101000;
		Coeff[4625] <= 15'b011011011101010;
		Coeff[4626] <= 15'b011011011101101;
		Coeff[4627] <= 15'b011011011110000;
		Coeff[4628] <= 15'b011011011110011;
		Coeff[4629] <= 15'b011011011110110;
		Coeff[4630] <= 15'b011011011111001;
		Coeff[4631] <= 15'b011011011111011;
		Coeff[4632] <= 15'b011011011111110;
		Coeff[4633] <= 15'b011011100000001;
		Coeff[4634] <= 15'b011011100000100;
		Coeff[4635] <= 15'b011011100000111;
		Coeff[4636] <= 15'b011011100001010;
		Coeff[4637] <= 15'b011011100001100;
		Coeff[4638] <= 15'b011011100001111;
		Coeff[4639] <= 15'b011011100010010;
		Coeff[4640] <= 15'b011011100010101;
		Coeff[4641] <= 15'b011011100011000;
		Coeff[4642] <= 15'b011011100011011;
		Coeff[4643] <= 15'b011011100011101;
		Coeff[4644] <= 15'b011011100100000;
		Coeff[4645] <= 15'b011011100100011;
		Coeff[4646] <= 15'b011011100100110;
		Coeff[4647] <= 15'b011011100101001;
		Coeff[4648] <= 15'b011011100101100;
		Coeff[4649] <= 15'b011011100101110;
		Coeff[4650] <= 15'b011011100110001;
		Coeff[4651] <= 15'b011011100110100;
		Coeff[4652] <= 15'b011011100110111;
		Coeff[4653] <= 15'b011011100111010;
		Coeff[4654] <= 15'b011011100111101;
		Coeff[4655] <= 15'b011011100111111;
		Coeff[4656] <= 15'b011011101000010;
		Coeff[4657] <= 15'b011011101000101;
		Coeff[4658] <= 15'b011011101001000;
		Coeff[4659] <= 15'b011011101001011;
		Coeff[4660] <= 15'b011011101001110;
		Coeff[4661] <= 15'b011011101010000;
		Coeff[4662] <= 15'b011011101010011;
		Coeff[4663] <= 15'b011011101010110;
		Coeff[4664] <= 15'b011011101011001;
		Coeff[4665] <= 15'b011011101011100;
		Coeff[4666] <= 15'b011011101011111;
		Coeff[4667] <= 15'b011011101100001;
		Coeff[4668] <= 15'b011011101100100;
		Coeff[4669] <= 15'b011011101100111;
		Coeff[4670] <= 15'b011011101101010;
		Coeff[4671] <= 15'b011011101101101;
		Coeff[4672] <= 15'b011011101110000;
		Coeff[4673] <= 15'b011011101110010;
		Coeff[4674] <= 15'b011011101110101;
		Coeff[4675] <= 15'b011011101111000;
		Coeff[4676] <= 15'b011011101111011;
		Coeff[4677] <= 15'b011011101111110;
		Coeff[4678] <= 15'b011011110000001;
		Coeff[4679] <= 15'b011011110000011;
		Coeff[4680] <= 15'b011011110000110;
		Coeff[4681] <= 15'b011011110001001;
		Coeff[4682] <= 15'b011011110001100;
		Coeff[4683] <= 15'b011011110001111;
		Coeff[4684] <= 15'b011011110010010;
		Coeff[4685] <= 15'b011011110010100;
		Coeff[4686] <= 15'b011011110010111;
		Coeff[4687] <= 15'b011011110011010;
		Coeff[4688] <= 15'b011011110011101;
		Coeff[4689] <= 15'b011011110100000;
		Coeff[4690] <= 15'b011011110100011;
		Coeff[4691] <= 15'b011011110100101;
		Coeff[4692] <= 15'b011011110101000;
		Coeff[4693] <= 15'b011011110101011;
		Coeff[4694] <= 15'b011011110101110;
		Coeff[4695] <= 15'b011011110110001;
		Coeff[4696] <= 15'b011011110110100;
		Coeff[4697] <= 15'b011011110110110;
		Coeff[4698] <= 15'b011011110111001;
		Coeff[4699] <= 15'b011011110111100;
		Coeff[4700] <= 15'b011011110111111;
		Coeff[4701] <= 15'b011011111000010;
		Coeff[4702] <= 15'b011011111000101;
		Coeff[4703] <= 15'b011011111000111;
		Coeff[4704] <= 15'b011011111001010;
		Coeff[4705] <= 15'b011011111001101;
		Coeff[4706] <= 15'b011011111010000;
		Coeff[4707] <= 15'b011011111010011;
		Coeff[4708] <= 15'b011011111010101;
		Coeff[4709] <= 15'b011011111011000;
		Coeff[4710] <= 15'b011011111011011;
		Coeff[4711] <= 15'b011011111011110;
		Coeff[4712] <= 15'b011011111100001;
		Coeff[4713] <= 15'b011011111100100;
		Coeff[4714] <= 15'b011011111100110;
		Coeff[4715] <= 15'b011011111101001;
		Coeff[4716] <= 15'b011011111101100;
		Coeff[4717] <= 15'b011011111101111;
		Coeff[4718] <= 15'b011011111110010;
		Coeff[4719] <= 15'b011011111110101;
		Coeff[4720] <= 15'b011011111110111;
		Coeff[4721] <= 15'b011011111111010;
		Coeff[4722] <= 15'b011011111111101;
		Coeff[4723] <= 15'b011100000000000;
		Coeff[4724] <= 15'b011100000000011;
		Coeff[4725] <= 15'b011100000000110;
		Coeff[4726] <= 15'b011100000001000;
		Coeff[4727] <= 15'b011100000001011;
		Coeff[4728] <= 15'b011100000001110;
		Coeff[4729] <= 15'b011100000010001;
		Coeff[4730] <= 15'b011100000010100;
		Coeff[4731] <= 15'b011100000010110;
		Coeff[4732] <= 15'b011100000011001;
		Coeff[4733] <= 15'b011100000011100;
		Coeff[4734] <= 15'b011100000011111;
		Coeff[4735] <= 15'b011100000100010;
		Coeff[4736] <= 15'b011100000100101;
		Coeff[4737] <= 15'b011100000100111;
		Coeff[4738] <= 15'b011100000101010;
		Coeff[4739] <= 15'b011100000101101;
		Coeff[4740] <= 15'b011100000110000;
		Coeff[4741] <= 15'b011100000110011;
		Coeff[4742] <= 15'b011100000110110;
		Coeff[4743] <= 15'b011100000111000;
		Coeff[4744] <= 15'b011100000111011;
		Coeff[4745] <= 15'b011100000111110;
		Coeff[4746] <= 15'b011100001000001;
		Coeff[4747] <= 15'b011100001000100;
		Coeff[4748] <= 15'b011100001000110;
		Coeff[4749] <= 15'b011100001001001;
		Coeff[4750] <= 15'b011100001001100;
		Coeff[4751] <= 15'b011100001001111;
		Coeff[4752] <= 15'b011100001010010;
		Coeff[4753] <= 15'b011100001010101;
		Coeff[4754] <= 15'b011100001010111;
		Coeff[4755] <= 15'b011100001011010;
		Coeff[4756] <= 15'b011100001011101;
		Coeff[4757] <= 15'b011100001100000;
		Coeff[4758] <= 15'b011100001100011;
		Coeff[4759] <= 15'b011100001100101;
		Coeff[4760] <= 15'b011100001101000;
		Coeff[4761] <= 15'b011100001101011;
		Coeff[4762] <= 15'b011100001101110;
		Coeff[4763] <= 15'b011100001110001;
		Coeff[4764] <= 15'b011100001110100;
		Coeff[4765] <= 15'b011100001110110;
		Coeff[4766] <= 15'b011100001111001;
		Coeff[4767] <= 15'b011100001111100;
		Coeff[4768] <= 15'b011100001111111;
		Coeff[4769] <= 15'b011100010000010;
		Coeff[4770] <= 15'b011100010000100;
		Coeff[4771] <= 15'b011100010000111;
		Coeff[4772] <= 15'b011100010001010;
		Coeff[4773] <= 15'b011100010001101;
		Coeff[4774] <= 15'b011100010010000;
		Coeff[4775] <= 15'b011100010010011;
		Coeff[4776] <= 15'b011100010010101;
		Coeff[4777] <= 15'b011100010011000;
		Coeff[4778] <= 15'b011100010011011;
		Coeff[4779] <= 15'b011100010011110;
		Coeff[4780] <= 15'b011100010100001;
		Coeff[4781] <= 15'b011100010100011;
		Coeff[4782] <= 15'b011100010100110;
		Coeff[4783] <= 15'b011100010101001;
		Coeff[4784] <= 15'b011100010101100;
		Coeff[4785] <= 15'b011100010101111;
		Coeff[4786] <= 15'b011100010110010;
		Coeff[4787] <= 15'b011100010110100;
		Coeff[4788] <= 15'b011100010110111;
		Coeff[4789] <= 15'b011100010111010;
		Coeff[4790] <= 15'b011100010111101;
		Coeff[4791] <= 15'b011100011000000;
		Coeff[4792] <= 15'b011100011000010;
		Coeff[4793] <= 15'b011100011000101;
		Coeff[4794] <= 15'b011100011001000;
		Coeff[4795] <= 15'b011100011001011;
		Coeff[4796] <= 15'b011100011001110;
		Coeff[4797] <= 15'b011100011010001;
		Coeff[4798] <= 15'b011100011010011;
		Coeff[4799] <= 15'b011100011010110;
		Coeff[4800] <= 15'b011100011011001;
		Coeff[4801] <= 15'b011100011011100;
		Coeff[4802] <= 15'b011100011011111;
		Coeff[4803] <= 15'b011100011100001;
		Coeff[4804] <= 15'b011100011100100;
		Coeff[4805] <= 15'b011100011100111;
		Coeff[4806] <= 15'b011100011101010;
		Coeff[4807] <= 15'b011100011101101;
		Coeff[4808] <= 15'b011100011110000;
		Coeff[4809] <= 15'b011100011110010;
		Coeff[4810] <= 15'b011100011110101;
		Coeff[4811] <= 15'b011100011111000;
		Coeff[4812] <= 15'b011100011111011;
		Coeff[4813] <= 15'b011100011111110;
		Coeff[4814] <= 15'b011100100000000;
		Coeff[4815] <= 15'b011100100000011;
		Coeff[4816] <= 15'b011100100000110;
		Coeff[4817] <= 15'b011100100001001;
		Coeff[4818] <= 15'b011100100001100;
		Coeff[4819] <= 15'b011100100001110;
		Coeff[4820] <= 15'b011100100010001;
		Coeff[4821] <= 15'b011100100010100;
		Coeff[4822] <= 15'b011100100010111;
		Coeff[4823] <= 15'b011100100011010;
		Coeff[4824] <= 15'b011100100011101;
		Coeff[4825] <= 15'b011100100011111;
		Coeff[4826] <= 15'b011100100100010;
		Coeff[4827] <= 15'b011100100100101;
		Coeff[4828] <= 15'b011100100101000;
		Coeff[4829] <= 15'b011100100101011;
		Coeff[4830] <= 15'b011100100101101;
		Coeff[4831] <= 15'b011100100110000;
		Coeff[4832] <= 15'b011100100110011;
		Coeff[4833] <= 15'b011100100110110;
		Coeff[4834] <= 15'b011100100111001;
		Coeff[4835] <= 15'b011100100111011;
		Coeff[4836] <= 15'b011100100111110;
		Coeff[4837] <= 15'b011100101000001;
		Coeff[4838] <= 15'b011100101000100;
		Coeff[4839] <= 15'b011100101000111;
		Coeff[4840] <= 15'b011100101001001;
		Coeff[4841] <= 15'b011100101001100;
		Coeff[4842] <= 15'b011100101001111;
		Coeff[4843] <= 15'b011100101010010;
		Coeff[4844] <= 15'b011100101010101;
		Coeff[4845] <= 15'b011100101011000;
		Coeff[4846] <= 15'b011100101011010;
		Coeff[4847] <= 15'b011100101011101;
		Coeff[4848] <= 15'b011100101100000;
		Coeff[4849] <= 15'b011100101100011;
		Coeff[4850] <= 15'b011100101100110;
		Coeff[4851] <= 15'b011100101101000;
		Coeff[4852] <= 15'b011100101101011;
		Coeff[4853] <= 15'b011100101101110;
		Coeff[4854] <= 15'b011100101110001;
		Coeff[4855] <= 15'b011100101110100;
		Coeff[4856] <= 15'b011100101110110;
		Coeff[4857] <= 15'b011100101111001;
		Coeff[4858] <= 15'b011100101111100;
		Coeff[4859] <= 15'b011100101111111;
		Coeff[4860] <= 15'b011100110000010;
		Coeff[4861] <= 15'b011100110000100;
		Coeff[4862] <= 15'b011100110000111;
		Coeff[4863] <= 15'b011100110001010;
		Coeff[4864] <= 15'b011100110001101;
		Coeff[4865] <= 15'b011100110010000;
		Coeff[4866] <= 15'b011100110010010;
		Coeff[4867] <= 15'b011100110010101;
		Coeff[4868] <= 15'b011100110011000;
		Coeff[4869] <= 15'b011100110011011;
		Coeff[4870] <= 15'b011100110011110;
		Coeff[4871] <= 15'b011100110100001;
		Coeff[4872] <= 15'b011100110100011;
		Coeff[4873] <= 15'b011100110100110;
		Coeff[4874] <= 15'b011100110101001;
		Coeff[4875] <= 15'b011100110101100;
		Coeff[4876] <= 15'b011100110101111;
		Coeff[4877] <= 15'b011100110110001;
		Coeff[4878] <= 15'b011100110110100;
		Coeff[4879] <= 15'b011100110110111;
		Coeff[4880] <= 15'b011100110111010;
		Coeff[4881] <= 15'b011100110111101;
		Coeff[4882] <= 15'b011100110111111;
		Coeff[4883] <= 15'b011100111000010;
		Coeff[4884] <= 15'b011100111000101;
		Coeff[4885] <= 15'b011100111001000;
		Coeff[4886] <= 15'b011100111001011;
		Coeff[4887] <= 15'b011100111001101;
		Coeff[4888] <= 15'b011100111010000;
		Coeff[4889] <= 15'b011100111010011;
		Coeff[4890] <= 15'b011100111010110;
		Coeff[4891] <= 15'b011100111011001;
		Coeff[4892] <= 15'b011100111011011;
		Coeff[4893] <= 15'b011100111011110;
		Coeff[4894] <= 15'b011100111100001;
		Coeff[4895] <= 15'b011100111100100;
		Coeff[4896] <= 15'b011100111100111;
		Coeff[4897] <= 15'b011100111101001;
		Coeff[4898] <= 15'b011100111101100;
		Coeff[4899] <= 15'b011100111101111;
		Coeff[4900] <= 15'b011100111110010;
		Coeff[4901] <= 15'b011100111110101;
		Coeff[4902] <= 15'b011100111110111;
		Coeff[4903] <= 15'b011100111111010;
		Coeff[4904] <= 15'b011100111111101;
		Coeff[4905] <= 15'b011101000000000;
		Coeff[4906] <= 15'b011101000000011;
		Coeff[4907] <= 15'b011101000000101;
		Coeff[4908] <= 15'b011101000001000;
		Coeff[4909] <= 15'b011101000001011;
		Coeff[4910] <= 15'b011101000001110;
		Coeff[4911] <= 15'b011101000010001;
		Coeff[4912] <= 15'b011101000010011;
		Coeff[4913] <= 15'b011101000010110;
		Coeff[4914] <= 15'b011101000011001;
		Coeff[4915] <= 15'b011101000011100;
		Coeff[4916] <= 15'b011101000011111;
		Coeff[4917] <= 15'b011101000100001;
		Coeff[4918] <= 15'b011101000100100;
		Coeff[4919] <= 15'b011101000100111;
		Coeff[4920] <= 15'b011101000101010;
		Coeff[4921] <= 15'b011101000101101;
		Coeff[4922] <= 15'b011101000101111;
		Coeff[4923] <= 15'b011101000110010;
		Coeff[4924] <= 15'b011101000110101;
		Coeff[4925] <= 15'b011101000111000;
		Coeff[4926] <= 15'b011101000111011;
		Coeff[4927] <= 15'b011101000111101;
		Coeff[4928] <= 15'b011101001000000;
		Coeff[4929] <= 15'b011101001000011;
		Coeff[4930] <= 15'b011101001000110;
		Coeff[4931] <= 15'b011101001001001;
		Coeff[4932] <= 15'b011101001001011;
		Coeff[4933] <= 15'b011101001001110;
		Coeff[4934] <= 15'b011101001010001;
		Coeff[4935] <= 15'b011101001010100;
		Coeff[4936] <= 15'b011101001010111;
		Coeff[4937] <= 15'b011101001011001;
		Coeff[4938] <= 15'b011101001011100;
		Coeff[4939] <= 15'b011101001011111;
		Coeff[4940] <= 15'b011101001100010;
		Coeff[4941] <= 15'b011101001100101;
		Coeff[4942] <= 15'b011101001100111;
		Coeff[4943] <= 15'b011101001101010;
		Coeff[4944] <= 15'b011101001101101;
		Coeff[4945] <= 15'b011101001110000;
		Coeff[4946] <= 15'b011101001110011;
		Coeff[4947] <= 15'b011101001110101;
		Coeff[4948] <= 15'b011101001111000;
		Coeff[4949] <= 15'b011101001111011;
		Coeff[4950] <= 15'b011101001111110;
		Coeff[4951] <= 15'b011101010000000;
		Coeff[4952] <= 15'b011101010000011;
		Coeff[4953] <= 15'b011101010000110;
		Coeff[4954] <= 15'b011101010001001;
		Coeff[4955] <= 15'b011101010001100;
		Coeff[4956] <= 15'b011101010001110;
		Coeff[4957] <= 15'b011101010010001;
		Coeff[4958] <= 15'b011101010010100;
		Coeff[4959] <= 15'b011101010010111;
		Coeff[4960] <= 15'b011101010011010;
		Coeff[4961] <= 15'b011101010011100;
		Coeff[4962] <= 15'b011101010011111;
		Coeff[4963] <= 15'b011101010100010;
		Coeff[4964] <= 15'b011101010100101;
		Coeff[4965] <= 15'b011101010101000;
		Coeff[4966] <= 15'b011101010101010;
		Coeff[4967] <= 15'b011101010101101;
		Coeff[4968] <= 15'b011101010110000;
		Coeff[4969] <= 15'b011101010110011;
		Coeff[4970] <= 15'b011101010110110;
		Coeff[4971] <= 15'b011101010111000;
		Coeff[4972] <= 15'b011101010111011;
		Coeff[4973] <= 15'b011101010111110;
		Coeff[4974] <= 15'b011101011000001;
		Coeff[4975] <= 15'b011101011000100;
		Coeff[4976] <= 15'b011101011000110;
		Coeff[4977] <= 15'b011101011001001;
		Coeff[4978] <= 15'b011101011001100;
		Coeff[4979] <= 15'b011101011001111;
		Coeff[4980] <= 15'b011101011010001;
		Coeff[4981] <= 15'b011101011010100;
		Coeff[4982] <= 15'b011101011010111;
		Coeff[4983] <= 15'b011101011011010;
		Coeff[4984] <= 15'b011101011011101;
		Coeff[4985] <= 15'b011101011011111;
		Coeff[4986] <= 15'b011101011100010;
		Coeff[4987] <= 15'b011101011100101;
		Coeff[4988] <= 15'b011101011101000;
		Coeff[4989] <= 15'b011101011101011;
		Coeff[4990] <= 15'b011101011101101;
		Coeff[4991] <= 15'b011101011110000;
		Coeff[4992] <= 15'b011101011110011;
		Coeff[4993] <= 15'b011101011110110;
		Coeff[4994] <= 15'b011101011111001;
		Coeff[4995] <= 15'b011101011111011;
		Coeff[4996] <= 15'b011101011111110;
		Coeff[4997] <= 15'b011101100000001;
		Coeff[4998] <= 15'b011101100000100;
		Coeff[4999] <= 15'b011101100000110;
		Coeff[5000] <= 15'b011101100001001;
		Coeff[5001] <= 15'b011101100001100;
		Coeff[5002] <= 15'b011101100001111;
		Coeff[5003] <= 15'b011101100010010;
		Coeff[5004] <= 15'b011101100010100;
		Coeff[5005] <= 15'b011101100010111;
		Coeff[5006] <= 15'b011101100011010;
		Coeff[5007] <= 15'b011101100011101;
		Coeff[5008] <= 15'b011101100100000;
		Coeff[5009] <= 15'b011101100100010;
		Coeff[5010] <= 15'b011101100100101;
		Coeff[5011] <= 15'b011101100101000;
		Coeff[5012] <= 15'b011101100101011;
		Coeff[5013] <= 15'b011101100101101;
		Coeff[5014] <= 15'b011101100110000;
		Coeff[5015] <= 15'b011101100110011;
		Coeff[5016] <= 15'b011101100110110;
		Coeff[5017] <= 15'b011101100111001;
		Coeff[5018] <= 15'b011101100111011;
		Coeff[5019] <= 15'b011101100111110;
		Coeff[5020] <= 15'b011101101000001;
		Coeff[5021] <= 15'b011101101000100;
		Coeff[5022] <= 15'b011101101000111;
		Coeff[5023] <= 15'b011101101001001;
		Coeff[5024] <= 15'b011101101001100;
		Coeff[5025] <= 15'b011101101001111;
		Coeff[5026] <= 15'b011101101010010;
		Coeff[5027] <= 15'b011101101010100;
		Coeff[5028] <= 15'b011101101010111;
		Coeff[5029] <= 15'b011101101011010;
		Coeff[5030] <= 15'b011101101011101;
		Coeff[5031] <= 15'b011101101100000;
		Coeff[5032] <= 15'b011101101100010;
		Coeff[5033] <= 15'b011101101100101;
		Coeff[5034] <= 15'b011101101101000;
		Coeff[5035] <= 15'b011101101101011;
		Coeff[5036] <= 15'b011101101101101;
		Coeff[5037] <= 15'b011101101110000;
		Coeff[5038] <= 15'b011101101110011;
		Coeff[5039] <= 15'b011101101110110;
		Coeff[5040] <= 15'b011101101111001;
		Coeff[5041] <= 15'b011101101111011;
		Coeff[5042] <= 15'b011101101111110;
		Coeff[5043] <= 15'b011101110000001;
		Coeff[5044] <= 15'b011101110000100;
		Coeff[5045] <= 15'b011101110000111;
		Coeff[5046] <= 15'b011101110001001;
		Coeff[5047] <= 15'b011101110001100;
		Coeff[5048] <= 15'b011101110001111;
		Coeff[5049] <= 15'b011101110010010;
		Coeff[5050] <= 15'b011101110010100;
		Coeff[5051] <= 15'b011101110010111;
		Coeff[5052] <= 15'b011101110011010;
		Coeff[5053] <= 15'b011101110011101;
		Coeff[5054] <= 15'b011101110100000;
		Coeff[5055] <= 15'b011101110100010;
		Coeff[5056] <= 15'b011101110100101;
		Coeff[5057] <= 15'b011101110101000;
		Coeff[5058] <= 15'b011101110101011;
		Coeff[5059] <= 15'b011101110101101;
		Coeff[5060] <= 15'b011101110110000;
		Coeff[5061] <= 15'b011101110110011;
		Coeff[5062] <= 15'b011101110110110;
		Coeff[5063] <= 15'b011101110111001;
		Coeff[5064] <= 15'b011101110111011;
		Coeff[5065] <= 15'b011101110111110;
		Coeff[5066] <= 15'b011101111000001;
		Coeff[5067] <= 15'b011101111000100;
		Coeff[5068] <= 15'b011101111000110;
		Coeff[5069] <= 15'b011101111001001;
		Coeff[5070] <= 15'b011101111001100;
		Coeff[5071] <= 15'b011101111001111;
		Coeff[5072] <= 15'b011101111010010;
		Coeff[5073] <= 15'b011101111010100;
		Coeff[5074] <= 15'b011101111010111;
		Coeff[5075] <= 15'b011101111011010;
		Coeff[5076] <= 15'b011101111011101;
		Coeff[5077] <= 15'b011101111011111;
		Coeff[5078] <= 15'b011101111100010;
		Coeff[5079] <= 15'b011101111100101;
		Coeff[5080] <= 15'b011101111101000;
		Coeff[5081] <= 15'b011101111101011;
		Coeff[5082] <= 15'b011101111101101;
		Coeff[5083] <= 15'b011101111110000;
		Coeff[5084] <= 15'b011101111110011;
		Coeff[5085] <= 15'b011101111110110;
		Coeff[5086] <= 15'b011101111111000;
		Coeff[5087] <= 15'b011101111111011;
		Coeff[5088] <= 15'b011101111111110;
		Coeff[5089] <= 15'b011110000000001;
		Coeff[5090] <= 15'b011110000000100;
		Coeff[5091] <= 15'b011110000000110;
		Coeff[5092] <= 15'b011110000001001;
		Coeff[5093] <= 15'b011110000001100;
		Coeff[5094] <= 15'b011110000001111;
		Coeff[5095] <= 15'b011110000010001;
		Coeff[5096] <= 15'b011110000010100;
		Coeff[5097] <= 15'b011110000010111;
		Coeff[5098] <= 15'b011110000011010;
		Coeff[5099] <= 15'b011110000011101;
		Coeff[5100] <= 15'b011110000011111;
		Coeff[5101] <= 15'b011110000100010;
		Coeff[5102] <= 15'b011110000100101;
		Coeff[5103] <= 15'b011110000101000;
		Coeff[5104] <= 15'b011110000101010;
		Coeff[5105] <= 15'b011110000101101;
		Coeff[5106] <= 15'b011110000110000;
		Coeff[5107] <= 15'b011110000110011;
		Coeff[5108] <= 15'b011110000110101;
		Coeff[5109] <= 15'b011110000111000;
		Coeff[5110] <= 15'b011110000111011;
		Coeff[5111] <= 15'b011110000111110;
		Coeff[5112] <= 15'b011110001000001;
		Coeff[5113] <= 15'b011110001000011;
		Coeff[5114] <= 15'b011110001000110;
		Coeff[5115] <= 15'b011110001001001;
		Coeff[5116] <= 15'b011110001001100;
		Coeff[5117] <= 15'b011110001001110;
		Coeff[5118] <= 15'b011110001010001;
		Coeff[5119] <= 15'b011110001010100;
		Coeff[5120] <= 15'b011110001010111;
		Coeff[5121] <= 15'b011110001011001;
		Coeff[5122] <= 15'b011110001011100;
		Coeff[5123] <= 15'b011110001011111;
		Coeff[5124] <= 15'b011110001100010;
		Coeff[5125] <= 15'b011110001100101;
		Coeff[5126] <= 15'b011110001100111;
		Coeff[5127] <= 15'b011110001101010;
		Coeff[5128] <= 15'b011110001101101;
		Coeff[5129] <= 15'b011110001110000;
		Coeff[5130] <= 15'b011110001110010;
		Coeff[5131] <= 15'b011110001110101;
		Coeff[5132] <= 15'b011110001111000;
		Coeff[5133] <= 15'b011110001111011;
		Coeff[5134] <= 15'b011110001111110;
		Coeff[5135] <= 15'b011110010000000;
		Coeff[5136] <= 15'b011110010000011;
		Coeff[5137] <= 15'b011110010000110;
		Coeff[5138] <= 15'b011110010001001;
		Coeff[5139] <= 15'b011110010001011;
		Coeff[5140] <= 15'b011110010001110;
		Coeff[5141] <= 15'b011110010010001;
		Coeff[5142] <= 15'b011110010010100;
		Coeff[5143] <= 15'b011110010010110;
		Coeff[5144] <= 15'b011110010011001;
		Coeff[5145] <= 15'b011110010011100;
		Coeff[5146] <= 15'b011110010011111;
		Coeff[5147] <= 15'b011110010100001;
		Coeff[5148] <= 15'b011110010100100;
		Coeff[5149] <= 15'b011110010100111;
		Coeff[5150] <= 15'b011110010101010;
		Coeff[5151] <= 15'b011110010101101;
		Coeff[5152] <= 15'b011110010101111;
		Coeff[5153] <= 15'b011110010110010;
		Coeff[5154] <= 15'b011110010110101;
		Coeff[5155] <= 15'b011110010111000;
		Coeff[5156] <= 15'b011110010111010;
		Coeff[5157] <= 15'b011110010111101;
		Coeff[5158] <= 15'b011110011000000;
		Coeff[5159] <= 15'b011110011000011;
		Coeff[5160] <= 15'b011110011000101;
		Coeff[5161] <= 15'b011110011001000;
		Coeff[5162] <= 15'b011110011001011;
		Coeff[5163] <= 15'b011110011001110;
		Coeff[5164] <= 15'b011110011010000;
		Coeff[5165] <= 15'b011110011010011;
		Coeff[5166] <= 15'b011110011010110;
		Coeff[5167] <= 15'b011110011011001;
		Coeff[5168] <= 15'b011110011011100;
		Coeff[5169] <= 15'b011110011011110;
		Coeff[5170] <= 15'b011110011100001;
		Coeff[5171] <= 15'b011110011100100;
		Coeff[5172] <= 15'b011110011100111;
		Coeff[5173] <= 15'b011110011101001;
		Coeff[5174] <= 15'b011110011101100;
		Coeff[5175] <= 15'b011110011101111;
		Coeff[5176] <= 15'b011110011110010;
		Coeff[5177] <= 15'b011110011110100;
		Coeff[5178] <= 15'b011110011110111;
		Coeff[5179] <= 15'b011110011111010;
		Coeff[5180] <= 15'b011110011111101;
		Coeff[5181] <= 15'b011110011111111;
		Coeff[5182] <= 15'b011110100000010;
		Coeff[5183] <= 15'b011110100000101;
		Coeff[5184] <= 15'b011110100001000;
		Coeff[5185] <= 15'b011110100001011;
		Coeff[5186] <= 15'b011110100001101;
		Coeff[5187] <= 15'b011110100010000;
		Coeff[5188] <= 15'b011110100010011;
		Coeff[5189] <= 15'b011110100010110;
		Coeff[5190] <= 15'b011110100011000;
		Coeff[5191] <= 15'b011110100011011;
		Coeff[5192] <= 15'b011110100011110;
		Coeff[5193] <= 15'b011110100100001;
		Coeff[5194] <= 15'b011110100100011;
		Coeff[5195] <= 15'b011110100100110;
		Coeff[5196] <= 15'b011110100101001;
		Coeff[5197] <= 15'b011110100101100;
		Coeff[5198] <= 15'b011110100101110;
		Coeff[5199] <= 15'b011110100110001;
		Coeff[5200] <= 15'b011110100110100;
		Coeff[5201] <= 15'b011110100110111;
		Coeff[5202] <= 15'b011110100111001;
		Coeff[5203] <= 15'b011110100111100;
		Coeff[5204] <= 15'b011110100111111;
		Coeff[5205] <= 15'b011110101000010;
		Coeff[5206] <= 15'b011110101000100;
		Coeff[5207] <= 15'b011110101000111;
		Coeff[5208] <= 15'b011110101001010;
		Coeff[5209] <= 15'b011110101001101;
		Coeff[5210] <= 15'b011110101010000;
		Coeff[5211] <= 15'b011110101010010;
		Coeff[5212] <= 15'b011110101010101;
		Coeff[5213] <= 15'b011110101011000;
		Coeff[5214] <= 15'b011110101011011;
		Coeff[5215] <= 15'b011110101011101;
		Coeff[5216] <= 15'b011110101100000;
		Coeff[5217] <= 15'b011110101100011;
		Coeff[5218] <= 15'b011110101100110;
		Coeff[5219] <= 15'b011110101101000;
		Coeff[5220] <= 15'b011110101101011;
		Coeff[5221] <= 15'b011110101101110;
		Coeff[5222] <= 15'b011110101110001;
		Coeff[5223] <= 15'b011110101110011;
		Coeff[5224] <= 15'b011110101110110;
		Coeff[5225] <= 15'b011110101111001;
		Coeff[5226] <= 15'b011110101111100;
		Coeff[5227] <= 15'b011110101111110;
		Coeff[5228] <= 15'b011110110000001;
		Coeff[5229] <= 15'b011110110000100;
		Coeff[5230] <= 15'b011110110000111;
		Coeff[5231] <= 15'b011110110001001;
		Coeff[5232] <= 15'b011110110001100;
		Coeff[5233] <= 15'b011110110001111;
		Coeff[5234] <= 15'b011110110010010;
		Coeff[5235] <= 15'b011110110010100;
		Coeff[5236] <= 15'b011110110010111;
		Coeff[5237] <= 15'b011110110011010;
		Coeff[5238] <= 15'b011110110011101;
		Coeff[5239] <= 15'b011110110011111;
		Coeff[5240] <= 15'b011110110100010;
		Coeff[5241] <= 15'b011110110100101;
		Coeff[5242] <= 15'b011110110101000;
		Coeff[5243] <= 15'b011110110101010;
		Coeff[5244] <= 15'b011110110101101;
		Coeff[5245] <= 15'b011110110110000;
		Coeff[5246] <= 15'b011110110110011;
		Coeff[5247] <= 15'b011110110110101;
		Coeff[5248] <= 15'b011110110111000;
		Coeff[5249] <= 15'b011110110111011;
		Coeff[5250] <= 15'b011110110111110;
		Coeff[5251] <= 15'b011110111000000;
		Coeff[5252] <= 15'b011110111000011;
		Coeff[5253] <= 15'b011110111000110;
		Coeff[5254] <= 15'b011110111001001;
		Coeff[5255] <= 15'b011110111001011;
		Coeff[5256] <= 15'b011110111001110;
		Coeff[5257] <= 15'b011110111010001;
		Coeff[5258] <= 15'b011110111010100;
		Coeff[5259] <= 15'b011110111010110;
		Coeff[5260] <= 15'b011110111011001;
		Coeff[5261] <= 15'b011110111011100;
		Coeff[5262] <= 15'b011110111011111;
		Coeff[5263] <= 15'b011110111100001;
		Coeff[5264] <= 15'b011110111100100;
		Coeff[5265] <= 15'b011110111100111;
		Coeff[5266] <= 15'b011110111101010;
		Coeff[5267] <= 15'b011110111101100;
		Coeff[5268] <= 15'b011110111101111;
		Coeff[5269] <= 15'b011110111110010;
		Coeff[5270] <= 15'b011110111110101;
		Coeff[5271] <= 15'b011110111110111;
		Coeff[5272] <= 15'b011110111111010;
		Coeff[5273] <= 15'b011110111111101;
		Coeff[5274] <= 15'b011111000000000;
		Coeff[5275] <= 15'b011111000000010;
		Coeff[5276] <= 15'b011111000000101;
		Coeff[5277] <= 15'b011111000001000;
		Coeff[5278] <= 15'b011111000001011;
		Coeff[5279] <= 15'b011111000001101;
		Coeff[5280] <= 15'b011111000010000;
		Coeff[5281] <= 15'b011111000010011;
		Coeff[5282] <= 15'b011111000010110;
		Coeff[5283] <= 15'b011111000011000;
		Coeff[5284] <= 15'b011111000011011;
		Coeff[5285] <= 15'b011111000011110;
		Coeff[5286] <= 15'b011111000100001;
		Coeff[5287] <= 15'b011111000100011;
		Coeff[5288] <= 15'b011111000100110;
		Coeff[5289] <= 15'b011111000101001;
		Coeff[5290] <= 15'b011111000101100;
		Coeff[5291] <= 15'b011111000101110;
		Coeff[5292] <= 15'b011111000110001;
		Coeff[5293] <= 15'b011111000110100;
		Coeff[5294] <= 15'b011111000110111;
		Coeff[5295] <= 15'b011111000111001;
		Coeff[5296] <= 15'b011111000111100;
		Coeff[5297] <= 15'b011111000111111;
		Coeff[5298] <= 15'b011111001000010;
		Coeff[5299] <= 15'b011111001000100;
		Coeff[5300] <= 15'b011111001000111;
		Coeff[5301] <= 15'b011111001001010;
		Coeff[5302] <= 15'b011111001001101;
		Coeff[5303] <= 15'b011111001001111;
		Coeff[5304] <= 15'b011111001010010;
		Coeff[5305] <= 15'b011111001010101;
		Coeff[5306] <= 15'b011111001011000;
		Coeff[5307] <= 15'b011111001011010;
		Coeff[5308] <= 15'b011111001011101;
		Coeff[5309] <= 15'b011111001100000;
		Coeff[5310] <= 15'b011111001100011;
		Coeff[5311] <= 15'b011111001100101;
		Coeff[5312] <= 15'b011111001101000;
		Coeff[5313] <= 15'b011111001101011;
		Coeff[5314] <= 15'b011111001101110;
		Coeff[5315] <= 15'b011111001110000;
		Coeff[5316] <= 15'b011111001110011;
		Coeff[5317] <= 15'b011111001110110;
		Coeff[5318] <= 15'b011111001111000;
		Coeff[5319] <= 15'b011111001111011;
		Coeff[5320] <= 15'b011111001111110;
		Coeff[5321] <= 15'b011111010000001;
		Coeff[5322] <= 15'b011111010000011;
		Coeff[5323] <= 15'b011111010000110;
		Coeff[5324] <= 15'b011111010001001;
		Coeff[5325] <= 15'b011111010001100;
		Coeff[5326] <= 15'b011111010001110;
		Coeff[5327] <= 15'b011111010010001;
		Coeff[5328] <= 15'b011111010010100;
		Coeff[5329] <= 15'b011111010010111;
		Coeff[5330] <= 15'b011111010011001;
		Coeff[5331] <= 15'b011111010011100;
		Coeff[5332] <= 15'b011111010011111;
		Coeff[5333] <= 15'b011111010100010;
		Coeff[5334] <= 15'b011111010100100;
		Coeff[5335] <= 15'b011111010100111;
		Coeff[5336] <= 15'b011111010101010;
		Coeff[5337] <= 15'b011111010101101;
		Coeff[5338] <= 15'b011111010101111;
		Coeff[5339] <= 15'b011111010110010;
		Coeff[5340] <= 15'b011111010110101;
		Coeff[5341] <= 15'b011111010111000;
		Coeff[5342] <= 15'b011111010111010;
		Coeff[5343] <= 15'b011111010111101;
		Coeff[5344] <= 15'b011111011000000;
		Coeff[5345] <= 15'b011111011000010;
		Coeff[5346] <= 15'b011111011000101;
		Coeff[5347] <= 15'b011111011001000;
		Coeff[5348] <= 15'b011111011001011;
		Coeff[5349] <= 15'b011111011001101;
		Coeff[5350] <= 15'b011111011010000;
		Coeff[5351] <= 15'b011111011010011;
		Coeff[5352] <= 15'b011111011010110;
		Coeff[5353] <= 15'b011111011011000;
		Coeff[5354] <= 15'b011111011011011;
		Coeff[5355] <= 15'b011111011011110;
		Coeff[5356] <= 15'b011111011100001;
		Coeff[5357] <= 15'b011111011100011;
		Coeff[5358] <= 15'b011111011100110;
		Coeff[5359] <= 15'b011111011101001;
		Coeff[5360] <= 15'b011111011101100;
		Coeff[5361] <= 15'b011111011101110;
		Coeff[5362] <= 15'b011111011110001;
		Coeff[5363] <= 15'b011111011110100;
		Coeff[5364] <= 15'b011111011110110;
		Coeff[5365] <= 15'b011111011111001;
		Coeff[5366] <= 15'b011111011111100;
		Coeff[5367] <= 15'b011111011111111;
		Coeff[5368] <= 15'b011111100000001;
		Coeff[5369] <= 15'b011111100000100;
		Coeff[5370] <= 15'b011111100000111;
		Coeff[5371] <= 15'b011111100001010;
		Coeff[5372] <= 15'b011111100001100;
		Coeff[5373] <= 15'b011111100001111;
		Coeff[5374] <= 15'b011111100010010;
		Coeff[5375] <= 15'b011111100010101;
		Coeff[5376] <= 15'b011111100010111;
		Coeff[5377] <= 15'b011111100011010;
		Coeff[5378] <= 15'b011111100011101;
		Coeff[5379] <= 15'b011111100011111;
		Coeff[5380] <= 15'b011111100100010;
		Coeff[5381] <= 15'b011111100100101;
		Coeff[5382] <= 15'b011111100101000;
		Coeff[5383] <= 15'b011111100101010;
		Coeff[5384] <= 15'b011111100101101;
		Coeff[5385] <= 15'b011111100110000;
		Coeff[5386] <= 15'b011111100110011;
		Coeff[5387] <= 15'b011111100110101;
		Coeff[5388] <= 15'b011111100111000;
		Coeff[5389] <= 15'b011111100111011;
		Coeff[5390] <= 15'b011111100111110;
		Coeff[5391] <= 15'b011111101000000;
		Coeff[5392] <= 15'b011111101000011;
		Coeff[5393] <= 15'b011111101000110;
		Coeff[5394] <= 15'b011111101001000;
		Coeff[5395] <= 15'b011111101001011;
		Coeff[5396] <= 15'b011111101001110;
		Coeff[5397] <= 15'b011111101010001;
		Coeff[5398] <= 15'b011111101010011;
		Coeff[5399] <= 15'b011111101010110;
		Coeff[5400] <= 15'b011111101011001;
		Coeff[5401] <= 15'b011111101011100;
		Coeff[5402] <= 15'b011111101011110;
		Coeff[5403] <= 15'b011111101100001;
		Coeff[5404] <= 15'b011111101100100;
		Coeff[5405] <= 15'b011111101100110;
		Coeff[5406] <= 15'b011111101101001;
		Coeff[5407] <= 15'b011111101101100;
		Coeff[5408] <= 15'b011111101101111;
		Coeff[5409] <= 15'b011111101110001;
		Coeff[5410] <= 15'b011111101110100;
		Coeff[5411] <= 15'b011111101110111;
		Coeff[5412] <= 15'b011111101111010;
		Coeff[5413] <= 15'b011111101111100;
		Coeff[5414] <= 15'b011111101111111;
		Coeff[5415] <= 15'b011111110000010;
		Coeff[5416] <= 15'b011111110000101;
		Coeff[5417] <= 15'b011111110000111;
		Coeff[5418] <= 15'b011111110001010;
		Coeff[5419] <= 15'b011111110001101;
		Coeff[5420] <= 15'b011111110001111;
		Coeff[5421] <= 15'b011111110010010;
		Coeff[5422] <= 15'b011111110010101;
		Coeff[5423] <= 15'b011111110011000;
		Coeff[5424] <= 15'b011111110011010;
		Coeff[5425] <= 15'b011111110011101;
		Coeff[5426] <= 15'b011111110100000;
		Coeff[5427] <= 15'b011111110100011;
		Coeff[5428] <= 15'b011111110100101;
		Coeff[5429] <= 15'b011111110101000;
		Coeff[5430] <= 15'b011111110101011;
		Coeff[5431] <= 15'b011111110101101;
		Coeff[5432] <= 15'b011111110110000;
		Coeff[5433] <= 15'b011111110110011;
		Coeff[5434] <= 15'b011111110110110;
		Coeff[5435] <= 15'b011111110111000;
		Coeff[5436] <= 15'b011111110111011;
		Coeff[5437] <= 15'b011111110111110;
		Coeff[5438] <= 15'b011111111000000;
		Coeff[5439] <= 15'b011111111000011;
		Coeff[5440] <= 15'b011111111000110;
		Coeff[5441] <= 15'b011111111001001;
		Coeff[5442] <= 15'b011111111001011;
		Coeff[5443] <= 15'b011111111001110;
		Coeff[5444] <= 15'b011111111010001;
		Coeff[5445] <= 15'b011111111010100;
		Coeff[5446] <= 15'b011111111010110;
		Coeff[5447] <= 15'b011111111011001;
		Coeff[5448] <= 15'b011111111011100;
		Coeff[5449] <= 15'b011111111011110;
		Coeff[5450] <= 15'b011111111100001;
		Coeff[5451] <= 15'b011111111100100;
		Coeff[5452] <= 15'b011111111100111;
		Coeff[5453] <= 15'b011111111101001;
		Coeff[5454] <= 15'b011111111101100;
		Coeff[5455] <= 15'b011111111101111;
		Coeff[5456] <= 15'b011111111110001;
		Coeff[5457] <= 15'b011111111110100;
		Coeff[5458] <= 15'b011111111110111;
		Coeff[5459] <= 15'b011111111111010;
		Coeff[5460] <= 15'b011111111111100;
		Coeff[5461] <= 15'b011111111111111;
		Coeff[5462] <= 15'b100000000000010;
		Coeff[5463] <= 15'b100000000000101;
		Coeff[5464] <= 15'b100000000000111;
		Coeff[5465] <= 15'b100000000001010;
		Coeff[5466] <= 15'b100000000001101;
		Coeff[5467] <= 15'b100000000001111;
		Coeff[5468] <= 15'b100000000010010;
		Coeff[5469] <= 15'b100000000010101;
		Coeff[5470] <= 15'b100000000011000;
		Coeff[5471] <= 15'b100000000011010;
		Coeff[5472] <= 15'b100000000011101;
		Coeff[5473] <= 15'b100000000100000;
		Coeff[5474] <= 15'b100000000100010;
		Coeff[5475] <= 15'b100000000100101;
		Coeff[5476] <= 15'b100000000101000;
		Coeff[5477] <= 15'b100000000101011;
		Coeff[5478] <= 15'b100000000101101;
		Coeff[5479] <= 15'b100000000110000;
		Coeff[5480] <= 15'b100000000110011;
		Coeff[5481] <= 15'b100000000110101;
		Coeff[5482] <= 15'b100000000111000;
		Coeff[5483] <= 15'b100000000111011;
		Coeff[5484] <= 15'b100000000111110;
		Coeff[5485] <= 15'b100000001000000;
		Coeff[5486] <= 15'b100000001000011;
		Coeff[5487] <= 15'b100000001000110;
		Coeff[5488] <= 15'b100000001001000;
		Coeff[5489] <= 15'b100000001001011;
		Coeff[5490] <= 15'b100000001001110;
		Coeff[5491] <= 15'b100000001010001;
		Coeff[5492] <= 15'b100000001010011;
		Coeff[5493] <= 15'b100000001010110;
		Coeff[5494] <= 15'b100000001011001;
		Coeff[5495] <= 15'b100000001011100;
		Coeff[5496] <= 15'b100000001011110;
		Coeff[5497] <= 15'b100000001100001;
		Coeff[5498] <= 15'b100000001100100;
		Coeff[5499] <= 15'b100000001100110;
		Coeff[5500] <= 15'b100000001101001;
		Coeff[5501] <= 15'b100000001101100;
		Coeff[5502] <= 15'b100000001101111;
		Coeff[5503] <= 15'b100000001110001;
		Coeff[5504] <= 15'b100000001110100;
		Coeff[5505] <= 15'b100000001110111;
		Coeff[5506] <= 15'b100000001111001;
		Coeff[5507] <= 15'b100000001111100;
		Coeff[5508] <= 15'b100000001111111;
		Coeff[5509] <= 15'b100000010000010;
		Coeff[5510] <= 15'b100000010000100;
		Coeff[5511] <= 15'b100000010000111;
		Coeff[5512] <= 15'b100000010001010;
		Coeff[5513] <= 15'b100000010001100;
		Coeff[5514] <= 15'b100000010001111;
		Coeff[5515] <= 15'b100000010010010;
		Coeff[5516] <= 15'b100000010010101;
		Coeff[5517] <= 15'b100000010010111;
		Coeff[5518] <= 15'b100000010011010;
		Coeff[5519] <= 15'b100000010011101;
		Coeff[5520] <= 15'b100000010011111;
		Coeff[5521] <= 15'b100000010100010;
		Coeff[5522] <= 15'b100000010100101;
		Coeff[5523] <= 15'b100000010100111;
		Coeff[5524] <= 15'b100000010101010;
		Coeff[5525] <= 15'b100000010101101;
		Coeff[5526] <= 15'b100000010110000;
		Coeff[5527] <= 15'b100000010110010;
		Coeff[5528] <= 15'b100000010110101;
		Coeff[5529] <= 15'b100000010111000;
		Coeff[5530] <= 15'b100000010111010;
		Coeff[5531] <= 15'b100000010111101;
		Coeff[5532] <= 15'b100000011000000;
		Coeff[5533] <= 15'b100000011000011;
		Coeff[5534] <= 15'b100000011000101;
		Coeff[5535] <= 15'b100000011001000;
		Coeff[5536] <= 15'b100000011001011;
		Coeff[5537] <= 15'b100000011001101;
		Coeff[5538] <= 15'b100000011010000;
		Coeff[5539] <= 15'b100000011010011;
		Coeff[5540] <= 15'b100000011010110;
		Coeff[5541] <= 15'b100000011011000;
		Coeff[5542] <= 15'b100000011011011;
		Coeff[5543] <= 15'b100000011011110;
		Coeff[5544] <= 15'b100000011100000;
		Coeff[5545] <= 15'b100000011100011;
		Coeff[5546] <= 15'b100000011100110;
		Coeff[5547] <= 15'b100000011101001;
		Coeff[5548] <= 15'b100000011101011;
		Coeff[5549] <= 15'b100000011101110;
		Coeff[5550] <= 15'b100000011110001;
		Coeff[5551] <= 15'b100000011110011;
		Coeff[5552] <= 15'b100000011110110;
		Coeff[5553] <= 15'b100000011111001;
		Coeff[5554] <= 15'b100000011111011;
		Coeff[5555] <= 15'b100000011111110;
		Coeff[5556] <= 15'b100000100000001;
		Coeff[5557] <= 15'b100000100000100;
		Coeff[5558] <= 15'b100000100000110;
		Coeff[5559] <= 15'b100000100001001;
		Coeff[5560] <= 15'b100000100001100;
		Coeff[5561] <= 15'b100000100001110;
		Coeff[5562] <= 15'b100000100010001;
		Coeff[5563] <= 15'b100000100010100;
		Coeff[5564] <= 15'b100000100010111;
		Coeff[5565] <= 15'b100000100011001;
		Coeff[5566] <= 15'b100000100011100;
		Coeff[5567] <= 15'b100000100011111;
		Coeff[5568] <= 15'b100000100100001;
		Coeff[5569] <= 15'b100000100100100;
		Coeff[5570] <= 15'b100000100100111;
		Coeff[5571] <= 15'b100000100101001;
		Coeff[5572] <= 15'b100000100101100;
		Coeff[5573] <= 15'b100000100101111;
		Coeff[5574] <= 15'b100000100110010;
		Coeff[5575] <= 15'b100000100110100;
		Coeff[5576] <= 15'b100000100110111;
		Coeff[5577] <= 15'b100000100111010;
		Coeff[5578] <= 15'b100000100111100;
		Coeff[5579] <= 15'b100000100111111;
		Coeff[5580] <= 15'b100000101000010;
		Coeff[5581] <= 15'b100000101000100;
		Coeff[5582] <= 15'b100000101000111;
		Coeff[5583] <= 15'b100000101001010;
		Coeff[5584] <= 15'b100000101001101;
		Coeff[5585] <= 15'b100000101001111;
		Coeff[5586] <= 15'b100000101010010;
		Coeff[5587] <= 15'b100000101010101;
		Coeff[5588] <= 15'b100000101010111;
		Coeff[5589] <= 15'b100000101011010;
		Coeff[5590] <= 15'b100000101011101;
		Coeff[5591] <= 15'b100000101100000;
		Coeff[5592] <= 15'b100000101100010;
		Coeff[5593] <= 15'b100000101100101;
		Coeff[5594] <= 15'b100000101101000;
		Coeff[5595] <= 15'b100000101101010;
		Coeff[5596] <= 15'b100000101101101;
		Coeff[5597] <= 15'b100000101110000;
		Coeff[5598] <= 15'b100000101110010;
		Coeff[5599] <= 15'b100000101110101;
		Coeff[5600] <= 15'b100000101111000;
		Coeff[5601] <= 15'b100000101111011;
		Coeff[5602] <= 15'b100000101111101;
		Coeff[5603] <= 15'b100000110000000;
		Coeff[5604] <= 15'b100000110000011;
		Coeff[5605] <= 15'b100000110000101;
		Coeff[5606] <= 15'b100000110001000;
		Coeff[5607] <= 15'b100000110001011;
		Coeff[5608] <= 15'b100000110001101;
		Coeff[5609] <= 15'b100000110010000;
		Coeff[5610] <= 15'b100000110010011;
		Coeff[5611] <= 15'b100000110010101;
		Coeff[5612] <= 15'b100000110011000;
		Coeff[5613] <= 15'b100000110011011;
		Coeff[5614] <= 15'b100000110011110;
		Coeff[5615] <= 15'b100000110100000;
		Coeff[5616] <= 15'b100000110100011;
		Coeff[5617] <= 15'b100000110100110;
		Coeff[5618] <= 15'b100000110101000;
		Coeff[5619] <= 15'b100000110101011;
		Coeff[5620] <= 15'b100000110101110;
		Coeff[5621] <= 15'b100000110110000;
		Coeff[5622] <= 15'b100000110110011;
		Coeff[5623] <= 15'b100000110110110;
		Coeff[5624] <= 15'b100000110111001;
		Coeff[5625] <= 15'b100000110111011;
		Coeff[5626] <= 15'b100000110111110;
		Coeff[5627] <= 15'b100000111000001;
		Coeff[5628] <= 15'b100000111000011;
		Coeff[5629] <= 15'b100000111000110;
		Coeff[5630] <= 15'b100000111001001;
		Coeff[5631] <= 15'b100000111001011;
		Coeff[5632] <= 15'b100000111001110;
		Coeff[5633] <= 15'b100000111010001;
		Coeff[5634] <= 15'b100000111010100;
		Coeff[5635] <= 15'b100000111010110;
		Coeff[5636] <= 15'b100000111011001;
		Coeff[5637] <= 15'b100000111011100;
		Coeff[5638] <= 15'b100000111011110;
		Coeff[5639] <= 15'b100000111100001;
		Coeff[5640] <= 15'b100000111100100;
		Coeff[5641] <= 15'b100000111100110;
		Coeff[5642] <= 15'b100000111101001;
		Coeff[5643] <= 15'b100000111101100;
		Coeff[5644] <= 15'b100000111101110;
		Coeff[5645] <= 15'b100000111110001;
		Coeff[5646] <= 15'b100000111110100;
		Coeff[5647] <= 15'b100000111110111;
		Coeff[5648] <= 15'b100000111111001;
		Coeff[5649] <= 15'b100000111111100;
		Coeff[5650] <= 15'b100000111111111;
		Coeff[5651] <= 15'b100001000000001;
		Coeff[5652] <= 15'b100001000000100;
		Coeff[5653] <= 15'b100001000000111;
		Coeff[5654] <= 15'b100001000001001;
		Coeff[5655] <= 15'b100001000001100;
		Coeff[5656] <= 15'b100001000001111;
		Coeff[5657] <= 15'b100001000010001;
		Coeff[5658] <= 15'b100001000010100;
		Coeff[5659] <= 15'b100001000010111;
		Coeff[5660] <= 15'b100001000011010;
		Coeff[5661] <= 15'b100001000011100;
		Coeff[5662] <= 15'b100001000011111;
		Coeff[5663] <= 15'b100001000100010;
		Coeff[5664] <= 15'b100001000100100;
		Coeff[5665] <= 15'b100001000100111;
		Coeff[5666] <= 15'b100001000101010;
		Coeff[5667] <= 15'b100001000101100;
		Coeff[5668] <= 15'b100001000101111;
		Coeff[5669] <= 15'b100001000110010;
		Coeff[5670] <= 15'b100001000110100;
		Coeff[5671] <= 15'b100001000110111;
		Coeff[5672] <= 15'b100001000111010;
		Coeff[5673] <= 15'b100001000111100;
		Coeff[5674] <= 15'b100001000111111;
		Coeff[5675] <= 15'b100001001000010;
		Coeff[5676] <= 15'b100001001000101;
		Coeff[5677] <= 15'b100001001000111;
		Coeff[5678] <= 15'b100001001001010;
		Coeff[5679] <= 15'b100001001001101;
		Coeff[5680] <= 15'b100001001001111;
		Coeff[5681] <= 15'b100001001010010;
		Coeff[5682] <= 15'b100001001010101;
		Coeff[5683] <= 15'b100001001010111;
		Coeff[5684] <= 15'b100001001011010;
		Coeff[5685] <= 15'b100001001011101;
		Coeff[5686] <= 15'b100001001011111;
		Coeff[5687] <= 15'b100001001100010;
		Coeff[5688] <= 15'b100001001100101;
		Coeff[5689] <= 15'b100001001100111;
		Coeff[5690] <= 15'b100001001101010;
		Coeff[5691] <= 15'b100001001101101;
		Coeff[5692] <= 15'b100001001110000;
		Coeff[5693] <= 15'b100001001110010;
		Coeff[5694] <= 15'b100001001110101;
		Coeff[5695] <= 15'b100001001111000;
		Coeff[5696] <= 15'b100001001111010;
		Coeff[5697] <= 15'b100001001111101;
		Coeff[5698] <= 15'b100001010000000;
		Coeff[5699] <= 15'b100001010000010;
		Coeff[5700] <= 15'b100001010000101;
		Coeff[5701] <= 15'b100001010001000;
		Coeff[5702] <= 15'b100001010001010;
		Coeff[5703] <= 15'b100001010001101;
		Coeff[5704] <= 15'b100001010010000;
		Coeff[5705] <= 15'b100001010010010;
		Coeff[5706] <= 15'b100001010010101;
		Coeff[5707] <= 15'b100001010011000;
		Coeff[5708] <= 15'b100001010011010;
		Coeff[5709] <= 15'b100001010011101;
		Coeff[5710] <= 15'b100001010100000;
		Coeff[5711] <= 15'b100001010100011;
		Coeff[5712] <= 15'b100001010100101;
		Coeff[5713] <= 15'b100001010101000;
		Coeff[5714] <= 15'b100001010101011;
		Coeff[5715] <= 15'b100001010101101;
		Coeff[5716] <= 15'b100001010110000;
		Coeff[5717] <= 15'b100001010110011;
		Coeff[5718] <= 15'b100001010110101;
		Coeff[5719] <= 15'b100001010111000;
		Coeff[5720] <= 15'b100001010111011;
		Coeff[5721] <= 15'b100001010111101;
		Coeff[5722] <= 15'b100001011000000;
		Coeff[5723] <= 15'b100001011000011;
		Coeff[5724] <= 15'b100001011000101;
		Coeff[5725] <= 15'b100001011001000;
		Coeff[5726] <= 15'b100001011001011;
		Coeff[5727] <= 15'b100001011001101;
		Coeff[5728] <= 15'b100001011010000;
		Coeff[5729] <= 15'b100001011010011;
		Coeff[5730] <= 15'b100001011010101;
		Coeff[5731] <= 15'b100001011011000;
		Coeff[5732] <= 15'b100001011011011;
		Coeff[5733] <= 15'b100001011011101;
		Coeff[5734] <= 15'b100001011100000;
		Coeff[5735] <= 15'b100001011100011;
		Coeff[5736] <= 15'b100001011100110;
		Coeff[5737] <= 15'b100001011101000;
		Coeff[5738] <= 15'b100001011101011;
		Coeff[5739] <= 15'b100001011101110;
		Coeff[5740] <= 15'b100001011110000;
		Coeff[5741] <= 15'b100001011110011;
		Coeff[5742] <= 15'b100001011110110;
		Coeff[5743] <= 15'b100001011111000;
		Coeff[5744] <= 15'b100001011111011;
		Coeff[5745] <= 15'b100001011111110;
		Coeff[5746] <= 15'b100001100000000;
		Coeff[5747] <= 15'b100001100000011;
		Coeff[5748] <= 15'b100001100000110;
		Coeff[5749] <= 15'b100001100001000;
		Coeff[5750] <= 15'b100001100001011;
		Coeff[5751] <= 15'b100001100001110;
		Coeff[5752] <= 15'b100001100010000;
		Coeff[5753] <= 15'b100001100010011;
		Coeff[5754] <= 15'b100001100010110;
		Coeff[5755] <= 15'b100001100011000;
		Coeff[5756] <= 15'b100001100011011;
		Coeff[5757] <= 15'b100001100011110;
		Coeff[5758] <= 15'b100001100100000;
		Coeff[5759] <= 15'b100001100100011;
		Coeff[5760] <= 15'b100001100100110;
		Coeff[5761] <= 15'b100001100101000;
		Coeff[5762] <= 15'b100001100101011;
		Coeff[5763] <= 15'b100001100101110;
		Coeff[5764] <= 15'b100001100110000;
		Coeff[5765] <= 15'b100001100110011;
		Coeff[5766] <= 15'b100001100110110;
		Coeff[5767] <= 15'b100001100111000;
		Coeff[5768] <= 15'b100001100111011;
		Coeff[5769] <= 15'b100001100111110;
		Coeff[5770] <= 15'b100001101000000;
		Coeff[5771] <= 15'b100001101000011;
		Coeff[5772] <= 15'b100001101000110;
		Coeff[5773] <= 15'b100001101001001;
		Coeff[5774] <= 15'b100001101001011;
		Coeff[5775] <= 15'b100001101001110;
		Coeff[5776] <= 15'b100001101010001;
		Coeff[5777] <= 15'b100001101010011;
		Coeff[5778] <= 15'b100001101010110;
		Coeff[5779] <= 15'b100001101011001;
		Coeff[5780] <= 15'b100001101011011;
		Coeff[5781] <= 15'b100001101011110;
		Coeff[5782] <= 15'b100001101100001;
		Coeff[5783] <= 15'b100001101100011;
		Coeff[5784] <= 15'b100001101100110;
		Coeff[5785] <= 15'b100001101101001;
		Coeff[5786] <= 15'b100001101101011;
		Coeff[5787] <= 15'b100001101101110;
		Coeff[5788] <= 15'b100001101110001;
		Coeff[5789] <= 15'b100001101110011;
		Coeff[5790] <= 15'b100001101110110;
		Coeff[5791] <= 15'b100001101111001;
		Coeff[5792] <= 15'b100001101111011;
		Coeff[5793] <= 15'b100001101111110;
		Coeff[5794] <= 15'b100001110000001;
		Coeff[5795] <= 15'b100001110000011;
		Coeff[5796] <= 15'b100001110000110;
		Coeff[5797] <= 15'b100001110001001;
		Coeff[5798] <= 15'b100001110001011;
		Coeff[5799] <= 15'b100001110001110;
		Coeff[5800] <= 15'b100001110010001;
		Coeff[5801] <= 15'b100001110010011;
		Coeff[5802] <= 15'b100001110010110;
		Coeff[5803] <= 15'b100001110011001;
		Coeff[5804] <= 15'b100001110011011;
		Coeff[5805] <= 15'b100001110011110;
		Coeff[5806] <= 15'b100001110100001;
		Coeff[5807] <= 15'b100001110100011;
		Coeff[5808] <= 15'b100001110100110;
		Coeff[5809] <= 15'b100001110101001;
		Coeff[5810] <= 15'b100001110101011;
		Coeff[5811] <= 15'b100001110101110;
		Coeff[5812] <= 15'b100001110110001;
		Coeff[5813] <= 15'b100001110110011;
		Coeff[5814] <= 15'b100001110110110;
		Coeff[5815] <= 15'b100001110111001;
		Coeff[5816] <= 15'b100001110111011;
		Coeff[5817] <= 15'b100001110111110;
		Coeff[5818] <= 15'b100001111000001;
		Coeff[5819] <= 15'b100001111000011;
		Coeff[5820] <= 15'b100001111000110;
		Coeff[5821] <= 15'b100001111001001;
		Coeff[5822] <= 15'b100001111001011;
		Coeff[5823] <= 15'b100001111001110;
		Coeff[5824] <= 15'b100001111010001;
		Coeff[5825] <= 15'b100001111010011;
		Coeff[5826] <= 15'b100001111010110;
		Coeff[5827] <= 15'b100001111011001;
		Coeff[5828] <= 15'b100001111011011;
		Coeff[5829] <= 15'b100001111011110;
		Coeff[5830] <= 15'b100001111100001;
		Coeff[5831] <= 15'b100001111100011;
		Coeff[5832] <= 15'b100001111100110;
		Coeff[5833] <= 15'b100001111101001;
		Coeff[5834] <= 15'b100001111101011;
		Coeff[5835] <= 15'b100001111101110;
		Coeff[5836] <= 15'b100001111110001;
		Coeff[5837] <= 15'b100001111110011;
		Coeff[5838] <= 15'b100001111110110;
		Coeff[5839] <= 15'b100001111111001;
		Coeff[5840] <= 15'b100001111111011;
		Coeff[5841] <= 15'b100001111111110;
		Coeff[5842] <= 15'b100010000000001;
		Coeff[5843] <= 15'b100010000000011;
		Coeff[5844] <= 15'b100010000000110;
		Coeff[5845] <= 15'b100010000001001;
		Coeff[5846] <= 15'b100010000001011;
		Coeff[5847] <= 15'b100010000001110;
		Coeff[5848] <= 15'b100010000010001;
		Coeff[5849] <= 15'b100010000010011;
		Coeff[5850] <= 15'b100010000010110;
		Coeff[5851] <= 15'b100010000011000;
		Coeff[5852] <= 15'b100010000011011;
		Coeff[5853] <= 15'b100010000011110;
		Coeff[5854] <= 15'b100010000100000;
		Coeff[5855] <= 15'b100010000100011;
		Coeff[5856] <= 15'b100010000100110;
		Coeff[5857] <= 15'b100010000101000;
		Coeff[5858] <= 15'b100010000101011;
		Coeff[5859] <= 15'b100010000101110;
		Coeff[5860] <= 15'b100010000110000;
		Coeff[5861] <= 15'b100010000110011;
		Coeff[5862] <= 15'b100010000110110;
		Coeff[5863] <= 15'b100010000111000;
		Coeff[5864] <= 15'b100010000111011;
		Coeff[5865] <= 15'b100010000111110;
		Coeff[5866] <= 15'b100010001000000;
		Coeff[5867] <= 15'b100010001000011;
		Coeff[5868] <= 15'b100010001000110;
		Coeff[5869] <= 15'b100010001001000;
		Coeff[5870] <= 15'b100010001001011;
		Coeff[5871] <= 15'b100010001001110;
		Coeff[5872] <= 15'b100010001010000;
		Coeff[5873] <= 15'b100010001010011;
		Coeff[5874] <= 15'b100010001010110;
		Coeff[5875] <= 15'b100010001011000;
		Coeff[5876] <= 15'b100010001011011;
		Coeff[5877] <= 15'b100010001011110;
		Coeff[5878] <= 15'b100010001100000;
		Coeff[5879] <= 15'b100010001100011;
		Coeff[5880] <= 15'b100010001100110;
		Coeff[5881] <= 15'b100010001101000;
		Coeff[5882] <= 15'b100010001101011;
		Coeff[5883] <= 15'b100010001101110;
		Coeff[5884] <= 15'b100010001110000;
		Coeff[5885] <= 15'b100010001110011;
		Coeff[5886] <= 15'b100010001110101;
		Coeff[5887] <= 15'b100010001111000;
		Coeff[5888] <= 15'b100010001111011;
		Coeff[5889] <= 15'b100010001111101;
		Coeff[5890] <= 15'b100010010000000;
		Coeff[5891] <= 15'b100010010000011;
		Coeff[5892] <= 15'b100010010000101;
		Coeff[5893] <= 15'b100010010001000;
		Coeff[5894] <= 15'b100010010001011;
		Coeff[5895] <= 15'b100010010001101;
		Coeff[5896] <= 15'b100010010010000;
		Coeff[5897] <= 15'b100010010010011;
		Coeff[5898] <= 15'b100010010010101;
		Coeff[5899] <= 15'b100010010011000;
		Coeff[5900] <= 15'b100010010011011;
		Coeff[5901] <= 15'b100010010011101;
		Coeff[5902] <= 15'b100010010100000;
		Coeff[5903] <= 15'b100010010100011;
		Coeff[5904] <= 15'b100010010100101;
		Coeff[5905] <= 15'b100010010101000;
		Coeff[5906] <= 15'b100010010101011;
		Coeff[5907] <= 15'b100010010101101;
		Coeff[5908] <= 15'b100010010110000;
		Coeff[5909] <= 15'b100010010110011;
		Coeff[5910] <= 15'b100010010110101;
		Coeff[5911] <= 15'b100010010111000;
		Coeff[5912] <= 15'b100010010111010;
		Coeff[5913] <= 15'b100010010111101;
		Coeff[5914] <= 15'b100010011000000;
		Coeff[5915] <= 15'b100010011000010;
		Coeff[5916] <= 15'b100010011000101;
		Coeff[5917] <= 15'b100010011001000;
		Coeff[5918] <= 15'b100010011001010;
		Coeff[5919] <= 15'b100010011001101;
		Coeff[5920] <= 15'b100010011010000;
		Coeff[5921] <= 15'b100010011010010;
		Coeff[5922] <= 15'b100010011010101;
		Coeff[5923] <= 15'b100010011011000;
		Coeff[5924] <= 15'b100010011011010;
		Coeff[5925] <= 15'b100010011011101;
		Coeff[5926] <= 15'b100010011100000;
		Coeff[5927] <= 15'b100010011100010;
		Coeff[5928] <= 15'b100010011100101;
		Coeff[5929] <= 15'b100010011100111;
		Coeff[5930] <= 15'b100010011101010;
		Coeff[5931] <= 15'b100010011101101;
		Coeff[5932] <= 15'b100010011101111;
		Coeff[5933] <= 15'b100010011110010;
		Coeff[5934] <= 15'b100010011110101;
		Coeff[5935] <= 15'b100010011110111;
		Coeff[5936] <= 15'b100010011111010;
		Coeff[5937] <= 15'b100010011111101;
		Coeff[5938] <= 15'b100010011111111;
		Coeff[5939] <= 15'b100010100000010;
		Coeff[5940] <= 15'b100010100000101;
		Coeff[5941] <= 15'b100010100000111;
		Coeff[5942] <= 15'b100010100001010;
		Coeff[5943] <= 15'b100010100001101;
		Coeff[5944] <= 15'b100010100001111;
		Coeff[5945] <= 15'b100010100010010;
		Coeff[5946] <= 15'b100010100010100;
		Coeff[5947] <= 15'b100010100010111;
		Coeff[5948] <= 15'b100010100011010;
		Coeff[5949] <= 15'b100010100011100;
		Coeff[5950] <= 15'b100010100011111;
		Coeff[5951] <= 15'b100010100100010;
		Coeff[5952] <= 15'b100010100100100;
		Coeff[5953] <= 15'b100010100100111;
		Coeff[5954] <= 15'b100010100101010;
		Coeff[5955] <= 15'b100010100101100;
		Coeff[5956] <= 15'b100010100101111;
		Coeff[5957] <= 15'b100010100110010;
		Coeff[5958] <= 15'b100010100110100;
		Coeff[5959] <= 15'b100010100110111;
		Coeff[5960] <= 15'b100010100111001;
		Coeff[5961] <= 15'b100010100111100;
		Coeff[5962] <= 15'b100010100111111;
		Coeff[5963] <= 15'b100010101000001;
		Coeff[5964] <= 15'b100010101000100;
		Coeff[5965] <= 15'b100010101000111;
		Coeff[5966] <= 15'b100010101001001;
		Coeff[5967] <= 15'b100010101001100;
		Coeff[5968] <= 15'b100010101001111;
		Coeff[5969] <= 15'b100010101010001;
		Coeff[5970] <= 15'b100010101010100;
		Coeff[5971] <= 15'b100010101010111;
		Coeff[5972] <= 15'b100010101011001;
		Coeff[5973] <= 15'b100010101011100;
		Coeff[5974] <= 15'b100010101011110;
		Coeff[5975] <= 15'b100010101100001;
		Coeff[5976] <= 15'b100010101100100;
		Coeff[5977] <= 15'b100010101100110;
		Coeff[5978] <= 15'b100010101101001;
		Coeff[5979] <= 15'b100010101101100;
		Coeff[5980] <= 15'b100010101101110;
		Coeff[5981] <= 15'b100010101110001;
		Coeff[5982] <= 15'b100010101110100;
		Coeff[5983] <= 15'b100010101110110;
		Coeff[5984] <= 15'b100010101111001;
		Coeff[5985] <= 15'b100010101111011;
		Coeff[5986] <= 15'b100010101111110;
		Coeff[5987] <= 15'b100010110000001;
		Coeff[5988] <= 15'b100010110000011;
		Coeff[5989] <= 15'b100010110000110;
		Coeff[5990] <= 15'b100010110001001;
		Coeff[5991] <= 15'b100010110001011;
		Coeff[5992] <= 15'b100010110001110;
		Coeff[5993] <= 15'b100010110010001;
		Coeff[5994] <= 15'b100010110010011;
		Coeff[5995] <= 15'b100010110010110;
		Coeff[5996] <= 15'b100010110011001;
		Coeff[5997] <= 15'b100010110011011;
		Coeff[5998] <= 15'b100010110011110;
		Coeff[5999] <= 15'b100010110100000;
		Coeff[6000] <= 15'b100010110100011;
		Coeff[6001] <= 15'b100010110100110;
		Coeff[6002] <= 15'b100010110101000;
		Coeff[6003] <= 15'b100010110101011;
		Coeff[6004] <= 15'b100010110101110;
		Coeff[6005] <= 15'b100010110110000;
		Coeff[6006] <= 15'b100010110110011;
		Coeff[6007] <= 15'b100010110110110;
		Coeff[6008] <= 15'b100010110111000;
		Coeff[6009] <= 15'b100010110111011;
		Coeff[6010] <= 15'b100010110111101;
		Coeff[6011] <= 15'b100010111000000;
		Coeff[6012] <= 15'b100010111000011;
		Coeff[6013] <= 15'b100010111000101;
		Coeff[6014] <= 15'b100010111001000;
		Coeff[6015] <= 15'b100010111001011;
		Coeff[6016] <= 15'b100010111001101;
		Coeff[6017] <= 15'b100010111010000;
		Coeff[6018] <= 15'b100010111010010;
		Coeff[6019] <= 15'b100010111010101;
		Coeff[6020] <= 15'b100010111011000;
		Coeff[6021] <= 15'b100010111011010;
		Coeff[6022] <= 15'b100010111011101;
		Coeff[6023] <= 15'b100010111100000;
		Coeff[6024] <= 15'b100010111100010;
		Coeff[6025] <= 15'b100010111100101;
		Coeff[6026] <= 15'b100010111101000;
		Coeff[6027] <= 15'b100010111101010;
		Coeff[6028] <= 15'b100010111101101;
		Coeff[6029] <= 15'b100010111101111;
		Coeff[6030] <= 15'b100010111110010;
		Coeff[6031] <= 15'b100010111110101;
		Coeff[6032] <= 15'b100010111110111;
		Coeff[6033] <= 15'b100010111111010;
		Coeff[6034] <= 15'b100010111111101;
		Coeff[6035] <= 15'b100010111111111;
		Coeff[6036] <= 15'b100011000000010;
		Coeff[6037] <= 15'b100011000000100;
		Coeff[6038] <= 15'b100011000000111;
		Coeff[6039] <= 15'b100011000001010;
		Coeff[6040] <= 15'b100011000001100;
		Coeff[6041] <= 15'b100011000001111;
		Coeff[6042] <= 15'b100011000010010;
		Coeff[6043] <= 15'b100011000010100;
		Coeff[6044] <= 15'b100011000010111;
		Coeff[6045] <= 15'b100011000011010;
		Coeff[6046] <= 15'b100011000011100;
		Coeff[6047] <= 15'b100011000011111;
		Coeff[6048] <= 15'b100011000100001;
		Coeff[6049] <= 15'b100011000100100;
		Coeff[6050] <= 15'b100011000100111;
		Coeff[6051] <= 15'b100011000101001;
		Coeff[6052] <= 15'b100011000101100;
		Coeff[6053] <= 15'b100011000101111;
		Coeff[6054] <= 15'b100011000110001;
		Coeff[6055] <= 15'b100011000110100;
		Coeff[6056] <= 15'b100011000110110;
		Coeff[6057] <= 15'b100011000111001;
		Coeff[6058] <= 15'b100011000111100;
		Coeff[6059] <= 15'b100011000111110;
		Coeff[6060] <= 15'b100011001000001;
		Coeff[6061] <= 15'b100011001000100;
		Coeff[6062] <= 15'b100011001000110;
		Coeff[6063] <= 15'b100011001001001;
		Coeff[6064] <= 15'b100011001001011;
		Coeff[6065] <= 15'b100011001001110;
		Coeff[6066] <= 15'b100011001010001;
		Coeff[6067] <= 15'b100011001010011;
		Coeff[6068] <= 15'b100011001010110;
		Coeff[6069] <= 15'b100011001011001;
		Coeff[6070] <= 15'b100011001011011;
		Coeff[6071] <= 15'b100011001011110;
		Coeff[6072] <= 15'b100011001100000;
		Coeff[6073] <= 15'b100011001100011;
		Coeff[6074] <= 15'b100011001100110;
		Coeff[6075] <= 15'b100011001101000;
		Coeff[6076] <= 15'b100011001101011;
		Coeff[6077] <= 15'b100011001101110;
		Coeff[6078] <= 15'b100011001110000;
		Coeff[6079] <= 15'b100011001110011;
		Coeff[6080] <= 15'b100011001110101;
		Coeff[6081] <= 15'b100011001111000;
		Coeff[6082] <= 15'b100011001111011;
		Coeff[6083] <= 15'b100011001111101;
		Coeff[6084] <= 15'b100011010000000;
		Coeff[6085] <= 15'b100011010000011;
		Coeff[6086] <= 15'b100011010000101;
		Coeff[6087] <= 15'b100011010001000;
		Coeff[6088] <= 15'b100011010001010;
		Coeff[6089] <= 15'b100011010001101;
		Coeff[6090] <= 15'b100011010010000;
		Coeff[6091] <= 15'b100011010010010;
		Coeff[6092] <= 15'b100011010010101;
		Coeff[6093] <= 15'b100011010010111;
		Coeff[6094] <= 15'b100011010011010;
		Coeff[6095] <= 15'b100011010011101;
		Coeff[6096] <= 15'b100011010011111;
		Coeff[6097] <= 15'b100011010100010;
		Coeff[6098] <= 15'b100011010100101;
		Coeff[6099] <= 15'b100011010100111;
		Coeff[6100] <= 15'b100011010101010;
		Coeff[6101] <= 15'b100011010101100;
		Coeff[6102] <= 15'b100011010101111;
		Coeff[6103] <= 15'b100011010110010;
		Coeff[6104] <= 15'b100011010110100;
		Coeff[6105] <= 15'b100011010110111;
		Coeff[6106] <= 15'b100011010111010;
		Coeff[6107] <= 15'b100011010111100;
		Coeff[6108] <= 15'b100011010111111;
		Coeff[6109] <= 15'b100011011000001;
		Coeff[6110] <= 15'b100011011000100;
		Coeff[6111] <= 15'b100011011000111;
		Coeff[6112] <= 15'b100011011001001;
		Coeff[6113] <= 15'b100011011001100;
		Coeff[6114] <= 15'b100011011001110;
		Coeff[6115] <= 15'b100011011010001;
		Coeff[6116] <= 15'b100011011010100;
		Coeff[6117] <= 15'b100011011010110;
		Coeff[6118] <= 15'b100011011011001;
		Coeff[6119] <= 15'b100011011011100;
		Coeff[6120] <= 15'b100011011011110;
		Coeff[6121] <= 15'b100011011100001;
		Coeff[6122] <= 15'b100011011100011;
		Coeff[6123] <= 15'b100011011100110;
		Coeff[6124] <= 15'b100011011101001;
		Coeff[6125] <= 15'b100011011101011;
		Coeff[6126] <= 15'b100011011101110;
		Coeff[6127] <= 15'b100011011110000;
		Coeff[6128] <= 15'b100011011110011;
		Coeff[6129] <= 15'b100011011110110;
		Coeff[6130] <= 15'b100011011111000;
		Coeff[6131] <= 15'b100011011111011;
		Coeff[6132] <= 15'b100011011111110;
		Coeff[6133] <= 15'b100011100000000;
		Coeff[6134] <= 15'b100011100000011;
		Coeff[6135] <= 15'b100011100000101;
		Coeff[6136] <= 15'b100011100001000;
		Coeff[6137] <= 15'b100011100001011;
		Coeff[6138] <= 15'b100011100001101;
		Coeff[6139] <= 15'b100011100010000;
		Coeff[6140] <= 15'b100011100010010;
		Coeff[6141] <= 15'b100011100010101;
		Coeff[6142] <= 15'b100011100011000;
		Coeff[6143] <= 15'b100011100011010;
		Coeff[6144] <= 15'b100011100011101;
		Coeff[6145] <= 15'b100011100100000;
		Coeff[6146] <= 15'b100011100100010;
		Coeff[6147] <= 15'b100011100100101;
		Coeff[6148] <= 15'b100011100100111;
		Coeff[6149] <= 15'b100011100101010;
		Coeff[6150] <= 15'b100011100101101;
		Coeff[6151] <= 15'b100011100101111;
		Coeff[6152] <= 15'b100011100110010;
		Coeff[6153] <= 15'b100011100110100;
		Coeff[6154] <= 15'b100011100110111;
		Coeff[6155] <= 15'b100011100111010;
		Coeff[6156] <= 15'b100011100111100;
		Coeff[6157] <= 15'b100011100111111;
		Coeff[6158] <= 15'b100011101000001;
		Coeff[6159] <= 15'b100011101000100;
		Coeff[6160] <= 15'b100011101000111;
		Coeff[6161] <= 15'b100011101001001;
		Coeff[6162] <= 15'b100011101001100;
		Coeff[6163] <= 15'b100011101001111;
		Coeff[6164] <= 15'b100011101010001;
		Coeff[6165] <= 15'b100011101010100;
		Coeff[6166] <= 15'b100011101010110;
		Coeff[6167] <= 15'b100011101011001;
		Coeff[6168] <= 15'b100011101011100;
		Coeff[6169] <= 15'b100011101011110;
		Coeff[6170] <= 15'b100011101100001;
		Coeff[6171] <= 15'b100011101100011;
		Coeff[6172] <= 15'b100011101100110;
		Coeff[6173] <= 15'b100011101101001;
		Coeff[6174] <= 15'b100011101101011;
		Coeff[6175] <= 15'b100011101101110;
		Coeff[6176] <= 15'b100011101110000;
		Coeff[6177] <= 15'b100011101110011;
		Coeff[6178] <= 15'b100011101110110;
		Coeff[6179] <= 15'b100011101111000;
		Coeff[6180] <= 15'b100011101111011;
		Coeff[6181] <= 15'b100011101111101;
		Coeff[6182] <= 15'b100011110000000;
		Coeff[6183] <= 15'b100011110000011;
		Coeff[6184] <= 15'b100011110000101;
		Coeff[6185] <= 15'b100011110001000;
		Coeff[6186] <= 15'b100011110001010;
		Coeff[6187] <= 15'b100011110001101;
		Coeff[6188] <= 15'b100011110010000;
		Coeff[6189] <= 15'b100011110010010;
		Coeff[6190] <= 15'b100011110010101;
		Coeff[6191] <= 15'b100011110011000;
		Coeff[6192] <= 15'b100011110011010;
		Coeff[6193] <= 15'b100011110011101;
		Coeff[6194] <= 15'b100011110011111;
		Coeff[6195] <= 15'b100011110100010;
		Coeff[6196] <= 15'b100011110100101;
		Coeff[6197] <= 15'b100011110100111;
		Coeff[6198] <= 15'b100011110101010;
		Coeff[6199] <= 15'b100011110101100;
		Coeff[6200] <= 15'b100011110101111;
		Coeff[6201] <= 15'b100011110110010;
		Coeff[6202] <= 15'b100011110110100;
		Coeff[6203] <= 15'b100011110110111;
		Coeff[6204] <= 15'b100011110111001;
		Coeff[6205] <= 15'b100011110111100;
		Coeff[6206] <= 15'b100011110111111;
		Coeff[6207] <= 15'b100011111000001;
		Coeff[6208] <= 15'b100011111000100;
		Coeff[6209] <= 15'b100011111000110;
		Coeff[6210] <= 15'b100011111001001;
		Coeff[6211] <= 15'b100011111001100;
		Coeff[6212] <= 15'b100011111001110;
		Coeff[6213] <= 15'b100011111010001;
		Coeff[6214] <= 15'b100011111010011;
		Coeff[6215] <= 15'b100011111010110;
		Coeff[6216] <= 15'b100011111011001;
		Coeff[6217] <= 15'b100011111011011;
		Coeff[6218] <= 15'b100011111011110;
		Coeff[6219] <= 15'b100011111100000;
		Coeff[6220] <= 15'b100011111100011;
		Coeff[6221] <= 15'b100011111100110;
		Coeff[6222] <= 15'b100011111101000;
		Coeff[6223] <= 15'b100011111101011;
		Coeff[6224] <= 15'b100011111101101;
		Coeff[6225] <= 15'b100011111110000;
		Coeff[6226] <= 15'b100011111110011;
		Coeff[6227] <= 15'b100011111110101;
		Coeff[6228] <= 15'b100011111111000;
		Coeff[6229] <= 15'b100011111111010;
		Coeff[6230] <= 15'b100011111111101;
		Coeff[6231] <= 15'b100100000000000;
		Coeff[6232] <= 15'b100100000000010;
		Coeff[6233] <= 15'b100100000000101;
		Coeff[6234] <= 15'b100100000000111;
		Coeff[6235] <= 15'b100100000001010;
		Coeff[6236] <= 15'b100100000001101;
		Coeff[6237] <= 15'b100100000001111;
		Coeff[6238] <= 15'b100100000010010;
		Coeff[6239] <= 15'b100100000010100;
		Coeff[6240] <= 15'b100100000010111;
		Coeff[6241] <= 15'b100100000011010;
		Coeff[6242] <= 15'b100100000011100;
		Coeff[6243] <= 15'b100100000011111;
		Coeff[6244] <= 15'b100100000100001;
		Coeff[6245] <= 15'b100100000100100;
		Coeff[6246] <= 15'b100100000100110;
		Coeff[6247] <= 15'b100100000101001;
		Coeff[6248] <= 15'b100100000101100;
		Coeff[6249] <= 15'b100100000101110;
		Coeff[6250] <= 15'b100100000110001;
		Coeff[6251] <= 15'b100100000110011;
		Coeff[6252] <= 15'b100100000110110;
		Coeff[6253] <= 15'b100100000111001;
		Coeff[6254] <= 15'b100100000111011;
		Coeff[6255] <= 15'b100100000111110;
		Coeff[6256] <= 15'b100100001000000;
		Coeff[6257] <= 15'b100100001000011;
		Coeff[6258] <= 15'b100100001000110;
		Coeff[6259] <= 15'b100100001001000;
		Coeff[6260] <= 15'b100100001001011;
		Coeff[6261] <= 15'b100100001001101;
		Coeff[6262] <= 15'b100100001010000;
		Coeff[6263] <= 15'b100100001010011;
		Coeff[6264] <= 15'b100100001010101;
		Coeff[6265] <= 15'b100100001011000;
		Coeff[6266] <= 15'b100100001011010;
		Coeff[6267] <= 15'b100100001011101;
		Coeff[6268] <= 15'b100100001100000;
		Coeff[6269] <= 15'b100100001100010;
		Coeff[6270] <= 15'b100100001100101;
		Coeff[6271] <= 15'b100100001100111;
		Coeff[6272] <= 15'b100100001101010;
		Coeff[6273] <= 15'b100100001101100;
		Coeff[6274] <= 15'b100100001101111;
		Coeff[6275] <= 15'b100100001110010;
		Coeff[6276] <= 15'b100100001110100;
		Coeff[6277] <= 15'b100100001110111;
		Coeff[6278] <= 15'b100100001111001;
		Coeff[6279] <= 15'b100100001111100;
		Coeff[6280] <= 15'b100100001111111;
		Coeff[6281] <= 15'b100100010000001;
		Coeff[6282] <= 15'b100100010000100;
		Coeff[6283] <= 15'b100100010000110;
		Coeff[6284] <= 15'b100100010001001;
		Coeff[6285] <= 15'b100100010001100;
		Coeff[6286] <= 15'b100100010001110;
		Coeff[6287] <= 15'b100100010010001;
		Coeff[6288] <= 15'b100100010010011;
		Coeff[6289] <= 15'b100100010010110;
		Coeff[6290] <= 15'b100100010011001;
		Coeff[6291] <= 15'b100100010011011;
		Coeff[6292] <= 15'b100100010011110;
		Coeff[6293] <= 15'b100100010100000;
		Coeff[6294] <= 15'b100100010100011;
		Coeff[6295] <= 15'b100100010100101;
		Coeff[6296] <= 15'b100100010101000;
		Coeff[6297] <= 15'b100100010101011;
		Coeff[6298] <= 15'b100100010101101;
		Coeff[6299] <= 15'b100100010110000;
		Coeff[6300] <= 15'b100100010110010;
		Coeff[6301] <= 15'b100100010110101;
		Coeff[6302] <= 15'b100100010111000;
		Coeff[6303] <= 15'b100100010111010;
		Coeff[6304] <= 15'b100100010111101;
		Coeff[6305] <= 15'b100100010111111;
		Coeff[6306] <= 15'b100100011000010;
		Coeff[6307] <= 15'b100100011000100;
		Coeff[6308] <= 15'b100100011000111;
		Coeff[6309] <= 15'b100100011001010;
		Coeff[6310] <= 15'b100100011001100;
		Coeff[6311] <= 15'b100100011001111;
		Coeff[6312] <= 15'b100100011010001;
		Coeff[6313] <= 15'b100100011010100;
		Coeff[6314] <= 15'b100100011010111;
		Coeff[6315] <= 15'b100100011011001;
		Coeff[6316] <= 15'b100100011011100;
		Coeff[6317] <= 15'b100100011011110;
		Coeff[6318] <= 15'b100100011100001;
		Coeff[6319] <= 15'b100100011100011;
		Coeff[6320] <= 15'b100100011100110;
		Coeff[6321] <= 15'b100100011101001;
		Coeff[6322] <= 15'b100100011101011;
		Coeff[6323] <= 15'b100100011101110;
		Coeff[6324] <= 15'b100100011110000;
		Coeff[6325] <= 15'b100100011110011;
		Coeff[6326] <= 15'b100100011110110;
		Coeff[6327] <= 15'b100100011111000;
		Coeff[6328] <= 15'b100100011111011;
		Coeff[6329] <= 15'b100100011111101;
		Coeff[6330] <= 15'b100100100000000;
		Coeff[6331] <= 15'b100100100000010;
		Coeff[6332] <= 15'b100100100000101;
		Coeff[6333] <= 15'b100100100001000;
		Coeff[6334] <= 15'b100100100001010;
		Coeff[6335] <= 15'b100100100001101;
		Coeff[6336] <= 15'b100100100001111;
		Coeff[6337] <= 15'b100100100010010;
		Coeff[6338] <= 15'b100100100010101;
		Coeff[6339] <= 15'b100100100010111;
		Coeff[6340] <= 15'b100100100011010;
		Coeff[6341] <= 15'b100100100011100;
		Coeff[6342] <= 15'b100100100011111;
		Coeff[6343] <= 15'b100100100100001;
		Coeff[6344] <= 15'b100100100100100;
		Coeff[6345] <= 15'b100100100100111;
		Coeff[6346] <= 15'b100100100101001;
		Coeff[6347] <= 15'b100100100101100;
		Coeff[6348] <= 15'b100100100101110;
		Coeff[6349] <= 15'b100100100110001;
		Coeff[6350] <= 15'b100100100110011;
		Coeff[6351] <= 15'b100100100110110;
		Coeff[6352] <= 15'b100100100111001;
		Coeff[6353] <= 15'b100100100111011;
		Coeff[6354] <= 15'b100100100111110;
		Coeff[6355] <= 15'b100100101000000;
		Coeff[6356] <= 15'b100100101000011;
		Coeff[6357] <= 15'b100100101000101;
		Coeff[6358] <= 15'b100100101001000;
		Coeff[6359] <= 15'b100100101001011;
		Coeff[6360] <= 15'b100100101001101;
		Coeff[6361] <= 15'b100100101010000;
		Coeff[6362] <= 15'b100100101010010;
		Coeff[6363] <= 15'b100100101010101;
		Coeff[6364] <= 15'b100100101011000;
		Coeff[6365] <= 15'b100100101011010;
		Coeff[6366] <= 15'b100100101011101;
		Coeff[6367] <= 15'b100100101011111;
		Coeff[6368] <= 15'b100100101100010;
		Coeff[6369] <= 15'b100100101100100;
		Coeff[6370] <= 15'b100100101100111;
		Coeff[6371] <= 15'b100100101101010;
		Coeff[6372] <= 15'b100100101101100;
		Coeff[6373] <= 15'b100100101101111;
		Coeff[6374] <= 15'b100100101110001;
		Coeff[6375] <= 15'b100100101110100;
		Coeff[6376] <= 15'b100100101110110;
		Coeff[6377] <= 15'b100100101111001;
		Coeff[6378] <= 15'b100100101111100;
		Coeff[6379] <= 15'b100100101111110;
		Coeff[6380] <= 15'b100100110000001;
		Coeff[6381] <= 15'b100100110000011;
		Coeff[6382] <= 15'b100100110000110;
		Coeff[6383] <= 15'b100100110001000;
		Coeff[6384] <= 15'b100100110001011;
		Coeff[6385] <= 15'b100100110001110;
		Coeff[6386] <= 15'b100100110010000;
		Coeff[6387] <= 15'b100100110010011;
		Coeff[6388] <= 15'b100100110010101;
		Coeff[6389] <= 15'b100100110011000;
		Coeff[6390] <= 15'b100100110011010;
		Coeff[6391] <= 15'b100100110011101;
		Coeff[6392] <= 15'b100100110100000;
		Coeff[6393] <= 15'b100100110100010;
		Coeff[6394] <= 15'b100100110100101;
		Coeff[6395] <= 15'b100100110100111;
		Coeff[6396] <= 15'b100100110101010;
		Coeff[6397] <= 15'b100100110101100;
		Coeff[6398] <= 15'b100100110101111;
		Coeff[6399] <= 15'b100100110110010;
		Coeff[6400] <= 15'b100100110110100;
		Coeff[6401] <= 15'b100100110110111;
		Coeff[6402] <= 15'b100100110111001;
		Coeff[6403] <= 15'b100100110111100;
		Coeff[6404] <= 15'b100100110111110;
		Coeff[6405] <= 15'b100100111000001;
		Coeff[6406] <= 15'b100100111000011;
		Coeff[6407] <= 15'b100100111000110;
		Coeff[6408] <= 15'b100100111001001;
		Coeff[6409] <= 15'b100100111001011;
		Coeff[6410] <= 15'b100100111001110;
		Coeff[6411] <= 15'b100100111010000;
		Coeff[6412] <= 15'b100100111010011;
		Coeff[6413] <= 15'b100100111010101;
		Coeff[6414] <= 15'b100100111011000;
		Coeff[6415] <= 15'b100100111011011;
		Coeff[6416] <= 15'b100100111011101;
		Coeff[6417] <= 15'b100100111100000;
		Coeff[6418] <= 15'b100100111100010;
		Coeff[6419] <= 15'b100100111100101;
		Coeff[6420] <= 15'b100100111100111;
		Coeff[6421] <= 15'b100100111101010;
		Coeff[6422] <= 15'b100100111101101;
		Coeff[6423] <= 15'b100100111101111;
		Coeff[6424] <= 15'b100100111110010;
		Coeff[6425] <= 15'b100100111110100;
		Coeff[6426] <= 15'b100100111110111;
		Coeff[6427] <= 15'b100100111111001;
		Coeff[6428] <= 15'b100100111111100;
		Coeff[6429] <= 15'b100100111111110;
		Coeff[6430] <= 15'b100101000000001;
		Coeff[6431] <= 15'b100101000000100;
		Coeff[6432] <= 15'b100101000000110;
		Coeff[6433] <= 15'b100101000001001;
		Coeff[6434] <= 15'b100101000001011;
		Coeff[6435] <= 15'b100101000001110;
		Coeff[6436] <= 15'b100101000010000;
		Coeff[6437] <= 15'b100101000010011;
		Coeff[6438] <= 15'b100101000010110;
		Coeff[6439] <= 15'b100101000011000;
		Coeff[6440] <= 15'b100101000011011;
		Coeff[6441] <= 15'b100101000011101;
		Coeff[6442] <= 15'b100101000100000;
		Coeff[6443] <= 15'b100101000100010;
		Coeff[6444] <= 15'b100101000100101;
		Coeff[6445] <= 15'b100101000100111;
		Coeff[6446] <= 15'b100101000101010;
		Coeff[6447] <= 15'b100101000101101;
		Coeff[6448] <= 15'b100101000101111;
		Coeff[6449] <= 15'b100101000110010;
		Coeff[6450] <= 15'b100101000110100;
		Coeff[6451] <= 15'b100101000110111;
		Coeff[6452] <= 15'b100101000111001;
		Coeff[6453] <= 15'b100101000111100;
		Coeff[6454] <= 15'b100101000111111;
		Coeff[6455] <= 15'b100101001000001;
		Coeff[6456] <= 15'b100101001000100;
		Coeff[6457] <= 15'b100101001000110;
		Coeff[6458] <= 15'b100101001001001;
		Coeff[6459] <= 15'b100101001001011;
		Coeff[6460] <= 15'b100101001001110;
		Coeff[6461] <= 15'b100101001010000;
		Coeff[6462] <= 15'b100101001010011;
		Coeff[6463] <= 15'b100101001010110;
		Coeff[6464] <= 15'b100101001011000;
		Coeff[6465] <= 15'b100101001011011;
		Coeff[6466] <= 15'b100101001011101;
		Coeff[6467] <= 15'b100101001100000;
		Coeff[6468] <= 15'b100101001100010;
		Coeff[6469] <= 15'b100101001100101;
		Coeff[6470] <= 15'b100101001100111;
		Coeff[6471] <= 15'b100101001101010;
		Coeff[6472] <= 15'b100101001101101;
		Coeff[6473] <= 15'b100101001101111;
		Coeff[6474] <= 15'b100101001110010;
		Coeff[6475] <= 15'b100101001110100;
		Coeff[6476] <= 15'b100101001110111;
		Coeff[6477] <= 15'b100101001111001;
		Coeff[6478] <= 15'b100101001111100;
		Coeff[6479] <= 15'b100101001111110;
		Coeff[6480] <= 15'b100101010000001;
		Coeff[6481] <= 15'b100101010000100;
		Coeff[6482] <= 15'b100101010000110;
		Coeff[6483] <= 15'b100101010001001;
		Coeff[6484] <= 15'b100101010001011;
		Coeff[6485] <= 15'b100101010001110;
		Coeff[6486] <= 15'b100101010010000;
		Coeff[6487] <= 15'b100101010010011;
		Coeff[6488] <= 15'b100101010010101;
		Coeff[6489] <= 15'b100101010011000;
		Coeff[6490] <= 15'b100101010011011;
		Coeff[6491] <= 15'b100101010011101;
		Coeff[6492] <= 15'b100101010100000;
		Coeff[6493] <= 15'b100101010100010;
		Coeff[6494] <= 15'b100101010100101;
		Coeff[6495] <= 15'b100101010100111;
		Coeff[6496] <= 15'b100101010101010;
		Coeff[6497] <= 15'b100101010101100;
		Coeff[6498] <= 15'b100101010101111;
		Coeff[6499] <= 15'b100101010110010;
		Coeff[6500] <= 15'b100101010110100;
		Coeff[6501] <= 15'b100101010110111;
		Coeff[6502] <= 15'b100101010111001;
		Coeff[6503] <= 15'b100101010111100;
		Coeff[6504] <= 15'b100101010111110;
		Coeff[6505] <= 15'b100101011000001;
		Coeff[6506] <= 15'b100101011000011;
		Coeff[6507] <= 15'b100101011000110;
		Coeff[6508] <= 15'b100101011001000;
		Coeff[6509] <= 15'b100101011001011;
		Coeff[6510] <= 15'b100101011001110;
		Coeff[6511] <= 15'b100101011010000;
		Coeff[6512] <= 15'b100101011010011;
		Coeff[6513] <= 15'b100101011010101;
		Coeff[6514] <= 15'b100101011011000;
		Coeff[6515] <= 15'b100101011011010;
		Coeff[6516] <= 15'b100101011011101;
		Coeff[6517] <= 15'b100101011011111;
		Coeff[6518] <= 15'b100101011100010;
		Coeff[6519] <= 15'b100101011100101;
		Coeff[6520] <= 15'b100101011100111;
		Coeff[6521] <= 15'b100101011101010;
		Coeff[6522] <= 15'b100101011101100;
		Coeff[6523] <= 15'b100101011101111;
		Coeff[6524] <= 15'b100101011110001;
		Coeff[6525] <= 15'b100101011110100;
		Coeff[6526] <= 15'b100101011110110;
		Coeff[6527] <= 15'b100101011111001;
		Coeff[6528] <= 15'b100101011111011;
		Coeff[6529] <= 15'b100101011111110;
		Coeff[6530] <= 15'b100101100000001;
		Coeff[6531] <= 15'b100101100000011;
		Coeff[6532] <= 15'b100101100000110;
		Coeff[6533] <= 15'b100101100001000;
		Coeff[6534] <= 15'b100101100001011;
		Coeff[6535] <= 15'b100101100001101;
		Coeff[6536] <= 15'b100101100010000;
		Coeff[6537] <= 15'b100101100010010;
		Coeff[6538] <= 15'b100101100010101;
		Coeff[6539] <= 15'b100101100010111;
		Coeff[6540] <= 15'b100101100011010;
		Coeff[6541] <= 15'b100101100011101;
		Coeff[6542] <= 15'b100101100011111;
		Coeff[6543] <= 15'b100101100100010;
		Coeff[6544] <= 15'b100101100100100;
		Coeff[6545] <= 15'b100101100100111;
		Coeff[6546] <= 15'b100101100101001;
		Coeff[6547] <= 15'b100101100101100;
		Coeff[6548] <= 15'b100101100101110;
		Coeff[6549] <= 15'b100101100110001;
		Coeff[6550] <= 15'b100101100110011;
		Coeff[6551] <= 15'b100101100110110;
		Coeff[6552] <= 15'b100101100111000;
		Coeff[6553] <= 15'b100101100111011;
		Coeff[6554] <= 15'b100101100111110;
		Coeff[6555] <= 15'b100101101000000;
		Coeff[6556] <= 15'b100101101000011;
		Coeff[6557] <= 15'b100101101000101;
		Coeff[6558] <= 15'b100101101001000;
		Coeff[6559] <= 15'b100101101001010;
		Coeff[6560] <= 15'b100101101001101;
		Coeff[6561] <= 15'b100101101001111;
		Coeff[6562] <= 15'b100101101010010;
		Coeff[6563] <= 15'b100101101010100;
		Coeff[6564] <= 15'b100101101010111;
		Coeff[6565] <= 15'b100101101011010;
		Coeff[6566] <= 15'b100101101011100;
		Coeff[6567] <= 15'b100101101011111;
		Coeff[6568] <= 15'b100101101100001;
		Coeff[6569] <= 15'b100101101100100;
		Coeff[6570] <= 15'b100101101100110;
		Coeff[6571] <= 15'b100101101101001;
		Coeff[6572] <= 15'b100101101101011;
		Coeff[6573] <= 15'b100101101101110;
		Coeff[6574] <= 15'b100101101110000;
		Coeff[6575] <= 15'b100101101110011;
		Coeff[6576] <= 15'b100101101110101;
		Coeff[6577] <= 15'b100101101111000;
		Coeff[6578] <= 15'b100101101111011;
		Coeff[6579] <= 15'b100101101111101;
		Coeff[6580] <= 15'b100101110000000;
		Coeff[6581] <= 15'b100101110000010;
		Coeff[6582] <= 15'b100101110000101;
		Coeff[6583] <= 15'b100101110000111;
		Coeff[6584] <= 15'b100101110001010;
		Coeff[6585] <= 15'b100101110001100;
		Coeff[6586] <= 15'b100101110001111;
		Coeff[6587] <= 15'b100101110010001;
		Coeff[6588] <= 15'b100101110010100;
		Coeff[6589] <= 15'b100101110010110;
		Coeff[6590] <= 15'b100101110011001;
		Coeff[6591] <= 15'b100101110011011;
		Coeff[6592] <= 15'b100101110011110;
		Coeff[6593] <= 15'b100101110100001;
		Coeff[6594] <= 15'b100101110100011;
		Coeff[6595] <= 15'b100101110100110;
		Coeff[6596] <= 15'b100101110101000;
		Coeff[6597] <= 15'b100101110101011;
		Coeff[6598] <= 15'b100101110101101;
		Coeff[6599] <= 15'b100101110110000;
		Coeff[6600] <= 15'b100101110110010;
		Coeff[6601] <= 15'b100101110110101;
		Coeff[6602] <= 15'b100101110110111;
		Coeff[6603] <= 15'b100101110111010;
		Coeff[6604] <= 15'b100101110111100;
		Coeff[6605] <= 15'b100101110111111;
		Coeff[6606] <= 15'b100101111000001;
		Coeff[6607] <= 15'b100101111000100;
		Coeff[6608] <= 15'b100101111000111;
		Coeff[6609] <= 15'b100101111001001;
		Coeff[6610] <= 15'b100101111001100;
		Coeff[6611] <= 15'b100101111001110;
		Coeff[6612] <= 15'b100101111010001;
		Coeff[6613] <= 15'b100101111010011;
		Coeff[6614] <= 15'b100101111010110;
		Coeff[6615] <= 15'b100101111011000;
		Coeff[6616] <= 15'b100101111011011;
		Coeff[6617] <= 15'b100101111011101;
		Coeff[6618] <= 15'b100101111100000;
		Coeff[6619] <= 15'b100101111100010;
		Coeff[6620] <= 15'b100101111100101;
		Coeff[6621] <= 15'b100101111100111;
		Coeff[6622] <= 15'b100101111101010;
		Coeff[6623] <= 15'b100101111101101;
		Coeff[6624] <= 15'b100101111101111;
		Coeff[6625] <= 15'b100101111110010;
		Coeff[6626] <= 15'b100101111110100;
		Coeff[6627] <= 15'b100101111110111;
		Coeff[6628] <= 15'b100101111111001;
		Coeff[6629] <= 15'b100101111111100;
		Coeff[6630] <= 15'b100101111111110;
		Coeff[6631] <= 15'b100110000000001;
		Coeff[6632] <= 15'b100110000000011;
		Coeff[6633] <= 15'b100110000000110;
		Coeff[6634] <= 15'b100110000001000;
		Coeff[6635] <= 15'b100110000001011;
		Coeff[6636] <= 15'b100110000001101;
		Coeff[6637] <= 15'b100110000010000;
		Coeff[6638] <= 15'b100110000010010;
		Coeff[6639] <= 15'b100110000010101;
		Coeff[6640] <= 15'b100110000010111;
		Coeff[6641] <= 15'b100110000011010;
		Coeff[6642] <= 15'b100110000011101;
		Coeff[6643] <= 15'b100110000011111;
		Coeff[6644] <= 15'b100110000100010;
		Coeff[6645] <= 15'b100110000100100;
		Coeff[6646] <= 15'b100110000100111;
		Coeff[6647] <= 15'b100110000101001;
		Coeff[6648] <= 15'b100110000101100;
		Coeff[6649] <= 15'b100110000101110;
		Coeff[6650] <= 15'b100110000110001;
		Coeff[6651] <= 15'b100110000110011;
		Coeff[6652] <= 15'b100110000110110;
		Coeff[6653] <= 15'b100110000111000;
		Coeff[6654] <= 15'b100110000111011;
		Coeff[6655] <= 15'b100110000111101;
		Coeff[6656] <= 15'b100110001000000;
		Coeff[6657] <= 15'b100110001000010;
		Coeff[6658] <= 15'b100110001000101;
		Coeff[6659] <= 15'b100110001000111;
		Coeff[6660] <= 15'b100110001001010;
		Coeff[6661] <= 15'b100110001001100;
		Coeff[6662] <= 15'b100110001001111;
		Coeff[6663] <= 15'b100110001010010;
		Coeff[6664] <= 15'b100110001010100;
		Coeff[6665] <= 15'b100110001010111;
		Coeff[6666] <= 15'b100110001011001;
		Coeff[6667] <= 15'b100110001011100;
		Coeff[6668] <= 15'b100110001011110;
		Coeff[6669] <= 15'b100110001100001;
		Coeff[6670] <= 15'b100110001100011;
		Coeff[6671] <= 15'b100110001100110;
		Coeff[6672] <= 15'b100110001101000;
		Coeff[6673] <= 15'b100110001101011;
		Coeff[6674] <= 15'b100110001101101;
		Coeff[6675] <= 15'b100110001110000;
		Coeff[6676] <= 15'b100110001110010;
		Coeff[6677] <= 15'b100110001110101;
		Coeff[6678] <= 15'b100110001110111;
		Coeff[6679] <= 15'b100110001111010;
		Coeff[6680] <= 15'b100110001111100;
		Coeff[6681] <= 15'b100110001111111;
		Coeff[6682] <= 15'b100110010000001;
		Coeff[6683] <= 15'b100110010000100;
		Coeff[6684] <= 15'b100110010000110;
		Coeff[6685] <= 15'b100110010001001;
		Coeff[6686] <= 15'b100110010001011;
		Coeff[6687] <= 15'b100110010001110;
		Coeff[6688] <= 15'b100110010010001;
		Coeff[6689] <= 15'b100110010010011;
		Coeff[6690] <= 15'b100110010010110;
		Coeff[6691] <= 15'b100110010011000;
		Coeff[6692] <= 15'b100110010011011;
		Coeff[6693] <= 15'b100110010011101;
		Coeff[6694] <= 15'b100110010100000;
		Coeff[6695] <= 15'b100110010100010;
		Coeff[6696] <= 15'b100110010100101;
		Coeff[6697] <= 15'b100110010100111;
		Coeff[6698] <= 15'b100110010101010;
		Coeff[6699] <= 15'b100110010101100;
		Coeff[6700] <= 15'b100110010101111;
		Coeff[6701] <= 15'b100110010110001;
		Coeff[6702] <= 15'b100110010110100;
		Coeff[6703] <= 15'b100110010110110;
		Coeff[6704] <= 15'b100110010111001;
		Coeff[6705] <= 15'b100110010111011;
		Coeff[6706] <= 15'b100110010111110;
		Coeff[6707] <= 15'b100110011000000;
		Coeff[6708] <= 15'b100110011000011;
		Coeff[6709] <= 15'b100110011000101;
		Coeff[6710] <= 15'b100110011001000;
		Coeff[6711] <= 15'b100110011001010;
		Coeff[6712] <= 15'b100110011001101;
		Coeff[6713] <= 15'b100110011001111;
		Coeff[6714] <= 15'b100110011010010;
		Coeff[6715] <= 15'b100110011010100;
		Coeff[6716] <= 15'b100110011010111;
		Coeff[6717] <= 15'b100110011011001;
		Coeff[6718] <= 15'b100110011011100;
		Coeff[6719] <= 15'b100110011011110;
		Coeff[6720] <= 15'b100110011100001;
		Coeff[6721] <= 15'b100110011100100;
		Coeff[6722] <= 15'b100110011100110;
		Coeff[6723] <= 15'b100110011101001;
		Coeff[6724] <= 15'b100110011101011;
		Coeff[6725] <= 15'b100110011101110;
		Coeff[6726] <= 15'b100110011110000;
		Coeff[6727] <= 15'b100110011110011;
		Coeff[6728] <= 15'b100110011110101;
		Coeff[6729] <= 15'b100110011111000;
		Coeff[6730] <= 15'b100110011111010;
		Coeff[6731] <= 15'b100110011111101;
		Coeff[6732] <= 15'b100110011111111;
		Coeff[6733] <= 15'b100110100000010;
		Coeff[6734] <= 15'b100110100000100;
		Coeff[6735] <= 15'b100110100000111;
		Coeff[6736] <= 15'b100110100001001;
		Coeff[6737] <= 15'b100110100001100;
		Coeff[6738] <= 15'b100110100001110;
		Coeff[6739] <= 15'b100110100010001;
		Coeff[6740] <= 15'b100110100010011;
		Coeff[6741] <= 15'b100110100010110;
		Coeff[6742] <= 15'b100110100011000;
		Coeff[6743] <= 15'b100110100011011;
		Coeff[6744] <= 15'b100110100011101;
		Coeff[6745] <= 15'b100110100100000;
		Coeff[6746] <= 15'b100110100100010;
		Coeff[6747] <= 15'b100110100100101;
		Coeff[6748] <= 15'b100110100100111;
		Coeff[6749] <= 15'b100110100101010;
		Coeff[6750] <= 15'b100110100101100;
		Coeff[6751] <= 15'b100110100101111;
		Coeff[6752] <= 15'b100110100110001;
		Coeff[6753] <= 15'b100110100110100;
		Coeff[6754] <= 15'b100110100110110;
		Coeff[6755] <= 15'b100110100111001;
		Coeff[6756] <= 15'b100110100111011;
		Coeff[6757] <= 15'b100110100111110;
		Coeff[6758] <= 15'b100110101000000;
		Coeff[6759] <= 15'b100110101000011;
		Coeff[6760] <= 15'b100110101000101;
		Coeff[6761] <= 15'b100110101001000;
		Coeff[6762] <= 15'b100110101001010;
		Coeff[6763] <= 15'b100110101001101;
		Coeff[6764] <= 15'b100110101001111;
		Coeff[6765] <= 15'b100110101010010;
		Coeff[6766] <= 15'b100110101010100;
		Coeff[6767] <= 15'b100110101010111;
		Coeff[6768] <= 15'b100110101011001;
		Coeff[6769] <= 15'b100110101011100;
		Coeff[6770] <= 15'b100110101011110;
		Coeff[6771] <= 15'b100110101100001;
		Coeff[6772] <= 15'b100110101100011;
		Coeff[6773] <= 15'b100110101100110;
		Coeff[6774] <= 15'b100110101101000;
		Coeff[6775] <= 15'b100110101101011;
		Coeff[6776] <= 15'b100110101101101;
		Coeff[6777] <= 15'b100110101110000;
		Coeff[6778] <= 15'b100110101110010;
		Coeff[6779] <= 15'b100110101110101;
		Coeff[6780] <= 15'b100110101110111;
		Coeff[6781] <= 15'b100110101111010;
		Coeff[6782] <= 15'b100110101111100;
		Coeff[6783] <= 15'b100110101111111;
		Coeff[6784] <= 15'b100110110000001;
		Coeff[6785] <= 15'b100110110000100;
		Coeff[6786] <= 15'b100110110000110;
		Coeff[6787] <= 15'b100110110001001;
		Coeff[6788] <= 15'b100110110001011;
		Coeff[6789] <= 15'b100110110001110;
		Coeff[6790] <= 15'b100110110010000;
		Coeff[6791] <= 15'b100110110010011;
		Coeff[6792] <= 15'b100110110010101;
		Coeff[6793] <= 15'b100110110011000;
		Coeff[6794] <= 15'b100110110011010;
		Coeff[6795] <= 15'b100110110011101;
		Coeff[6796] <= 15'b100110110011111;
		Coeff[6797] <= 15'b100110110100010;
		Coeff[6798] <= 15'b100110110100100;
		Coeff[6799] <= 15'b100110110100111;
		Coeff[6800] <= 15'b100110110101001;
		Coeff[6801] <= 15'b100110110101100;
		Coeff[6802] <= 15'b100110110101110;
		Coeff[6803] <= 15'b100110110110001;
		Coeff[6804] <= 15'b100110110110011;
		Coeff[6805] <= 15'b100110110110110;
		Coeff[6806] <= 15'b100110110111000;
		Coeff[6807] <= 15'b100110110111011;
		Coeff[6808] <= 15'b100110110111101;
		Coeff[6809] <= 15'b100110111000000;
		Coeff[6810] <= 15'b100110111000010;
		Coeff[6811] <= 15'b100110111000101;
		Coeff[6812] <= 15'b100110111000111;
		Coeff[6813] <= 15'b100110111001010;
		Coeff[6814] <= 15'b100110111001100;
		Coeff[6815] <= 15'b100110111001111;
		Coeff[6816] <= 15'b100110111010001;
		Coeff[6817] <= 15'b100110111010100;
		Coeff[6818] <= 15'b100110111010110;
		Coeff[6819] <= 15'b100110111011001;
		Coeff[6820] <= 15'b100110111011011;
		Coeff[6821] <= 15'b100110111011110;
		Coeff[6822] <= 15'b100110111100000;
		Coeff[6823] <= 15'b100110111100011;
		Coeff[6824] <= 15'b100110111100101;
		Coeff[6825] <= 15'b100110111101000;
		Coeff[6826] <= 15'b100110111101010;
		Coeff[6827] <= 15'b100110111101101;
		Coeff[6828] <= 15'b100110111101111;
		Coeff[6829] <= 15'b100110111110010;
		Coeff[6830] <= 15'b100110111110100;
		Coeff[6831] <= 15'b100110111110111;
		Coeff[6832] <= 15'b100110111111001;
		Coeff[6833] <= 15'b100110111111100;
		Coeff[6834] <= 15'b100110111111110;
		Coeff[6835] <= 15'b100111000000001;
		Coeff[6836] <= 15'b100111000000011;
		Coeff[6837] <= 15'b100111000000110;
		Coeff[6838] <= 15'b100111000001000;
		Coeff[6839] <= 15'b100111000001011;
		Coeff[6840] <= 15'b100111000001101;
		Coeff[6841] <= 15'b100111000010000;
		Coeff[6842] <= 15'b100111000010010;
		Coeff[6843] <= 15'b100111000010101;
		Coeff[6844] <= 15'b100111000010111;
		Coeff[6845] <= 15'b100111000011010;
		Coeff[6846] <= 15'b100111000011100;
		Coeff[6847] <= 15'b100111000011111;
		Coeff[6848] <= 15'b100111000100001;
		Coeff[6849] <= 15'b100111000100100;
		Coeff[6850] <= 15'b100111000100110;
		Coeff[6851] <= 15'b100111000101000;
		Coeff[6852] <= 15'b100111000101011;
		Coeff[6853] <= 15'b100111000101101;
		Coeff[6854] <= 15'b100111000110000;
		Coeff[6855] <= 15'b100111000110010;
		Coeff[6856] <= 15'b100111000110101;
		Coeff[6857] <= 15'b100111000110111;
		Coeff[6858] <= 15'b100111000111010;
		Coeff[6859] <= 15'b100111000111100;
		Coeff[6860] <= 15'b100111000111111;
		Coeff[6861] <= 15'b100111001000001;
		Coeff[6862] <= 15'b100111001000100;
		Coeff[6863] <= 15'b100111001000110;
		Coeff[6864] <= 15'b100111001001001;
		Coeff[6865] <= 15'b100111001001011;
		Coeff[6866] <= 15'b100111001001110;
		Coeff[6867] <= 15'b100111001010000;
		Coeff[6868] <= 15'b100111001010011;
		Coeff[6869] <= 15'b100111001010101;
		Coeff[6870] <= 15'b100111001011000;
		Coeff[6871] <= 15'b100111001011010;
		Coeff[6872] <= 15'b100111001011101;
		Coeff[6873] <= 15'b100111001011111;
		Coeff[6874] <= 15'b100111001100010;
		Coeff[6875] <= 15'b100111001100100;
		Coeff[6876] <= 15'b100111001100111;
		Coeff[6877] <= 15'b100111001101001;
		Coeff[6878] <= 15'b100111001101100;
		Coeff[6879] <= 15'b100111001101110;
		Coeff[6880] <= 15'b100111001110001;
		Coeff[6881] <= 15'b100111001110011;
		Coeff[6882] <= 15'b100111001110110;
		Coeff[6883] <= 15'b100111001111000;
		Coeff[6884] <= 15'b100111001111010;
		Coeff[6885] <= 15'b100111001111101;
		Coeff[6886] <= 15'b100111001111111;
		Coeff[6887] <= 15'b100111010000010;
		Coeff[6888] <= 15'b100111010000100;
		Coeff[6889] <= 15'b100111010000111;
		Coeff[6890] <= 15'b100111010001001;
		Coeff[6891] <= 15'b100111010001100;
		Coeff[6892] <= 15'b100111010001110;
		Coeff[6893] <= 15'b100111010010001;
		Coeff[6894] <= 15'b100111010010011;
		Coeff[6895] <= 15'b100111010010110;
		Coeff[6896] <= 15'b100111010011000;
		Coeff[6897] <= 15'b100111010011011;
		Coeff[6898] <= 15'b100111010011101;
		Coeff[6899] <= 15'b100111010100000;
		Coeff[6900] <= 15'b100111010100010;
		Coeff[6901] <= 15'b100111010100101;
		Coeff[6902] <= 15'b100111010100111;
		Coeff[6903] <= 15'b100111010101010;
		Coeff[6904] <= 15'b100111010101100;
		Coeff[6905] <= 15'b100111010101111;
		Coeff[6906] <= 15'b100111010110001;
		Coeff[6907] <= 15'b100111010110100;
		Coeff[6908] <= 15'b100111010110110;
		Coeff[6909] <= 15'b100111010111000;
		Coeff[6910] <= 15'b100111010111011;
		Coeff[6911] <= 15'b100111010111101;
		Coeff[6912] <= 15'b100111011000000;
		Coeff[6913] <= 15'b100111011000010;
		Coeff[6914] <= 15'b100111011000101;
		Coeff[6915] <= 15'b100111011000111;
		Coeff[6916] <= 15'b100111011001010;
		Coeff[6917] <= 15'b100111011001100;
		Coeff[6918] <= 15'b100111011001111;
		Coeff[6919] <= 15'b100111011010001;
		Coeff[6920] <= 15'b100111011010100;
		Coeff[6921] <= 15'b100111011010110;
		Coeff[6922] <= 15'b100111011011001;
		Coeff[6923] <= 15'b100111011011011;
		Coeff[6924] <= 15'b100111011011110;
		Coeff[6925] <= 15'b100111011100000;
		Coeff[6926] <= 15'b100111011100011;
		Coeff[6927] <= 15'b100111011100101;
		Coeff[6928] <= 15'b100111011101000;
		Coeff[6929] <= 15'b100111011101010;
		Coeff[6930] <= 15'b100111011101100;
		Coeff[6931] <= 15'b100111011101111;
		Coeff[6932] <= 15'b100111011110001;
		Coeff[6933] <= 15'b100111011110100;
		Coeff[6934] <= 15'b100111011110110;
		Coeff[6935] <= 15'b100111011111001;
		Coeff[6936] <= 15'b100111011111011;
		Coeff[6937] <= 15'b100111011111110;
		Coeff[6938] <= 15'b100111100000000;
		Coeff[6939] <= 15'b100111100000011;
		Coeff[6940] <= 15'b100111100000101;
		Coeff[6941] <= 15'b100111100001000;
		Coeff[6942] <= 15'b100111100001010;
		Coeff[6943] <= 15'b100111100001101;
		Coeff[6944] <= 15'b100111100001111;
		Coeff[6945] <= 15'b100111100010010;
		Coeff[6946] <= 15'b100111100010100;
		Coeff[6947] <= 15'b100111100010110;
		Coeff[6948] <= 15'b100111100011001;
		Coeff[6949] <= 15'b100111100011011;
		Coeff[6950] <= 15'b100111100011110;
		Coeff[6951] <= 15'b100111100100000;
		Coeff[6952] <= 15'b100111100100011;
		Coeff[6953] <= 15'b100111100100101;
		Coeff[6954] <= 15'b100111100101000;
		Coeff[6955] <= 15'b100111100101010;
		Coeff[6956] <= 15'b100111100101101;
		Coeff[6957] <= 15'b100111100101111;
		Coeff[6958] <= 15'b100111100110010;
		Coeff[6959] <= 15'b100111100110100;
		Coeff[6960] <= 15'b100111100110111;
		Coeff[6961] <= 15'b100111100111001;
		Coeff[6962] <= 15'b100111100111100;
		Coeff[6963] <= 15'b100111100111110;
		Coeff[6964] <= 15'b100111101000000;
		Coeff[6965] <= 15'b100111101000011;
		Coeff[6966] <= 15'b100111101000101;
		Coeff[6967] <= 15'b100111101001000;
		Coeff[6968] <= 15'b100111101001010;
		Coeff[6969] <= 15'b100111101001101;
		Coeff[6970] <= 15'b100111101001111;
		Coeff[6971] <= 15'b100111101010010;
		Coeff[6972] <= 15'b100111101010100;
		Coeff[6973] <= 15'b100111101010111;
		Coeff[6974] <= 15'b100111101011001;
		Coeff[6975] <= 15'b100111101011100;
		Coeff[6976] <= 15'b100111101011110;
		Coeff[6977] <= 15'b100111101100000;
		Coeff[6978] <= 15'b100111101100011;
		Coeff[6979] <= 15'b100111101100101;
		Coeff[6980] <= 15'b100111101101000;
		Coeff[6981] <= 15'b100111101101010;
		Coeff[6982] <= 15'b100111101101101;
		Coeff[6983] <= 15'b100111101101111;
		Coeff[6984] <= 15'b100111101110010;
		Coeff[6985] <= 15'b100111101110100;
		Coeff[6986] <= 15'b100111101110111;
		Coeff[6987] <= 15'b100111101111001;
		Coeff[6988] <= 15'b100111101111100;
		Coeff[6989] <= 15'b100111101111110;
		Coeff[6990] <= 15'b100111110000001;
		Coeff[6991] <= 15'b100111110000011;
		Coeff[6992] <= 15'b100111110000101;
		Coeff[6993] <= 15'b100111110001000;
		Coeff[6994] <= 15'b100111110001010;
		Coeff[6995] <= 15'b100111110001101;
		Coeff[6996] <= 15'b100111110001111;
		Coeff[6997] <= 15'b100111110010010;
		Coeff[6998] <= 15'b100111110010100;
		Coeff[6999] <= 15'b100111110010111;
		Coeff[7000] <= 15'b100111110011001;
		Coeff[7001] <= 15'b100111110011100;
		Coeff[7002] <= 15'b100111110011110;
		Coeff[7003] <= 15'b100111110100001;
		Coeff[7004] <= 15'b100111110100011;
		Coeff[7005] <= 15'b100111110100101;
		Coeff[7006] <= 15'b100111110101000;
		Coeff[7007] <= 15'b100111110101010;
		Coeff[7008] <= 15'b100111110101101;
		Coeff[7009] <= 15'b100111110101111;
		Coeff[7010] <= 15'b100111110110010;
		Coeff[7011] <= 15'b100111110110100;
		Coeff[7012] <= 15'b100111110110111;
		Coeff[7013] <= 15'b100111110111001;
		Coeff[7014] <= 15'b100111110111100;
		Coeff[7015] <= 15'b100111110111110;
		Coeff[7016] <= 15'b100111111000000;
		Coeff[7017] <= 15'b100111111000011;
		Coeff[7018] <= 15'b100111111000101;
		Coeff[7019] <= 15'b100111111001000;
		Coeff[7020] <= 15'b100111111001010;
		Coeff[7021] <= 15'b100111111001101;
		Coeff[7022] <= 15'b100111111001111;
		Coeff[7023] <= 15'b100111111010010;
		Coeff[7024] <= 15'b100111111010100;
		Coeff[7025] <= 15'b100111111010111;
		Coeff[7026] <= 15'b100111111011001;
		Coeff[7027] <= 15'b100111111011011;
		Coeff[7028] <= 15'b100111111011110;
		Coeff[7029] <= 15'b100111111100000;
		Coeff[7030] <= 15'b100111111100011;
		Coeff[7031] <= 15'b100111111100101;
		Coeff[7032] <= 15'b100111111101000;
		Coeff[7033] <= 15'b100111111101010;
		Coeff[7034] <= 15'b100111111101101;
		Coeff[7035] <= 15'b100111111101111;
		Coeff[7036] <= 15'b100111111110010;
		Coeff[7037] <= 15'b100111111110100;
		Coeff[7038] <= 15'b100111111110110;
		Coeff[7039] <= 15'b100111111111001;
		Coeff[7040] <= 15'b100111111111011;
		Coeff[7041] <= 15'b100111111111110;
		Coeff[7042] <= 15'b101000000000000;
		Coeff[7043] <= 15'b101000000000011;
		Coeff[7044] <= 15'b101000000000101;
		Coeff[7045] <= 15'b101000000001000;
		Coeff[7046] <= 15'b101000000001010;
		Coeff[7047] <= 15'b101000000001101;
		Coeff[7048] <= 15'b101000000001111;
		Coeff[7049] <= 15'b101000000010001;
		Coeff[7050] <= 15'b101000000010100;
		Coeff[7051] <= 15'b101000000010110;
		Coeff[7052] <= 15'b101000000011001;
		Coeff[7053] <= 15'b101000000011011;
		Coeff[7054] <= 15'b101000000011110;
		Coeff[7055] <= 15'b101000000100000;
		Coeff[7056] <= 15'b101000000100011;
		Coeff[7057] <= 15'b101000000100101;
		Coeff[7058] <= 15'b101000000101000;
		Coeff[7059] <= 15'b101000000101010;
		Coeff[7060] <= 15'b101000000101100;
		Coeff[7061] <= 15'b101000000101111;
		Coeff[7062] <= 15'b101000000110001;
		Coeff[7063] <= 15'b101000000110100;
		Coeff[7064] <= 15'b101000000110110;
		Coeff[7065] <= 15'b101000000111001;
		Coeff[7066] <= 15'b101000000111011;
		Coeff[7067] <= 15'b101000000111110;
		Coeff[7068] <= 15'b101000001000000;
		Coeff[7069] <= 15'b101000001000010;
		Coeff[7070] <= 15'b101000001000101;
		Coeff[7071] <= 15'b101000001000111;
		Coeff[7072] <= 15'b101000001001010;
		Coeff[7073] <= 15'b101000001001100;
		Coeff[7074] <= 15'b101000001001111;
		Coeff[7075] <= 15'b101000001010001;
		Coeff[7076] <= 15'b101000001010100;
		Coeff[7077] <= 15'b101000001010110;
		Coeff[7078] <= 15'b101000001011000;
		Coeff[7079] <= 15'b101000001011011;
		Coeff[7080] <= 15'b101000001011101;
		Coeff[7081] <= 15'b101000001100000;
		Coeff[7082] <= 15'b101000001100010;
		Coeff[7083] <= 15'b101000001100101;
		Coeff[7084] <= 15'b101000001100111;
		Coeff[7085] <= 15'b101000001101010;
		Coeff[7086] <= 15'b101000001101100;
		Coeff[7087] <= 15'b101000001101110;
		Coeff[7088] <= 15'b101000001110001;
		Coeff[7089] <= 15'b101000001110011;
		Coeff[7090] <= 15'b101000001110110;
		Coeff[7091] <= 15'b101000001111000;
		Coeff[7092] <= 15'b101000001111011;
		Coeff[7093] <= 15'b101000001111101;
		Coeff[7094] <= 15'b101000010000000;
		Coeff[7095] <= 15'b101000010000010;
		Coeff[7096] <= 15'b101000010000100;
		Coeff[7097] <= 15'b101000010000111;
		Coeff[7098] <= 15'b101000010001001;
		Coeff[7099] <= 15'b101000010001100;
		Coeff[7100] <= 15'b101000010001110;
		Coeff[7101] <= 15'b101000010010001;
		Coeff[7102] <= 15'b101000010010011;
		Coeff[7103] <= 15'b101000010010110;
		Coeff[7104] <= 15'b101000010011000;
		Coeff[7105] <= 15'b101000010011010;
		Coeff[7106] <= 15'b101000010011101;
		Coeff[7107] <= 15'b101000010011111;
		Coeff[7108] <= 15'b101000010100010;
		Coeff[7109] <= 15'b101000010100100;
		Coeff[7110] <= 15'b101000010100111;
		Coeff[7111] <= 15'b101000010101001;
		Coeff[7112] <= 15'b101000010101100;
		Coeff[7113] <= 15'b101000010101110;
		Coeff[7114] <= 15'b101000010110000;
		Coeff[7115] <= 15'b101000010110011;
		Coeff[7116] <= 15'b101000010110101;
		Coeff[7117] <= 15'b101000010111000;
		Coeff[7118] <= 15'b101000010111010;
		Coeff[7119] <= 15'b101000010111101;
		Coeff[7120] <= 15'b101000010111111;
		Coeff[7121] <= 15'b101000011000001;
		Coeff[7122] <= 15'b101000011000100;
		Coeff[7123] <= 15'b101000011000110;
		Coeff[7124] <= 15'b101000011001001;
		Coeff[7125] <= 15'b101000011001011;
		Coeff[7126] <= 15'b101000011001110;
		Coeff[7127] <= 15'b101000011010000;
		Coeff[7128] <= 15'b101000011010011;
		Coeff[7129] <= 15'b101000011010101;
		Coeff[7130] <= 15'b101000011010111;
		Coeff[7131] <= 15'b101000011011010;
		Coeff[7132] <= 15'b101000011011100;
		Coeff[7133] <= 15'b101000011011111;
		Coeff[7134] <= 15'b101000011100001;
		Coeff[7135] <= 15'b101000011100100;
		Coeff[7136] <= 15'b101000011100110;
		Coeff[7137] <= 15'b101000011101000;
		Coeff[7138] <= 15'b101000011101011;
		Coeff[7139] <= 15'b101000011101101;
		Coeff[7140] <= 15'b101000011110000;
		Coeff[7141] <= 15'b101000011110010;
		Coeff[7142] <= 15'b101000011110101;
		Coeff[7143] <= 15'b101000011110111;
		Coeff[7144] <= 15'b101000011111001;
		Coeff[7145] <= 15'b101000011111100;
		Coeff[7146] <= 15'b101000011111110;
		Coeff[7147] <= 15'b101000100000001;
		Coeff[7148] <= 15'b101000100000011;
		Coeff[7149] <= 15'b101000100000110;
		Coeff[7150] <= 15'b101000100001000;
		Coeff[7151] <= 15'b101000100001010;
		Coeff[7152] <= 15'b101000100001101;
		Coeff[7153] <= 15'b101000100001111;
		Coeff[7154] <= 15'b101000100010010;
		Coeff[7155] <= 15'b101000100010100;
		Coeff[7156] <= 15'b101000100010111;
		Coeff[7157] <= 15'b101000100011001;
		Coeff[7158] <= 15'b101000100011100;
		Coeff[7159] <= 15'b101000100011110;
		Coeff[7160] <= 15'b101000100100000;
		Coeff[7161] <= 15'b101000100100011;
		Coeff[7162] <= 15'b101000100100101;
		Coeff[7163] <= 15'b101000100101000;
		Coeff[7164] <= 15'b101000100101010;
		Coeff[7165] <= 15'b101000100101101;
		Coeff[7166] <= 15'b101000100101111;
		Coeff[7167] <= 15'b101000100110001;
		Coeff[7168] <= 15'b101000100110100;
		Coeff[7169] <= 15'b101000100110110;
		Coeff[7170] <= 15'b101000100111001;
		Coeff[7171] <= 15'b101000100111011;
		Coeff[7172] <= 15'b101000100111110;
		Coeff[7173] <= 15'b101000101000000;
		Coeff[7174] <= 15'b101000101000010;
		Coeff[7175] <= 15'b101000101000101;
		Coeff[7176] <= 15'b101000101000111;
		Coeff[7177] <= 15'b101000101001010;
		Coeff[7178] <= 15'b101000101001100;
		Coeff[7179] <= 15'b101000101001111;
		Coeff[7180] <= 15'b101000101010001;
		Coeff[7181] <= 15'b101000101010011;
		Coeff[7182] <= 15'b101000101010110;
		Coeff[7183] <= 15'b101000101011000;
		Coeff[7184] <= 15'b101000101011011;
		Coeff[7185] <= 15'b101000101011101;
		Coeff[7186] <= 15'b101000101011111;
		Coeff[7187] <= 15'b101000101100010;
		Coeff[7188] <= 15'b101000101100100;
		Coeff[7189] <= 15'b101000101100111;
		Coeff[7190] <= 15'b101000101101001;
		Coeff[7191] <= 15'b101000101101100;
		Coeff[7192] <= 15'b101000101101110;
		Coeff[7193] <= 15'b101000101110000;
		Coeff[7194] <= 15'b101000101110011;
		Coeff[7195] <= 15'b101000101110101;
		Coeff[7196] <= 15'b101000101111000;
		Coeff[7197] <= 15'b101000101111010;
		Coeff[7198] <= 15'b101000101111101;
		Coeff[7199] <= 15'b101000101111111;
		Coeff[7200] <= 15'b101000110000001;
		Coeff[7201] <= 15'b101000110000100;
		Coeff[7202] <= 15'b101000110000110;
		Coeff[7203] <= 15'b101000110001001;
		Coeff[7204] <= 15'b101000110001011;
		Coeff[7205] <= 15'b101000110001110;
		Coeff[7206] <= 15'b101000110010000;
		Coeff[7207] <= 15'b101000110010010;
		Coeff[7208] <= 15'b101000110010101;
		Coeff[7209] <= 15'b101000110010111;
		Coeff[7210] <= 15'b101000110011010;
		Coeff[7211] <= 15'b101000110011100;
		Coeff[7212] <= 15'b101000110011110;
		Coeff[7213] <= 15'b101000110100001;
		Coeff[7214] <= 15'b101000110100011;
		Coeff[7215] <= 15'b101000110100110;
		Coeff[7216] <= 15'b101000110101000;
		Coeff[7217] <= 15'b101000110101011;
		Coeff[7218] <= 15'b101000110101101;
		Coeff[7219] <= 15'b101000110101111;
		Coeff[7220] <= 15'b101000110110010;
		Coeff[7221] <= 15'b101000110110100;
		Coeff[7222] <= 15'b101000110110111;
		Coeff[7223] <= 15'b101000110111001;
		Coeff[7224] <= 15'b101000110111011;
		Coeff[7225] <= 15'b101000110111110;
		Coeff[7226] <= 15'b101000111000000;
		Coeff[7227] <= 15'b101000111000011;
		Coeff[7228] <= 15'b101000111000101;
		Coeff[7229] <= 15'b101000111001000;
		Coeff[7230] <= 15'b101000111001010;
		Coeff[7231] <= 15'b101000111001100;
		Coeff[7232] <= 15'b101000111001111;
		Coeff[7233] <= 15'b101000111010001;
		Coeff[7234] <= 15'b101000111010100;
		Coeff[7235] <= 15'b101000111010110;
		Coeff[7236] <= 15'b101000111011000;
		Coeff[7237] <= 15'b101000111011011;
		Coeff[7238] <= 15'b101000111011101;
		Coeff[7239] <= 15'b101000111100000;
		Coeff[7240] <= 15'b101000111100010;
		Coeff[7241] <= 15'b101000111100101;
		Coeff[7242] <= 15'b101000111100111;
		Coeff[7243] <= 15'b101000111101001;
		Coeff[7244] <= 15'b101000111101100;
		Coeff[7245] <= 15'b101000111101110;
		Coeff[7246] <= 15'b101000111110001;
		Coeff[7247] <= 15'b101000111110011;
		Coeff[7248] <= 15'b101000111110101;
		Coeff[7249] <= 15'b101000111111000;
		Coeff[7250] <= 15'b101000111111010;
		Coeff[7251] <= 15'b101000111111101;
		Coeff[7252] <= 15'b101000111111111;
		Coeff[7253] <= 15'b101001000000010;
		Coeff[7254] <= 15'b101001000000100;
		Coeff[7255] <= 15'b101001000000110;
		Coeff[7256] <= 15'b101001000001001;
		Coeff[7257] <= 15'b101001000001011;
		Coeff[7258] <= 15'b101001000001110;
		Coeff[7259] <= 15'b101001000010000;
		Coeff[7260] <= 15'b101001000010010;
		Coeff[7261] <= 15'b101001000010101;
		Coeff[7262] <= 15'b101001000010111;
		Coeff[7263] <= 15'b101001000011010;
		Coeff[7264] <= 15'b101001000011100;
		Coeff[7265] <= 15'b101001000011110;
		Coeff[7266] <= 15'b101001000100001;
		Coeff[7267] <= 15'b101001000100011;
		Coeff[7268] <= 15'b101001000100110;
		Coeff[7269] <= 15'b101001000101000;
		Coeff[7270] <= 15'b101001000101011;
		Coeff[7271] <= 15'b101001000101101;
		Coeff[7272] <= 15'b101001000101111;
		Coeff[7273] <= 15'b101001000110010;
		Coeff[7274] <= 15'b101001000110100;
		Coeff[7275] <= 15'b101001000110111;
		Coeff[7276] <= 15'b101001000111001;
		Coeff[7277] <= 15'b101001000111011;
		Coeff[7278] <= 15'b101001000111110;
		Coeff[7279] <= 15'b101001001000000;
		Coeff[7280] <= 15'b101001001000011;
		Coeff[7281] <= 15'b101001001000101;
		Coeff[7282] <= 15'b101001001000111;
		Coeff[7283] <= 15'b101001001001010;
		Coeff[7284] <= 15'b101001001001100;
		Coeff[7285] <= 15'b101001001001111;
		Coeff[7286] <= 15'b101001001010001;
		Coeff[7287] <= 15'b101001001010011;
		Coeff[7288] <= 15'b101001001010110;
		Coeff[7289] <= 15'b101001001011000;
		Coeff[7290] <= 15'b101001001011011;
		Coeff[7291] <= 15'b101001001011101;
		Coeff[7292] <= 15'b101001001011111;
		Coeff[7293] <= 15'b101001001100010;
		Coeff[7294] <= 15'b101001001100100;
		Coeff[7295] <= 15'b101001001100111;
		Coeff[7296] <= 15'b101001001101001;
		Coeff[7297] <= 15'b101001001101011;
		Coeff[7298] <= 15'b101001001101110;
		Coeff[7299] <= 15'b101001001110000;
		Coeff[7300] <= 15'b101001001110011;
		Coeff[7301] <= 15'b101001001110101;
		Coeff[7302] <= 15'b101001001110111;
		Coeff[7303] <= 15'b101001001111010;
		Coeff[7304] <= 15'b101001001111100;
		Coeff[7305] <= 15'b101001001111111;
		Coeff[7306] <= 15'b101001010000001;
		Coeff[7307] <= 15'b101001010000100;
		Coeff[7308] <= 15'b101001010000110;
		Coeff[7309] <= 15'b101001010001000;
		Coeff[7310] <= 15'b101001010001011;
		Coeff[7311] <= 15'b101001010001101;
		Coeff[7312] <= 15'b101001010010000;
		Coeff[7313] <= 15'b101001010010010;
		Coeff[7314] <= 15'b101001010010100;
		Coeff[7315] <= 15'b101001010010111;
		Coeff[7316] <= 15'b101001010011001;
		Coeff[7317] <= 15'b101001010011100;
		Coeff[7318] <= 15'b101001010011110;
		Coeff[7319] <= 15'b101001010100000;
		Coeff[7320] <= 15'b101001010100011;
		Coeff[7321] <= 15'b101001010100101;
		Coeff[7322] <= 15'b101001010101000;
		Coeff[7323] <= 15'b101001010101010;
		Coeff[7324] <= 15'b101001010101100;
		Coeff[7325] <= 15'b101001010101111;
		Coeff[7326] <= 15'b101001010110001;
		Coeff[7327] <= 15'b101001010110011;
		Coeff[7328] <= 15'b101001010110110;
		Coeff[7329] <= 15'b101001010111000;
		Coeff[7330] <= 15'b101001010111011;
		Coeff[7331] <= 15'b101001010111101;
		Coeff[7332] <= 15'b101001010111111;
		Coeff[7333] <= 15'b101001011000010;
		Coeff[7334] <= 15'b101001011000100;
		Coeff[7335] <= 15'b101001011000111;
		Coeff[7336] <= 15'b101001011001001;
		Coeff[7337] <= 15'b101001011001011;
		Coeff[7338] <= 15'b101001011001110;
		Coeff[7339] <= 15'b101001011010000;
		Coeff[7340] <= 15'b101001011010011;
		Coeff[7341] <= 15'b101001011010101;
		Coeff[7342] <= 15'b101001011010111;
		Coeff[7343] <= 15'b101001011011010;
		Coeff[7344] <= 15'b101001011011100;
		Coeff[7345] <= 15'b101001011011111;
		Coeff[7346] <= 15'b101001011100001;
		Coeff[7347] <= 15'b101001011100011;
		Coeff[7348] <= 15'b101001011100110;
		Coeff[7349] <= 15'b101001011101000;
		Coeff[7350] <= 15'b101001011101011;
		Coeff[7351] <= 15'b101001011101101;
		Coeff[7352] <= 15'b101001011101111;
		Coeff[7353] <= 15'b101001011110010;
		Coeff[7354] <= 15'b101001011110100;
		Coeff[7355] <= 15'b101001011110111;
		Coeff[7356] <= 15'b101001011111001;
		Coeff[7357] <= 15'b101001011111011;
		Coeff[7358] <= 15'b101001011111110;
		Coeff[7359] <= 15'b101001100000000;
		Coeff[7360] <= 15'b101001100000011;
		Coeff[7361] <= 15'b101001100000101;
		Coeff[7362] <= 15'b101001100000111;
		Coeff[7363] <= 15'b101001100001010;
		Coeff[7364] <= 15'b101001100001100;
		Coeff[7365] <= 15'b101001100001110;
		Coeff[7366] <= 15'b101001100010001;
		Coeff[7367] <= 15'b101001100010011;
		Coeff[7368] <= 15'b101001100010110;
		Coeff[7369] <= 15'b101001100011000;
		Coeff[7370] <= 15'b101001100011010;
		Coeff[7371] <= 15'b101001100011101;
		Coeff[7372] <= 15'b101001100011111;
		Coeff[7373] <= 15'b101001100100010;
		Coeff[7374] <= 15'b101001100100100;
		Coeff[7375] <= 15'b101001100100110;
		Coeff[7376] <= 15'b101001100101001;
		Coeff[7377] <= 15'b101001100101011;
		Coeff[7378] <= 15'b101001100101110;
		Coeff[7379] <= 15'b101001100110000;
		Coeff[7380] <= 15'b101001100110010;
		Coeff[7381] <= 15'b101001100110101;
		Coeff[7382] <= 15'b101001100110111;
		Coeff[7383] <= 15'b101001100111001;
		Coeff[7384] <= 15'b101001100111100;
		Coeff[7385] <= 15'b101001100111110;
		Coeff[7386] <= 15'b101001101000001;
		Coeff[7387] <= 15'b101001101000011;
		Coeff[7388] <= 15'b101001101000101;
		Coeff[7389] <= 15'b101001101001000;
		Coeff[7390] <= 15'b101001101001010;
		Coeff[7391] <= 15'b101001101001101;
		Coeff[7392] <= 15'b101001101001111;
		Coeff[7393] <= 15'b101001101010001;
		Coeff[7394] <= 15'b101001101010100;
		Coeff[7395] <= 15'b101001101010110;
		Coeff[7396] <= 15'b101001101011000;
		Coeff[7397] <= 15'b101001101011011;
		Coeff[7398] <= 15'b101001101011101;
		Coeff[7399] <= 15'b101001101100000;
		Coeff[7400] <= 15'b101001101100010;
		Coeff[7401] <= 15'b101001101100100;
		Coeff[7402] <= 15'b101001101100111;
		Coeff[7403] <= 15'b101001101101001;
		Coeff[7404] <= 15'b101001101101100;
		Coeff[7405] <= 15'b101001101101110;
		Coeff[7406] <= 15'b101001101110000;
		Coeff[7407] <= 15'b101001101110011;
		Coeff[7408] <= 15'b101001101110101;
		Coeff[7409] <= 15'b101001101110111;
		Coeff[7410] <= 15'b101001101111010;
		Coeff[7411] <= 15'b101001101111100;
		Coeff[7412] <= 15'b101001101111111;
		Coeff[7413] <= 15'b101001110000001;
		Coeff[7414] <= 15'b101001110000011;
		Coeff[7415] <= 15'b101001110000110;
		Coeff[7416] <= 15'b101001110001000;
		Coeff[7417] <= 15'b101001110001011;
		Coeff[7418] <= 15'b101001110001101;
		Coeff[7419] <= 15'b101001110001111;
		Coeff[7420] <= 15'b101001110010010;
		Coeff[7421] <= 15'b101001110010100;
		Coeff[7422] <= 15'b101001110010110;
		Coeff[7423] <= 15'b101001110011001;
		Coeff[7424] <= 15'b101001110011011;
		Coeff[7425] <= 15'b101001110011110;
		Coeff[7426] <= 15'b101001110100000;
		Coeff[7427] <= 15'b101001110100010;
		Coeff[7428] <= 15'b101001110100101;
		Coeff[7429] <= 15'b101001110100111;
		Coeff[7430] <= 15'b101001110101001;
		Coeff[7431] <= 15'b101001110101100;
		Coeff[7432] <= 15'b101001110101110;
		Coeff[7433] <= 15'b101001110110001;
		Coeff[7434] <= 15'b101001110110011;
		Coeff[7435] <= 15'b101001110110101;
		Coeff[7436] <= 15'b101001110111000;
		Coeff[7437] <= 15'b101001110111010;
		Coeff[7438] <= 15'b101001110111100;
		Coeff[7439] <= 15'b101001110111111;
		Coeff[7440] <= 15'b101001111000001;
		Coeff[7441] <= 15'b101001111000100;
		Coeff[7442] <= 15'b101001111000110;
		Coeff[7443] <= 15'b101001111001000;
		Coeff[7444] <= 15'b101001111001011;
		Coeff[7445] <= 15'b101001111001101;
		Coeff[7446] <= 15'b101001111001111;
		Coeff[7447] <= 15'b101001111010010;
		Coeff[7448] <= 15'b101001111010100;
		Coeff[7449] <= 15'b101001111010111;
		Coeff[7450] <= 15'b101001111011001;
		Coeff[7451] <= 15'b101001111011011;
		Coeff[7452] <= 15'b101001111011110;
		Coeff[7453] <= 15'b101001111100000;
		Coeff[7454] <= 15'b101001111100010;
		Coeff[7455] <= 15'b101001111100101;
		Coeff[7456] <= 15'b101001111100111;
		Coeff[7457] <= 15'b101001111101010;
		Coeff[7458] <= 15'b101001111101100;
		Coeff[7459] <= 15'b101001111101110;
		Coeff[7460] <= 15'b101001111110001;
		Coeff[7461] <= 15'b101001111110011;
		Coeff[7462] <= 15'b101001111110101;
		Coeff[7463] <= 15'b101001111111000;
		Coeff[7464] <= 15'b101001111111010;
		Coeff[7465] <= 15'b101001111111101;
		Coeff[7466] <= 15'b101001111111111;
		Coeff[7467] <= 15'b101010000000001;
		Coeff[7468] <= 15'b101010000000100;
		Coeff[7469] <= 15'b101010000000110;
		Coeff[7470] <= 15'b101010000001000;
		Coeff[7471] <= 15'b101010000001011;
		Coeff[7472] <= 15'b101010000001101;
		Coeff[7473] <= 15'b101010000001111;
		Coeff[7474] <= 15'b101010000010010;
		Coeff[7475] <= 15'b101010000010100;
		Coeff[7476] <= 15'b101010000010111;
		Coeff[7477] <= 15'b101010000011001;
		Coeff[7478] <= 15'b101010000011011;
		Coeff[7479] <= 15'b101010000011110;
		Coeff[7480] <= 15'b101010000100000;
		Coeff[7481] <= 15'b101010000100010;
		Coeff[7482] <= 15'b101010000100101;
		Coeff[7483] <= 15'b101010000100111;
		Coeff[7484] <= 15'b101010000101010;
		Coeff[7485] <= 15'b101010000101100;
		Coeff[7486] <= 15'b101010000101110;
		Coeff[7487] <= 15'b101010000110001;
		Coeff[7488] <= 15'b101010000110011;
		Coeff[7489] <= 15'b101010000110101;
		Coeff[7490] <= 15'b101010000111000;
		Coeff[7491] <= 15'b101010000111010;
		Coeff[7492] <= 15'b101010000111100;
		Coeff[7493] <= 15'b101010000111111;
		Coeff[7494] <= 15'b101010001000001;
		Coeff[7495] <= 15'b101010001000100;
		Coeff[7496] <= 15'b101010001000110;
		Coeff[7497] <= 15'b101010001001000;
		Coeff[7498] <= 15'b101010001001011;
		Coeff[7499] <= 15'b101010001001101;
		Coeff[7500] <= 15'b101010001001111;
		Coeff[7501] <= 15'b101010001010010;
		Coeff[7502] <= 15'b101010001010100;
		Coeff[7503] <= 15'b101010001010110;
		Coeff[7504] <= 15'b101010001011001;
		Coeff[7505] <= 15'b101010001011011;
		Coeff[7506] <= 15'b101010001011110;
		Coeff[7507] <= 15'b101010001100000;
		Coeff[7508] <= 15'b101010001100010;
		Coeff[7509] <= 15'b101010001100101;
		Coeff[7510] <= 15'b101010001100111;
		Coeff[7511] <= 15'b101010001101001;
		Coeff[7512] <= 15'b101010001101100;
		Coeff[7513] <= 15'b101010001101110;
		Coeff[7514] <= 15'b101010001110000;
		Coeff[7515] <= 15'b101010001110011;
		Coeff[7516] <= 15'b101010001110101;
		Coeff[7517] <= 15'b101010001111000;
		Coeff[7518] <= 15'b101010001111010;
		Coeff[7519] <= 15'b101010001111100;
		Coeff[7520] <= 15'b101010001111111;
		Coeff[7521] <= 15'b101010010000001;
		Coeff[7522] <= 15'b101010010000011;
		Coeff[7523] <= 15'b101010010000110;
		Coeff[7524] <= 15'b101010010001000;
		Coeff[7525] <= 15'b101010010001010;
		Coeff[7526] <= 15'b101010010001101;
		Coeff[7527] <= 15'b101010010001111;
		Coeff[7528] <= 15'b101010010010001;
		Coeff[7529] <= 15'b101010010010100;
		Coeff[7530] <= 15'b101010010010110;
		Coeff[7531] <= 15'b101010010011001;
		Coeff[7532] <= 15'b101010010011011;
		Coeff[7533] <= 15'b101010010011101;
		Coeff[7534] <= 15'b101010010100000;
		Coeff[7535] <= 15'b101010010100010;
		Coeff[7536] <= 15'b101010010100100;
		Coeff[7537] <= 15'b101010010100111;
		Coeff[7538] <= 15'b101010010101001;
		Coeff[7539] <= 15'b101010010101011;
		Coeff[7540] <= 15'b101010010101110;
		Coeff[7541] <= 15'b101010010110000;
		Coeff[7542] <= 15'b101010010110010;
		Coeff[7543] <= 15'b101010010110101;
		Coeff[7544] <= 15'b101010010110111;
		Coeff[7545] <= 15'b101010010111010;
		Coeff[7546] <= 15'b101010010111100;
		Coeff[7547] <= 15'b101010010111110;
		Coeff[7548] <= 15'b101010011000001;
		Coeff[7549] <= 15'b101010011000011;
		Coeff[7550] <= 15'b101010011000101;
		Coeff[7551] <= 15'b101010011001000;
		Coeff[7552] <= 15'b101010011001010;
		Coeff[7553] <= 15'b101010011001100;
		Coeff[7554] <= 15'b101010011001111;
		Coeff[7555] <= 15'b101010011010001;
		Coeff[7556] <= 15'b101010011010011;
		Coeff[7557] <= 15'b101010011010110;
		Coeff[7558] <= 15'b101010011011000;
		Coeff[7559] <= 15'b101010011011011;
		Coeff[7560] <= 15'b101010011011101;
		Coeff[7561] <= 15'b101010011011111;
		Coeff[7562] <= 15'b101010011100010;
		Coeff[7563] <= 15'b101010011100100;
		Coeff[7564] <= 15'b101010011100110;
		Coeff[7565] <= 15'b101010011101001;
		Coeff[7566] <= 15'b101010011101011;
		Coeff[7567] <= 15'b101010011101101;
		Coeff[7568] <= 15'b101010011110000;
		Coeff[7569] <= 15'b101010011110010;
		Coeff[7570] <= 15'b101010011110100;
		Coeff[7571] <= 15'b101010011110111;
		Coeff[7572] <= 15'b101010011111001;
		Coeff[7573] <= 15'b101010011111011;
		Coeff[7574] <= 15'b101010011111110;
		Coeff[7575] <= 15'b101010100000000;
		Coeff[7576] <= 15'b101010100000010;
		Coeff[7577] <= 15'b101010100000101;
		Coeff[7578] <= 15'b101010100000111;
		Coeff[7579] <= 15'b101010100001010;
		Coeff[7580] <= 15'b101010100001100;
		Coeff[7581] <= 15'b101010100001110;
		Coeff[7582] <= 15'b101010100010001;
		Coeff[7583] <= 15'b101010100010011;
		Coeff[7584] <= 15'b101010100010101;
		Coeff[7585] <= 15'b101010100011000;
		Coeff[7586] <= 15'b101010100011010;
		Coeff[7587] <= 15'b101010100011100;
		Coeff[7588] <= 15'b101010100011111;
		Coeff[7589] <= 15'b101010100100001;
		Coeff[7590] <= 15'b101010100100011;
		Coeff[7591] <= 15'b101010100100110;
		Coeff[7592] <= 15'b101010100101000;
		Coeff[7593] <= 15'b101010100101010;
		Coeff[7594] <= 15'b101010100101101;
		Coeff[7595] <= 15'b101010100101111;
		Coeff[7596] <= 15'b101010100110001;
		Coeff[7597] <= 15'b101010100110100;
		Coeff[7598] <= 15'b101010100110110;
		Coeff[7599] <= 15'b101010100111000;
		Coeff[7600] <= 15'b101010100111011;
		Coeff[7601] <= 15'b101010100111101;
		Coeff[7602] <= 15'b101010100111111;
		Coeff[7603] <= 15'b101010101000010;
		Coeff[7604] <= 15'b101010101000100;
		Coeff[7605] <= 15'b101010101000110;
		Coeff[7606] <= 15'b101010101001001;
		Coeff[7607] <= 15'b101010101001011;
		Coeff[7608] <= 15'b101010101001110;
		Coeff[7609] <= 15'b101010101010000;
		Coeff[7610] <= 15'b101010101010010;
		Coeff[7611] <= 15'b101010101010101;
		Coeff[7612] <= 15'b101010101010111;
		Coeff[7613] <= 15'b101010101011001;
		Coeff[7614] <= 15'b101010101011100;
		Coeff[7615] <= 15'b101010101011110;
		Coeff[7616] <= 15'b101010101100000;
		Coeff[7617] <= 15'b101010101100011;
		Coeff[7618] <= 15'b101010101100101;
		Coeff[7619] <= 15'b101010101100111;
		Coeff[7620] <= 15'b101010101101010;
		Coeff[7621] <= 15'b101010101101100;
		Coeff[7622] <= 15'b101010101101110;
		Coeff[7623] <= 15'b101010101110001;
		Coeff[7624] <= 15'b101010101110011;
		Coeff[7625] <= 15'b101010101110101;
		Coeff[7626] <= 15'b101010101111000;
		Coeff[7627] <= 15'b101010101111010;
		Coeff[7628] <= 15'b101010101111100;
		Coeff[7629] <= 15'b101010101111111;
		Coeff[7630] <= 15'b101010110000001;
		Coeff[7631] <= 15'b101010110000011;
		Coeff[7632] <= 15'b101010110000110;
		Coeff[7633] <= 15'b101010110001000;
		Coeff[7634] <= 15'b101010110001010;
		Coeff[7635] <= 15'b101010110001101;
		Coeff[7636] <= 15'b101010110001111;
		Coeff[7637] <= 15'b101010110010001;
		Coeff[7638] <= 15'b101010110010100;
		Coeff[7639] <= 15'b101010110010110;
		Coeff[7640] <= 15'b101010110011000;
		Coeff[7641] <= 15'b101010110011011;
		Coeff[7642] <= 15'b101010110011101;
		Coeff[7643] <= 15'b101010110011111;
		Coeff[7644] <= 15'b101010110100010;
		Coeff[7645] <= 15'b101010110100100;
		Coeff[7646] <= 15'b101010110100110;
		Coeff[7647] <= 15'b101010110101001;
		Coeff[7648] <= 15'b101010110101011;
		Coeff[7649] <= 15'b101010110101101;
		Coeff[7650] <= 15'b101010110110000;
		Coeff[7651] <= 15'b101010110110010;
		Coeff[7652] <= 15'b101010110110100;
		Coeff[7653] <= 15'b101010110110111;
		Coeff[7654] <= 15'b101010110111001;
		Coeff[7655] <= 15'b101010110111011;
		Coeff[7656] <= 15'b101010110111110;
		Coeff[7657] <= 15'b101010111000000;
		Coeff[7658] <= 15'b101010111000010;
		Coeff[7659] <= 15'b101010111000101;
		Coeff[7660] <= 15'b101010111000111;
		Coeff[7661] <= 15'b101010111001001;
		Coeff[7662] <= 15'b101010111001100;
		Coeff[7663] <= 15'b101010111001110;
		Coeff[7664] <= 15'b101010111010000;
		Coeff[7665] <= 15'b101010111010011;
		Coeff[7666] <= 15'b101010111010101;
		Coeff[7667] <= 15'b101010111010111;
		Coeff[7668] <= 15'b101010111011010;
		Coeff[7669] <= 15'b101010111011100;
		Coeff[7670] <= 15'b101010111011110;
		Coeff[7671] <= 15'b101010111100001;
		Coeff[7672] <= 15'b101010111100011;
		Coeff[7673] <= 15'b101010111100101;
		Coeff[7674] <= 15'b101010111101000;
		Coeff[7675] <= 15'b101010111101010;
		Coeff[7676] <= 15'b101010111101100;
		Coeff[7677] <= 15'b101010111101111;
		Coeff[7678] <= 15'b101010111110001;
		Coeff[7679] <= 15'b101010111110011;
		Coeff[7680] <= 15'b101010111110110;
		Coeff[7681] <= 15'b101010111111000;
		Coeff[7682] <= 15'b101010111111010;
		Coeff[7683] <= 15'b101010111111101;
		Coeff[7684] <= 15'b101010111111111;
		Coeff[7685] <= 15'b101011000000001;
		Coeff[7686] <= 15'b101011000000100;
		Coeff[7687] <= 15'b101011000000110;
		Coeff[7688] <= 15'b101011000001000;
		Coeff[7689] <= 15'b101011000001011;
		Coeff[7690] <= 15'b101011000001101;
		Coeff[7691] <= 15'b101011000001111;
		Coeff[7692] <= 15'b101011000010010;
		Coeff[7693] <= 15'b101011000010100;
		Coeff[7694] <= 15'b101011000010110;
		Coeff[7695] <= 15'b101011000011001;
		Coeff[7696] <= 15'b101011000011011;
		Coeff[7697] <= 15'b101011000011101;
		Coeff[7698] <= 15'b101011000100000;
		Coeff[7699] <= 15'b101011000100010;
		Coeff[7700] <= 15'b101011000100100;
		Coeff[7701] <= 15'b101011000100110;
		Coeff[7702] <= 15'b101011000101001;
		Coeff[7703] <= 15'b101011000101011;
		Coeff[7704] <= 15'b101011000101101;
		Coeff[7705] <= 15'b101011000110000;
		Coeff[7706] <= 15'b101011000110010;
		Coeff[7707] <= 15'b101011000110100;
		Coeff[7708] <= 15'b101011000110111;
		Coeff[7709] <= 15'b101011000111001;
		Coeff[7710] <= 15'b101011000111011;
		Coeff[7711] <= 15'b101011000111110;
		Coeff[7712] <= 15'b101011001000000;
		Coeff[7713] <= 15'b101011001000010;
		Coeff[7714] <= 15'b101011001000101;
		Coeff[7715] <= 15'b101011001000111;
		Coeff[7716] <= 15'b101011001001001;
		Coeff[7717] <= 15'b101011001001100;
		Coeff[7718] <= 15'b101011001001110;
		Coeff[7719] <= 15'b101011001010000;
		Coeff[7720] <= 15'b101011001010011;
		Coeff[7721] <= 15'b101011001010101;
		Coeff[7722] <= 15'b101011001010111;
		Coeff[7723] <= 15'b101011001011010;
		Coeff[7724] <= 15'b101011001011100;
		Coeff[7725] <= 15'b101011001011110;
		Coeff[7726] <= 15'b101011001100001;
		Coeff[7727] <= 15'b101011001100011;
		Coeff[7728] <= 15'b101011001100101;
		Coeff[7729] <= 15'b101011001100111;
		Coeff[7730] <= 15'b101011001101010;
		Coeff[7731] <= 15'b101011001101100;
		Coeff[7732] <= 15'b101011001101110;
		Coeff[7733] <= 15'b101011001110001;
		Coeff[7734] <= 15'b101011001110011;
		Coeff[7735] <= 15'b101011001110101;
		Coeff[7736] <= 15'b101011001111000;
		Coeff[7737] <= 15'b101011001111010;
		Coeff[7738] <= 15'b101011001111100;
		Coeff[7739] <= 15'b101011001111111;
		Coeff[7740] <= 15'b101011010000001;
		Coeff[7741] <= 15'b101011010000011;
		Coeff[7742] <= 15'b101011010000110;
		Coeff[7743] <= 15'b101011010001000;
		Coeff[7744] <= 15'b101011010001010;
		Coeff[7745] <= 15'b101011010001101;
		Coeff[7746] <= 15'b101011010001111;
		Coeff[7747] <= 15'b101011010010001;
		Coeff[7748] <= 15'b101011010010011;
		Coeff[7749] <= 15'b101011010010110;
		Coeff[7750] <= 15'b101011010011000;
		Coeff[7751] <= 15'b101011010011010;
		Coeff[7752] <= 15'b101011010011101;
		Coeff[7753] <= 15'b101011010011111;
		Coeff[7754] <= 15'b101011010100001;
		Coeff[7755] <= 15'b101011010100100;
		Coeff[7756] <= 15'b101011010100110;
		Coeff[7757] <= 15'b101011010101000;
		Coeff[7758] <= 15'b101011010101011;
		Coeff[7759] <= 15'b101011010101101;
		Coeff[7760] <= 15'b101011010101111;
		Coeff[7761] <= 15'b101011010110010;
		Coeff[7762] <= 15'b101011010110100;
		Coeff[7763] <= 15'b101011010110110;
		Coeff[7764] <= 15'b101011010111000;
		Coeff[7765] <= 15'b101011010111011;
		Coeff[7766] <= 15'b101011010111101;
		Coeff[7767] <= 15'b101011010111111;
		Coeff[7768] <= 15'b101011011000010;
		Coeff[7769] <= 15'b101011011000100;
		Coeff[7770] <= 15'b101011011000110;
		Coeff[7771] <= 15'b101011011001001;
		Coeff[7772] <= 15'b101011011001011;
		Coeff[7773] <= 15'b101011011001101;
		Coeff[7774] <= 15'b101011011010000;
		Coeff[7775] <= 15'b101011011010010;
		Coeff[7776] <= 15'b101011011010100;
		Coeff[7777] <= 15'b101011011010110;
		Coeff[7778] <= 15'b101011011011001;
		Coeff[7779] <= 15'b101011011011011;
		Coeff[7780] <= 15'b101011011011101;
		Coeff[7781] <= 15'b101011011100000;
		Coeff[7782] <= 15'b101011011100010;
		Coeff[7783] <= 15'b101011011100100;
		Coeff[7784] <= 15'b101011011100111;
		Coeff[7785] <= 15'b101011011101001;
		Coeff[7786] <= 15'b101011011101011;
		Coeff[7787] <= 15'b101011011101110;
		Coeff[7788] <= 15'b101011011110000;
		Coeff[7789] <= 15'b101011011110010;
		Coeff[7790] <= 15'b101011011110100;
		Coeff[7791] <= 15'b101011011110111;
		Coeff[7792] <= 15'b101011011111001;
		Coeff[7793] <= 15'b101011011111011;
		Coeff[7794] <= 15'b101011011111110;
		Coeff[7795] <= 15'b101011100000000;
		Coeff[7796] <= 15'b101011100000010;
		Coeff[7797] <= 15'b101011100000101;
		Coeff[7798] <= 15'b101011100000111;
		Coeff[7799] <= 15'b101011100001001;
		Coeff[7800] <= 15'b101011100001100;
		Coeff[7801] <= 15'b101011100001110;
		Coeff[7802] <= 15'b101011100010000;
		Coeff[7803] <= 15'b101011100010010;
		Coeff[7804] <= 15'b101011100010101;
		Coeff[7805] <= 15'b101011100010111;
		Coeff[7806] <= 15'b101011100011001;
		Coeff[7807] <= 15'b101011100011100;
		Coeff[7808] <= 15'b101011100011110;
		Coeff[7809] <= 15'b101011100100000;
		Coeff[7810] <= 15'b101011100100011;
		Coeff[7811] <= 15'b101011100100101;
		Coeff[7812] <= 15'b101011100100111;
		Coeff[7813] <= 15'b101011100101001;
		Coeff[7814] <= 15'b101011100101100;
		Coeff[7815] <= 15'b101011100101110;
		Coeff[7816] <= 15'b101011100110000;
		Coeff[7817] <= 15'b101011100110011;
		Coeff[7818] <= 15'b101011100110101;
		Coeff[7819] <= 15'b101011100110111;
		Coeff[7820] <= 15'b101011100111010;
		Coeff[7821] <= 15'b101011100111100;
		Coeff[7822] <= 15'b101011100111110;
		Coeff[7823] <= 15'b101011101000000;
		Coeff[7824] <= 15'b101011101000011;
		Coeff[7825] <= 15'b101011101000101;
		Coeff[7826] <= 15'b101011101000111;
		Coeff[7827] <= 15'b101011101001010;
		Coeff[7828] <= 15'b101011101001100;
		Coeff[7829] <= 15'b101011101001110;
		Coeff[7830] <= 15'b101011101010001;
		Coeff[7831] <= 15'b101011101010011;
		Coeff[7832] <= 15'b101011101010101;
		Coeff[7833] <= 15'b101011101010111;
		Coeff[7834] <= 15'b101011101011010;
		Coeff[7835] <= 15'b101011101011100;
		Coeff[7836] <= 15'b101011101011110;
		Coeff[7837] <= 15'b101011101100001;
		Coeff[7838] <= 15'b101011101100011;
		Coeff[7839] <= 15'b101011101100101;
		Coeff[7840] <= 15'b101011101100111;
		Coeff[7841] <= 15'b101011101101010;
		Coeff[7842] <= 15'b101011101101100;
		Coeff[7843] <= 15'b101011101101110;
		Coeff[7844] <= 15'b101011101110001;
		Coeff[7845] <= 15'b101011101110011;
		Coeff[7846] <= 15'b101011101110101;
		Coeff[7847] <= 15'b101011101111000;
		Coeff[7848] <= 15'b101011101111010;
		Coeff[7849] <= 15'b101011101111100;
		Coeff[7850] <= 15'b101011101111110;
		Coeff[7851] <= 15'b101011110000001;
		Coeff[7852] <= 15'b101011110000011;
		Coeff[7853] <= 15'b101011110000101;
		Coeff[7854] <= 15'b101011110001000;
		Coeff[7855] <= 15'b101011110001010;
		Coeff[7856] <= 15'b101011110001100;
		Coeff[7857] <= 15'b101011110001110;
		Coeff[7858] <= 15'b101011110010001;
		Coeff[7859] <= 15'b101011110010011;
		Coeff[7860] <= 15'b101011110010101;
		Coeff[7861] <= 15'b101011110011000;
		Coeff[7862] <= 15'b101011110011010;
		Coeff[7863] <= 15'b101011110011100;
		Coeff[7864] <= 15'b101011110011111;
		Coeff[7865] <= 15'b101011110100001;
		Coeff[7866] <= 15'b101011110100011;
		Coeff[7867] <= 15'b101011110100101;
		Coeff[7868] <= 15'b101011110101000;
		Coeff[7869] <= 15'b101011110101010;
		Coeff[7870] <= 15'b101011110101100;
		Coeff[7871] <= 15'b101011110101111;
		Coeff[7872] <= 15'b101011110110001;
		Coeff[7873] <= 15'b101011110110011;
		Coeff[7874] <= 15'b101011110110101;
		Coeff[7875] <= 15'b101011110111000;
		Coeff[7876] <= 15'b101011110111010;
		Coeff[7877] <= 15'b101011110111100;
		Coeff[7878] <= 15'b101011110111111;
		Coeff[7879] <= 15'b101011111000001;
		Coeff[7880] <= 15'b101011111000011;
		Coeff[7881] <= 15'b101011111000101;
		Coeff[7882] <= 15'b101011111001000;
		Coeff[7883] <= 15'b101011111001010;
		Coeff[7884] <= 15'b101011111001100;
		Coeff[7885] <= 15'b101011111001111;
		Coeff[7886] <= 15'b101011111010001;
		Coeff[7887] <= 15'b101011111010011;
		Coeff[7888] <= 15'b101011111010101;
		Coeff[7889] <= 15'b101011111011000;
		Coeff[7890] <= 15'b101011111011010;
		Coeff[7891] <= 15'b101011111011100;
		Coeff[7892] <= 15'b101011111011111;
		Coeff[7893] <= 15'b101011111100001;
		Coeff[7894] <= 15'b101011111100011;
		Coeff[7895] <= 15'b101011111100101;
		Coeff[7896] <= 15'b101011111101000;
		Coeff[7897] <= 15'b101011111101010;
		Coeff[7898] <= 15'b101011111101100;
		Coeff[7899] <= 15'b101011111101111;
		Coeff[7900] <= 15'b101011111110001;
		Coeff[7901] <= 15'b101011111110011;
		Coeff[7902] <= 15'b101011111110101;
		Coeff[7903] <= 15'b101011111111000;
		Coeff[7904] <= 15'b101011111111010;
		Coeff[7905] <= 15'b101011111111100;
		Coeff[7906] <= 15'b101011111111111;
		Coeff[7907] <= 15'b101100000000001;
		Coeff[7908] <= 15'b101100000000011;
		Coeff[7909] <= 15'b101100000000101;
		Coeff[7910] <= 15'b101100000001000;
		Coeff[7911] <= 15'b101100000001010;
		Coeff[7912] <= 15'b101100000001100;
		Coeff[7913] <= 15'b101100000001110;
		Coeff[7914] <= 15'b101100000010001;
		Coeff[7915] <= 15'b101100000010011;
		Coeff[7916] <= 15'b101100000010101;
		Coeff[7917] <= 15'b101100000011000;
		Coeff[7918] <= 15'b101100000011010;
		Coeff[7919] <= 15'b101100000011100;
		Coeff[7920] <= 15'b101100000011110;
		Coeff[7921] <= 15'b101100000100001;
		Coeff[7922] <= 15'b101100000100011;
		Coeff[7923] <= 15'b101100000100101;
		Coeff[7924] <= 15'b101100000101000;
		Coeff[7925] <= 15'b101100000101010;
		Coeff[7926] <= 15'b101100000101100;
		Coeff[7927] <= 15'b101100000101110;
		Coeff[7928] <= 15'b101100000110001;
		Coeff[7929] <= 15'b101100000110011;
		Coeff[7930] <= 15'b101100000110101;
		Coeff[7931] <= 15'b101100000110111;
		Coeff[7932] <= 15'b101100000111010;
		Coeff[7933] <= 15'b101100000111100;
		Coeff[7934] <= 15'b101100000111110;
		Coeff[7935] <= 15'b101100001000001;
		Coeff[7936] <= 15'b101100001000011;
		Coeff[7937] <= 15'b101100001000101;
		Coeff[7938] <= 15'b101100001000111;
		Coeff[7939] <= 15'b101100001001010;
		Coeff[7940] <= 15'b101100001001100;
		Coeff[7941] <= 15'b101100001001110;
		Coeff[7942] <= 15'b101100001010001;
		Coeff[7943] <= 15'b101100001010011;
		Coeff[7944] <= 15'b101100001010101;
		Coeff[7945] <= 15'b101100001010111;
		Coeff[7946] <= 15'b101100001011010;
		Coeff[7947] <= 15'b101100001011100;
		Coeff[7948] <= 15'b101100001011110;
		Coeff[7949] <= 15'b101100001100000;
		Coeff[7950] <= 15'b101100001100011;
		Coeff[7951] <= 15'b101100001100101;
		Coeff[7952] <= 15'b101100001100111;
		Coeff[7953] <= 15'b101100001101010;
		Coeff[7954] <= 15'b101100001101100;
		Coeff[7955] <= 15'b101100001101110;
		Coeff[7956] <= 15'b101100001110000;
		Coeff[7957] <= 15'b101100001110011;
		Coeff[7958] <= 15'b101100001110101;
		Coeff[7959] <= 15'b101100001110111;
		Coeff[7960] <= 15'b101100001111001;
		Coeff[7961] <= 15'b101100001111100;
		Coeff[7962] <= 15'b101100001111110;
		Coeff[7963] <= 15'b101100010000000;
		Coeff[7964] <= 15'b101100010000010;
		Coeff[7965] <= 15'b101100010000101;
		Coeff[7966] <= 15'b101100010000111;
		Coeff[7967] <= 15'b101100010001001;
		Coeff[7968] <= 15'b101100010001100;
		Coeff[7969] <= 15'b101100010001110;
		Coeff[7970] <= 15'b101100010010000;
		Coeff[7971] <= 15'b101100010010010;
		Coeff[7972] <= 15'b101100010010101;
		Coeff[7973] <= 15'b101100010010111;
		Coeff[7974] <= 15'b101100010011001;
		Coeff[7975] <= 15'b101100010011011;
		Coeff[7976] <= 15'b101100010011110;
		Coeff[7977] <= 15'b101100010100000;
		Coeff[7978] <= 15'b101100010100010;
		Coeff[7979] <= 15'b101100010100101;
		Coeff[7980] <= 15'b101100010100111;
		Coeff[7981] <= 15'b101100010101001;
		Coeff[7982] <= 15'b101100010101011;
		Coeff[7983] <= 15'b101100010101110;
		Coeff[7984] <= 15'b101100010110000;
		Coeff[7985] <= 15'b101100010110010;
		Coeff[7986] <= 15'b101100010110100;
		Coeff[7987] <= 15'b101100010110111;
		Coeff[7988] <= 15'b101100010111001;
		Coeff[7989] <= 15'b101100010111011;
		Coeff[7990] <= 15'b101100010111101;
		Coeff[7991] <= 15'b101100011000000;
		Coeff[7992] <= 15'b101100011000010;
		Coeff[7993] <= 15'b101100011000100;
		Coeff[7994] <= 15'b101100011000110;
		Coeff[7995] <= 15'b101100011001001;
		Coeff[7996] <= 15'b101100011001011;
		Coeff[7997] <= 15'b101100011001101;
		Coeff[7998] <= 15'b101100011010000;
		Coeff[7999] <= 15'b101100011010010;
		Coeff[8000] <= 15'b101100011010100;
		Coeff[8001] <= 15'b101100011010110;
		Coeff[8002] <= 15'b101100011011001;
		Coeff[8003] <= 15'b101100011011011;
		Coeff[8004] <= 15'b101100011011101;
		Coeff[8005] <= 15'b101100011011111;
		Coeff[8006] <= 15'b101100011100010;
		Coeff[8007] <= 15'b101100011100100;
		Coeff[8008] <= 15'b101100011100110;
		Coeff[8009] <= 15'b101100011101000;
		Coeff[8010] <= 15'b101100011101011;
		Coeff[8011] <= 15'b101100011101101;
		Coeff[8012] <= 15'b101100011101111;
		Coeff[8013] <= 15'b101100011110001;
		Coeff[8014] <= 15'b101100011110100;
		Coeff[8015] <= 15'b101100011110110;
		Coeff[8016] <= 15'b101100011111000;
		Coeff[8017] <= 15'b101100011111010;
		Coeff[8018] <= 15'b101100011111101;
		Coeff[8019] <= 15'b101100011111111;
		Coeff[8020] <= 15'b101100100000001;
		Coeff[8021] <= 15'b101100100000100;
		Coeff[8022] <= 15'b101100100000110;
		Coeff[8023] <= 15'b101100100001000;
		Coeff[8024] <= 15'b101100100001010;
		Coeff[8025] <= 15'b101100100001101;
		Coeff[8026] <= 15'b101100100001111;
		Coeff[8027] <= 15'b101100100010001;
		Coeff[8028] <= 15'b101100100010011;
		Coeff[8029] <= 15'b101100100010110;
		Coeff[8030] <= 15'b101100100011000;
		Coeff[8031] <= 15'b101100100011010;
		Coeff[8032] <= 15'b101100100011100;
		Coeff[8033] <= 15'b101100100011111;
		Coeff[8034] <= 15'b101100100100001;
		Coeff[8035] <= 15'b101100100100011;
		Coeff[8036] <= 15'b101100100100101;
		Coeff[8037] <= 15'b101100100101000;
		Coeff[8038] <= 15'b101100100101010;
		Coeff[8039] <= 15'b101100100101100;
		Coeff[8040] <= 15'b101100100101110;
		Coeff[8041] <= 15'b101100100110001;
		Coeff[8042] <= 15'b101100100110011;
		Coeff[8043] <= 15'b101100100110101;
		Coeff[8044] <= 15'b101100100110111;
		Coeff[8045] <= 15'b101100100111010;
		Coeff[8046] <= 15'b101100100111100;
		Coeff[8047] <= 15'b101100100111110;
		Coeff[8048] <= 15'b101100101000000;
		Coeff[8049] <= 15'b101100101000011;
		Coeff[8050] <= 15'b101100101000101;
		Coeff[8051] <= 15'b101100101000111;
		Coeff[8052] <= 15'b101100101001001;
		Coeff[8053] <= 15'b101100101001100;
		Coeff[8054] <= 15'b101100101001110;
		Coeff[8055] <= 15'b101100101010000;
		Coeff[8056] <= 15'b101100101010010;
		Coeff[8057] <= 15'b101100101010101;
		Coeff[8058] <= 15'b101100101010111;
		Coeff[8059] <= 15'b101100101011001;
		Coeff[8060] <= 15'b101100101011011;
		Coeff[8061] <= 15'b101100101011110;
		Coeff[8062] <= 15'b101100101100000;
		Coeff[8063] <= 15'b101100101100010;
		Coeff[8064] <= 15'b101100101100100;
		Coeff[8065] <= 15'b101100101100111;
		Coeff[8066] <= 15'b101100101101001;
		Coeff[8067] <= 15'b101100101101011;
		Coeff[8068] <= 15'b101100101101101;
		Coeff[8069] <= 15'b101100101110000;
		Coeff[8070] <= 15'b101100101110010;
		Coeff[8071] <= 15'b101100101110100;
		Coeff[8072] <= 15'b101100101110110;
		Coeff[8073] <= 15'b101100101111001;
		Coeff[8074] <= 15'b101100101111011;
		Coeff[8075] <= 15'b101100101111101;
		Coeff[8076] <= 15'b101100101111111;
		Coeff[8077] <= 15'b101100110000010;
		Coeff[8078] <= 15'b101100110000100;
		Coeff[8079] <= 15'b101100110000110;
		Coeff[8080] <= 15'b101100110001000;
		Coeff[8081] <= 15'b101100110001011;
		Coeff[8082] <= 15'b101100110001101;
		Coeff[8083] <= 15'b101100110001111;
		Coeff[8084] <= 15'b101100110010001;
		Coeff[8085] <= 15'b101100110010100;
		Coeff[8086] <= 15'b101100110010110;
		Coeff[8087] <= 15'b101100110011000;
		Coeff[8088] <= 15'b101100110011010;
		Coeff[8089] <= 15'b101100110011101;
		Coeff[8090] <= 15'b101100110011111;
		Coeff[8091] <= 15'b101100110100001;
		Coeff[8092] <= 15'b101100110100011;
		Coeff[8093] <= 15'b101100110100110;
		Coeff[8094] <= 15'b101100110101000;
		Coeff[8095] <= 15'b101100110101010;
		Coeff[8096] <= 15'b101100110101100;
		Coeff[8097] <= 15'b101100110101110;
		Coeff[8098] <= 15'b101100110110001;
		Coeff[8099] <= 15'b101100110110011;
		Coeff[8100] <= 15'b101100110110101;
		Coeff[8101] <= 15'b101100110110111;
		Coeff[8102] <= 15'b101100110111010;
		Coeff[8103] <= 15'b101100110111100;
		Coeff[8104] <= 15'b101100110111110;
		Coeff[8105] <= 15'b101100111000000;
		Coeff[8106] <= 15'b101100111000011;
		Coeff[8107] <= 15'b101100111000101;
		Coeff[8108] <= 15'b101100111000111;
		Coeff[8109] <= 15'b101100111001001;
		Coeff[8110] <= 15'b101100111001100;
		Coeff[8111] <= 15'b101100111001110;
		Coeff[8112] <= 15'b101100111010000;
		Coeff[8113] <= 15'b101100111010010;
		Coeff[8114] <= 15'b101100111010101;
		Coeff[8115] <= 15'b101100111010111;
		Coeff[8116] <= 15'b101100111011001;
		Coeff[8117] <= 15'b101100111011011;
		Coeff[8118] <= 15'b101100111011110;
		Coeff[8119] <= 15'b101100111100000;
		Coeff[8120] <= 15'b101100111100010;
		Coeff[8121] <= 15'b101100111100100;
		Coeff[8122] <= 15'b101100111100110;
		Coeff[8123] <= 15'b101100111101001;
		Coeff[8124] <= 15'b101100111101011;
		Coeff[8125] <= 15'b101100111101101;
		Coeff[8126] <= 15'b101100111101111;
		Coeff[8127] <= 15'b101100111110010;
		Coeff[8128] <= 15'b101100111110100;
		Coeff[8129] <= 15'b101100111110110;
		Coeff[8130] <= 15'b101100111111000;
		Coeff[8131] <= 15'b101100111111011;
		Coeff[8132] <= 15'b101100111111101;
		Coeff[8133] <= 15'b101100111111111;
		Coeff[8134] <= 15'b101101000000001;
		Coeff[8135] <= 15'b101101000000100;
		Coeff[8136] <= 15'b101101000000110;
		Coeff[8137] <= 15'b101101000001000;
		Coeff[8138] <= 15'b101101000001010;
		Coeff[8139] <= 15'b101101000001100;
		Coeff[8140] <= 15'b101101000001111;
		Coeff[8141] <= 15'b101101000010001;
		Coeff[8142] <= 15'b101101000010011;
		Coeff[8143] <= 15'b101101000010101;
		Coeff[8144] <= 15'b101101000011000;
		Coeff[8145] <= 15'b101101000011010;
		Coeff[8146] <= 15'b101101000011100;
		Coeff[8147] <= 15'b101101000011110;
		Coeff[8148] <= 15'b101101000100001;
		Coeff[8149] <= 15'b101101000100011;
		Coeff[8150] <= 15'b101101000100101;
		Coeff[8151] <= 15'b101101000100111;
		Coeff[8152] <= 15'b101101000101001;
		Coeff[8153] <= 15'b101101000101100;
		Coeff[8154] <= 15'b101101000101110;
		Coeff[8155] <= 15'b101101000110000;
		Coeff[8156] <= 15'b101101000110010;
		Coeff[8157] <= 15'b101101000110101;
		Coeff[8158] <= 15'b101101000110111;
		Coeff[8159] <= 15'b101101000111001;
		Coeff[8160] <= 15'b101101000111011;
		Coeff[8161] <= 15'b101101000111110;
		Coeff[8162] <= 15'b101101001000000;
		Coeff[8163] <= 15'b101101001000010;
		Coeff[8164] <= 15'b101101001000100;
		Coeff[8165] <= 15'b101101001000110;
		Coeff[8166] <= 15'b101101001001001;
		Coeff[8167] <= 15'b101101001001011;
		Coeff[8168] <= 15'b101101001001101;
		Coeff[8169] <= 15'b101101001001111;
		Coeff[8170] <= 15'b101101001010010;
		Coeff[8171] <= 15'b101101001010100;
		Coeff[8172] <= 15'b101101001010110;
		Coeff[8173] <= 15'b101101001011000;
		Coeff[8174] <= 15'b101101001011010;
		Coeff[8175] <= 15'b101101001011101;
		Coeff[8176] <= 15'b101101001011111;
		Coeff[8177] <= 15'b101101001100001;
		Coeff[8178] <= 15'b101101001100011;
		Coeff[8179] <= 15'b101101001100110;
		Coeff[8180] <= 15'b101101001101000;
		Coeff[8181] <= 15'b101101001101010;
		Coeff[8182] <= 15'b101101001101100;
		Coeff[8183] <= 15'b101101001101110;
		Coeff[8184] <= 15'b101101001110001;
		Coeff[8185] <= 15'b101101001110011;
		Coeff[8186] <= 15'b101101001110101;
		Coeff[8187] <= 15'b101101001110111;
		Coeff[8188] <= 15'b101101001111010;
		Coeff[8189] <= 15'b101101001111100;
		Coeff[8190] <= 15'b101101001111110;
		Coeff[8191] <= 15'b101101010000000;
		Coeff[8192] <= 15'b101101010000010;
		Coeff[8193] <= 15'b101101010000101;
		Coeff[8194] <= 15'b101101010000111;
		Coeff[8195] <= 15'b101101010001001;
		Coeff[8196] <= 15'b101101010001011;
		Coeff[8197] <= 15'b101101010001110;
		Coeff[8198] <= 15'b101101010010000;
		Coeff[8199] <= 15'b101101010010010;
		Coeff[8200] <= 15'b101101010010100;
		Coeff[8201] <= 15'b101101010010110;
		Coeff[8202] <= 15'b101101010011001;
		Coeff[8203] <= 15'b101101010011011;
		Coeff[8204] <= 15'b101101010011101;
		Coeff[8205] <= 15'b101101010011111;
		Coeff[8206] <= 15'b101101010100010;
		Coeff[8207] <= 15'b101101010100100;
		Coeff[8208] <= 15'b101101010100110;
		Coeff[8209] <= 15'b101101010101000;
		Coeff[8210] <= 15'b101101010101010;
		Coeff[8211] <= 15'b101101010101101;
		Coeff[8212] <= 15'b101101010101111;
		Coeff[8213] <= 15'b101101010110001;
		Coeff[8214] <= 15'b101101010110011;
		Coeff[8215] <= 15'b101101010110110;
		Coeff[8216] <= 15'b101101010111000;
		Coeff[8217] <= 15'b101101010111010;
		Coeff[8218] <= 15'b101101010111100;
		Coeff[8219] <= 15'b101101010111110;
		Coeff[8220] <= 15'b101101011000001;
		Coeff[8221] <= 15'b101101011000011;
		Coeff[8222] <= 15'b101101011000101;
		Coeff[8223] <= 15'b101101011000111;
		Coeff[8224] <= 15'b101101011001001;
		Coeff[8225] <= 15'b101101011001100;
		Coeff[8226] <= 15'b101101011001110;
		Coeff[8227] <= 15'b101101011010000;
		Coeff[8228] <= 15'b101101011010010;
		Coeff[8229] <= 15'b101101011010101;
		Coeff[8230] <= 15'b101101011010111;
		Coeff[8231] <= 15'b101101011011001;
		Coeff[8232] <= 15'b101101011011011;
		Coeff[8233] <= 15'b101101011011101;
		Coeff[8234] <= 15'b101101011100000;
		Coeff[8235] <= 15'b101101011100010;
		Coeff[8236] <= 15'b101101011100100;
		Coeff[8237] <= 15'b101101011100110;
		Coeff[8238] <= 15'b101101011101000;
		Coeff[8239] <= 15'b101101011101011;
		Coeff[8240] <= 15'b101101011101101;
		Coeff[8241] <= 15'b101101011101111;
		Coeff[8242] <= 15'b101101011110001;
		Coeff[8243] <= 15'b101101011110011;
		Coeff[8244] <= 15'b101101011110110;
		Coeff[8245] <= 15'b101101011111000;
		Coeff[8246] <= 15'b101101011111010;
		Coeff[8247] <= 15'b101101011111100;
		Coeff[8248] <= 15'b101101011111111;
		Coeff[8249] <= 15'b101101100000001;
		Coeff[8250] <= 15'b101101100000011;
		Coeff[8251] <= 15'b101101100000101;
		Coeff[8252] <= 15'b101101100000111;
		Coeff[8253] <= 15'b101101100001010;
		Coeff[8254] <= 15'b101101100001100;
		Coeff[8255] <= 15'b101101100001110;
		Coeff[8256] <= 15'b101101100010000;
		Coeff[8257] <= 15'b101101100010010;
		Coeff[8258] <= 15'b101101100010101;
		Coeff[8259] <= 15'b101101100010111;
		Coeff[8260] <= 15'b101101100011001;
		Coeff[8261] <= 15'b101101100011011;
		Coeff[8262] <= 15'b101101100011101;
		Coeff[8263] <= 15'b101101100100000;
		Coeff[8264] <= 15'b101101100100010;
		Coeff[8265] <= 15'b101101100100100;
		Coeff[8266] <= 15'b101101100100110;
		Coeff[8267] <= 15'b101101100101000;
		Coeff[8268] <= 15'b101101100101011;
		Coeff[8269] <= 15'b101101100101101;
		Coeff[8270] <= 15'b101101100101111;
		Coeff[8271] <= 15'b101101100110001;
		Coeff[8272] <= 15'b101101100110100;
		Coeff[8273] <= 15'b101101100110110;
		Coeff[8274] <= 15'b101101100111000;
		Coeff[8275] <= 15'b101101100111010;
		Coeff[8276] <= 15'b101101100111100;
		Coeff[8277] <= 15'b101101100111111;
		Coeff[8278] <= 15'b101101101000001;
		Coeff[8279] <= 15'b101101101000011;
		Coeff[8280] <= 15'b101101101000101;
		Coeff[8281] <= 15'b101101101000111;
		Coeff[8282] <= 15'b101101101001010;
		Coeff[8283] <= 15'b101101101001100;
		Coeff[8284] <= 15'b101101101001110;
		Coeff[8285] <= 15'b101101101010000;
		Coeff[8286] <= 15'b101101101010010;
		Coeff[8287] <= 15'b101101101010101;
		Coeff[8288] <= 15'b101101101010111;
		Coeff[8289] <= 15'b101101101011001;
		Coeff[8290] <= 15'b101101101011011;
		Coeff[8291] <= 15'b101101101011101;
		Coeff[8292] <= 15'b101101101100000;
		Coeff[8293] <= 15'b101101101100010;
		Coeff[8294] <= 15'b101101101100100;
		Coeff[8295] <= 15'b101101101100110;
		Coeff[8296] <= 15'b101101101101000;
		Coeff[8297] <= 15'b101101101101011;
		Coeff[8298] <= 15'b101101101101101;
		Coeff[8299] <= 15'b101101101101111;
		Coeff[8300] <= 15'b101101101110001;
		Coeff[8301] <= 15'b101101101110011;
		Coeff[8302] <= 15'b101101101110110;
		Coeff[8303] <= 15'b101101101111000;
		Coeff[8304] <= 15'b101101101111010;
		Coeff[8305] <= 15'b101101101111100;
		Coeff[8306] <= 15'b101101101111110;
		Coeff[8307] <= 15'b101101110000001;
		Coeff[8308] <= 15'b101101110000011;
		Coeff[8309] <= 15'b101101110000101;
		Coeff[8310] <= 15'b101101110000111;
		Coeff[8311] <= 15'b101101110001001;
		Coeff[8312] <= 15'b101101110001100;
		Coeff[8313] <= 15'b101101110001110;
		Coeff[8314] <= 15'b101101110010000;
		Coeff[8315] <= 15'b101101110010010;
		Coeff[8316] <= 15'b101101110010100;
		Coeff[8317] <= 15'b101101110010110;
		Coeff[8318] <= 15'b101101110011001;
		Coeff[8319] <= 15'b101101110011011;
		Coeff[8320] <= 15'b101101110011101;
		Coeff[8321] <= 15'b101101110011111;
		Coeff[8322] <= 15'b101101110100001;
		Coeff[8323] <= 15'b101101110100100;
		Coeff[8324] <= 15'b101101110100110;
		Coeff[8325] <= 15'b101101110101000;
		Coeff[8326] <= 15'b101101110101010;
		Coeff[8327] <= 15'b101101110101100;
		Coeff[8328] <= 15'b101101110101111;
		Coeff[8329] <= 15'b101101110110001;
		Coeff[8330] <= 15'b101101110110011;
		Coeff[8331] <= 15'b101101110110101;
		Coeff[8332] <= 15'b101101110110111;
		Coeff[8333] <= 15'b101101110111010;
		Coeff[8334] <= 15'b101101110111100;
		Coeff[8335] <= 15'b101101110111110;
		Coeff[8336] <= 15'b101101111000000;
		Coeff[8337] <= 15'b101101111000010;
		Coeff[8338] <= 15'b101101111000101;
		Coeff[8339] <= 15'b101101111000111;
		Coeff[8340] <= 15'b101101111001001;
		Coeff[8341] <= 15'b101101111001011;
		Coeff[8342] <= 15'b101101111001101;
		Coeff[8343] <= 15'b101101111001111;
		Coeff[8344] <= 15'b101101111010010;
		Coeff[8345] <= 15'b101101111010100;
		Coeff[8346] <= 15'b101101111010110;
		Coeff[8347] <= 15'b101101111011000;
		Coeff[8348] <= 15'b101101111011010;
		Coeff[8349] <= 15'b101101111011101;
		Coeff[8350] <= 15'b101101111011111;
		Coeff[8351] <= 15'b101101111100001;
		Coeff[8352] <= 15'b101101111100011;
		Coeff[8353] <= 15'b101101111100101;
		Coeff[8354] <= 15'b101101111101000;
		Coeff[8355] <= 15'b101101111101010;
		Coeff[8356] <= 15'b101101111101100;
		Coeff[8357] <= 15'b101101111101110;
		Coeff[8358] <= 15'b101101111110000;
		Coeff[8359] <= 15'b101101111110010;
		Coeff[8360] <= 15'b101101111110101;
		Coeff[8361] <= 15'b101101111110111;
		Coeff[8362] <= 15'b101101111111001;
		Coeff[8363] <= 15'b101101111111011;
		Coeff[8364] <= 15'b101101111111101;
		Coeff[8365] <= 15'b101110000000000;
		Coeff[8366] <= 15'b101110000000010;
		Coeff[8367] <= 15'b101110000000100;
		Coeff[8368] <= 15'b101110000000110;
		Coeff[8369] <= 15'b101110000001000;
		Coeff[8370] <= 15'b101110000001010;
		Coeff[8371] <= 15'b101110000001101;
		Coeff[8372] <= 15'b101110000001111;
		Coeff[8373] <= 15'b101110000010001;
		Coeff[8374] <= 15'b101110000010011;
		Coeff[8375] <= 15'b101110000010101;
		Coeff[8376] <= 15'b101110000011000;
		Coeff[8377] <= 15'b101110000011010;
		Coeff[8378] <= 15'b101110000011100;
		Coeff[8379] <= 15'b101110000011110;
		Coeff[8380] <= 15'b101110000100000;
		Coeff[8381] <= 15'b101110000100011;
		Coeff[8382] <= 15'b101110000100101;
		Coeff[8383] <= 15'b101110000100111;
		Coeff[8384] <= 15'b101110000101001;
		Coeff[8385] <= 15'b101110000101011;
		Coeff[8386] <= 15'b101110000101101;
		Coeff[8387] <= 15'b101110000110000;
		Coeff[8388] <= 15'b101110000110010;
		Coeff[8389] <= 15'b101110000110100;
		Coeff[8390] <= 15'b101110000110110;
		Coeff[8391] <= 15'b101110000111000;
		Coeff[8392] <= 15'b101110000111010;
		Coeff[8393] <= 15'b101110000111101;
		Coeff[8394] <= 15'b101110000111111;
		Coeff[8395] <= 15'b101110001000001;
		Coeff[8396] <= 15'b101110001000011;
		Coeff[8397] <= 15'b101110001000101;
		Coeff[8398] <= 15'b101110001001000;
		Coeff[8399] <= 15'b101110001001010;
		Coeff[8400] <= 15'b101110001001100;
		Coeff[8401] <= 15'b101110001001110;
		Coeff[8402] <= 15'b101110001010000;
		Coeff[8403] <= 15'b101110001010010;
		Coeff[8404] <= 15'b101110001010101;
		Coeff[8405] <= 15'b101110001010111;
		Coeff[8406] <= 15'b101110001011001;
		Coeff[8407] <= 15'b101110001011011;
		Coeff[8408] <= 15'b101110001011101;
		Coeff[8409] <= 15'b101110001011111;
		Coeff[8410] <= 15'b101110001100010;
		Coeff[8411] <= 15'b101110001100100;
		Coeff[8412] <= 15'b101110001100110;
		Coeff[8413] <= 15'b101110001101000;
		Coeff[8414] <= 15'b101110001101010;
		Coeff[8415] <= 15'b101110001101101;
		Coeff[8416] <= 15'b101110001101111;
		Coeff[8417] <= 15'b101110001110001;
		Coeff[8418] <= 15'b101110001110011;
		Coeff[8419] <= 15'b101110001110101;
		Coeff[8420] <= 15'b101110001110111;
		Coeff[8421] <= 15'b101110001111010;
		Coeff[8422] <= 15'b101110001111100;
		Coeff[8423] <= 15'b101110001111110;
		Coeff[8424] <= 15'b101110010000000;
		Coeff[8425] <= 15'b101110010000010;
		Coeff[8426] <= 15'b101110010000100;
		Coeff[8427] <= 15'b101110010000111;
		Coeff[8428] <= 15'b101110010001001;
		Coeff[8429] <= 15'b101110010001011;
		Coeff[8430] <= 15'b101110010001101;
		Coeff[8431] <= 15'b101110010001111;
		Coeff[8432] <= 15'b101110010010001;
		Coeff[8433] <= 15'b101110010010100;
		Coeff[8434] <= 15'b101110010010110;
		Coeff[8435] <= 15'b101110010011000;
		Coeff[8436] <= 15'b101110010011010;
		Coeff[8437] <= 15'b101110010011100;
		Coeff[8438] <= 15'b101110010011110;
		Coeff[8439] <= 15'b101110010100001;
		Coeff[8440] <= 15'b101110010100011;
		Coeff[8441] <= 15'b101110010100101;
		Coeff[8442] <= 15'b101110010100111;
		Coeff[8443] <= 15'b101110010101001;
		Coeff[8444] <= 15'b101110010101011;
		Coeff[8445] <= 15'b101110010101110;
		Coeff[8446] <= 15'b101110010110000;
		Coeff[8447] <= 15'b101110010110010;
		Coeff[8448] <= 15'b101110010110100;
		Coeff[8449] <= 15'b101110010110110;
		Coeff[8450] <= 15'b101110010111000;
		Coeff[8451] <= 15'b101110010111011;
		Coeff[8452] <= 15'b101110010111101;
		Coeff[8453] <= 15'b101110010111111;
		Coeff[8454] <= 15'b101110011000001;
		Coeff[8455] <= 15'b101110011000011;
		Coeff[8456] <= 15'b101110011000101;
		Coeff[8457] <= 15'b101110011001000;
		Coeff[8458] <= 15'b101110011001010;
		Coeff[8459] <= 15'b101110011001100;
		Coeff[8460] <= 15'b101110011001110;
		Coeff[8461] <= 15'b101110011010000;
		Coeff[8462] <= 15'b101110011010010;
		Coeff[8463] <= 15'b101110011010101;
		Coeff[8464] <= 15'b101110011010111;
		Coeff[8465] <= 15'b101110011011001;
		Coeff[8466] <= 15'b101110011011011;
		Coeff[8467] <= 15'b101110011011101;
		Coeff[8468] <= 15'b101110011011111;
		Coeff[8469] <= 15'b101110011100010;
		Coeff[8470] <= 15'b101110011100100;
		Coeff[8471] <= 15'b101110011100110;
		Coeff[8472] <= 15'b101110011101000;
		Coeff[8473] <= 15'b101110011101010;
		Coeff[8474] <= 15'b101110011101100;
		Coeff[8475] <= 15'b101110011101111;
		Coeff[8476] <= 15'b101110011110001;
		Coeff[8477] <= 15'b101110011110011;
		Coeff[8478] <= 15'b101110011110101;
		Coeff[8479] <= 15'b101110011110111;
		Coeff[8480] <= 15'b101110011111001;
		Coeff[8481] <= 15'b101110011111011;
		Coeff[8482] <= 15'b101110011111110;
		Coeff[8483] <= 15'b101110100000000;
		Coeff[8484] <= 15'b101110100000010;
		Coeff[8485] <= 15'b101110100000100;
		Coeff[8486] <= 15'b101110100000110;
		Coeff[8487] <= 15'b101110100001000;
		Coeff[8488] <= 15'b101110100001011;
		Coeff[8489] <= 15'b101110100001101;
		Coeff[8490] <= 15'b101110100001111;
		Coeff[8491] <= 15'b101110100010001;
		Coeff[8492] <= 15'b101110100010011;
		Coeff[8493] <= 15'b101110100010101;
		Coeff[8494] <= 15'b101110100011000;
		Coeff[8495] <= 15'b101110100011010;
		Coeff[8496] <= 15'b101110100011100;
		Coeff[8497] <= 15'b101110100011110;
		Coeff[8498] <= 15'b101110100100000;
		Coeff[8499] <= 15'b101110100100010;
		Coeff[8500] <= 15'b101110100100100;
		Coeff[8501] <= 15'b101110100100111;
		Coeff[8502] <= 15'b101110100101001;
		Coeff[8503] <= 15'b101110100101011;
		Coeff[8504] <= 15'b101110100101101;
		Coeff[8505] <= 15'b101110100101111;
		Coeff[8506] <= 15'b101110100110001;
		Coeff[8507] <= 15'b101110100110100;
		Coeff[8508] <= 15'b101110100110110;
		Coeff[8509] <= 15'b101110100111000;
		Coeff[8510] <= 15'b101110100111010;
		Coeff[8511] <= 15'b101110100111100;
		Coeff[8512] <= 15'b101110100111110;
		Coeff[8513] <= 15'b101110101000000;
		Coeff[8514] <= 15'b101110101000011;
		Coeff[8515] <= 15'b101110101000101;
		Coeff[8516] <= 15'b101110101000111;
		Coeff[8517] <= 15'b101110101001001;
		Coeff[8518] <= 15'b101110101001011;
		Coeff[8519] <= 15'b101110101001101;
		Coeff[8520] <= 15'b101110101010000;
		Coeff[8521] <= 15'b101110101010010;
		Coeff[8522] <= 15'b101110101010100;
		Coeff[8523] <= 15'b101110101010110;
		Coeff[8524] <= 15'b101110101011000;
		Coeff[8525] <= 15'b101110101011010;
		Coeff[8526] <= 15'b101110101011100;
		Coeff[8527] <= 15'b101110101011111;
		Coeff[8528] <= 15'b101110101100001;
		Coeff[8529] <= 15'b101110101100011;
		Coeff[8530] <= 15'b101110101100101;
		Coeff[8531] <= 15'b101110101100111;
		Coeff[8532] <= 15'b101110101101001;
		Coeff[8533] <= 15'b101110101101011;
		Coeff[8534] <= 15'b101110101101110;
		Coeff[8535] <= 15'b101110101110000;
		Coeff[8536] <= 15'b101110101110010;
		Coeff[8537] <= 15'b101110101110100;
		Coeff[8538] <= 15'b101110101110110;
		Coeff[8539] <= 15'b101110101111000;
		Coeff[8540] <= 15'b101110101111010;
		Coeff[8541] <= 15'b101110101111101;
		Coeff[8542] <= 15'b101110101111111;
		Coeff[8543] <= 15'b101110110000001;
		Coeff[8544] <= 15'b101110110000011;
		Coeff[8545] <= 15'b101110110000101;
		Coeff[8546] <= 15'b101110110000111;
		Coeff[8547] <= 15'b101110110001010;
		Coeff[8548] <= 15'b101110110001100;
		Coeff[8549] <= 15'b101110110001110;
		Coeff[8550] <= 15'b101110110010000;
		Coeff[8551] <= 15'b101110110010010;
		Coeff[8552] <= 15'b101110110010100;
		Coeff[8553] <= 15'b101110110010110;
		Coeff[8554] <= 15'b101110110011001;
		Coeff[8555] <= 15'b101110110011011;
		Coeff[8556] <= 15'b101110110011101;
		Coeff[8557] <= 15'b101110110011111;
		Coeff[8558] <= 15'b101110110100001;
		Coeff[8559] <= 15'b101110110100011;
		Coeff[8560] <= 15'b101110110100101;
		Coeff[8561] <= 15'b101110110101000;
		Coeff[8562] <= 15'b101110110101010;
		Coeff[8563] <= 15'b101110110101100;
		Coeff[8564] <= 15'b101110110101110;
		Coeff[8565] <= 15'b101110110110000;
		Coeff[8566] <= 15'b101110110110010;
		Coeff[8567] <= 15'b101110110110100;
		Coeff[8568] <= 15'b101110110110111;
		Coeff[8569] <= 15'b101110110111001;
		Coeff[8570] <= 15'b101110110111011;
		Coeff[8571] <= 15'b101110110111101;
		Coeff[8572] <= 15'b101110110111111;
		Coeff[8573] <= 15'b101110111000001;
		Coeff[8574] <= 15'b101110111000011;
		Coeff[8575] <= 15'b101110111000101;
		Coeff[8576] <= 15'b101110111001000;
		Coeff[8577] <= 15'b101110111001010;
		Coeff[8578] <= 15'b101110111001100;
		Coeff[8579] <= 15'b101110111001110;
		Coeff[8580] <= 15'b101110111010000;
		Coeff[8581] <= 15'b101110111010010;
		Coeff[8582] <= 15'b101110111010100;
		Coeff[8583] <= 15'b101110111010111;
		Coeff[8584] <= 15'b101110111011001;
		Coeff[8585] <= 15'b101110111011011;
		Coeff[8586] <= 15'b101110111011101;
		Coeff[8587] <= 15'b101110111011111;
		Coeff[8588] <= 15'b101110111100001;
		Coeff[8589] <= 15'b101110111100011;
		Coeff[8590] <= 15'b101110111100110;
		Coeff[8591] <= 15'b101110111101000;
		Coeff[8592] <= 15'b101110111101010;
		Coeff[8593] <= 15'b101110111101100;
		Coeff[8594] <= 15'b101110111101110;
		Coeff[8595] <= 15'b101110111110000;
		Coeff[8596] <= 15'b101110111110010;
		Coeff[8597] <= 15'b101110111110100;
		Coeff[8598] <= 15'b101110111110111;
		Coeff[8599] <= 15'b101110111111001;
		Coeff[8600] <= 15'b101110111111011;
		Coeff[8601] <= 15'b101110111111101;
		Coeff[8602] <= 15'b101110111111111;
		Coeff[8603] <= 15'b101111000000001;
		Coeff[8604] <= 15'b101111000000011;
		Coeff[8605] <= 15'b101111000000110;
		Coeff[8606] <= 15'b101111000001000;
		Coeff[8607] <= 15'b101111000001010;
		Coeff[8608] <= 15'b101111000001100;
		Coeff[8609] <= 15'b101111000001110;
		Coeff[8610] <= 15'b101111000010000;
		Coeff[8611] <= 15'b101111000010010;
		Coeff[8612] <= 15'b101111000010100;
		Coeff[8613] <= 15'b101111000010111;
		Coeff[8614] <= 15'b101111000011001;
		Coeff[8615] <= 15'b101111000011011;
		Coeff[8616] <= 15'b101111000011101;
		Coeff[8617] <= 15'b101111000011111;
		Coeff[8618] <= 15'b101111000100001;
		Coeff[8619] <= 15'b101111000100011;
		Coeff[8620] <= 15'b101111000100101;
		Coeff[8621] <= 15'b101111000101000;
		Coeff[8622] <= 15'b101111000101010;
		Coeff[8623] <= 15'b101111000101100;
		Coeff[8624] <= 15'b101111000101110;
		Coeff[8625] <= 15'b101111000110000;
		Coeff[8626] <= 15'b101111000110010;
		Coeff[8627] <= 15'b101111000110100;
		Coeff[8628] <= 15'b101111000110111;
		Coeff[8629] <= 15'b101111000111001;
		Coeff[8630] <= 15'b101111000111011;
		Coeff[8631] <= 15'b101111000111101;
		Coeff[8632] <= 15'b101111000111111;
		Coeff[8633] <= 15'b101111001000001;
		Coeff[8634] <= 15'b101111001000011;
		Coeff[8635] <= 15'b101111001000101;
		Coeff[8636] <= 15'b101111001001000;
		Coeff[8637] <= 15'b101111001001010;
		Coeff[8638] <= 15'b101111001001100;
		Coeff[8639] <= 15'b101111001001110;
		Coeff[8640] <= 15'b101111001010000;
		Coeff[8641] <= 15'b101111001010010;
		Coeff[8642] <= 15'b101111001010100;
		Coeff[8643] <= 15'b101111001010110;
		Coeff[8644] <= 15'b101111001011000;
		Coeff[8645] <= 15'b101111001011011;
		Coeff[8646] <= 15'b101111001011101;
		Coeff[8647] <= 15'b101111001011111;
		Coeff[8648] <= 15'b101111001100001;
		Coeff[8649] <= 15'b101111001100011;
		Coeff[8650] <= 15'b101111001100101;
		Coeff[8651] <= 15'b101111001100111;
		Coeff[8652] <= 15'b101111001101001;
		Coeff[8653] <= 15'b101111001101100;
		Coeff[8654] <= 15'b101111001101110;
		Coeff[8655] <= 15'b101111001110000;
		Coeff[8656] <= 15'b101111001110010;
		Coeff[8657] <= 15'b101111001110100;
		Coeff[8658] <= 15'b101111001110110;
		Coeff[8659] <= 15'b101111001111000;
		Coeff[8660] <= 15'b101111001111010;
		Coeff[8661] <= 15'b101111001111101;
		Coeff[8662] <= 15'b101111001111111;
		Coeff[8663] <= 15'b101111010000001;
		Coeff[8664] <= 15'b101111010000011;
		Coeff[8665] <= 15'b101111010000101;
		Coeff[8666] <= 15'b101111010000111;
		Coeff[8667] <= 15'b101111010001001;
		Coeff[8668] <= 15'b101111010001011;
		Coeff[8669] <= 15'b101111010001110;
		Coeff[8670] <= 15'b101111010010000;
		Coeff[8671] <= 15'b101111010010010;
		Coeff[8672] <= 15'b101111010010100;
		Coeff[8673] <= 15'b101111010010110;
		Coeff[8674] <= 15'b101111010011000;
		Coeff[8675] <= 15'b101111010011010;
		Coeff[8676] <= 15'b101111010011100;
		Coeff[8677] <= 15'b101111010011110;
		Coeff[8678] <= 15'b101111010100001;
		Coeff[8679] <= 15'b101111010100011;
		Coeff[8680] <= 15'b101111010100101;
		Coeff[8681] <= 15'b101111010100111;
		Coeff[8682] <= 15'b101111010101001;
		Coeff[8683] <= 15'b101111010101011;
		Coeff[8684] <= 15'b101111010101101;
		Coeff[8685] <= 15'b101111010101111;
		Coeff[8686] <= 15'b101111010110001;
		Coeff[8687] <= 15'b101111010110100;
		Coeff[8688] <= 15'b101111010110110;
		Coeff[8689] <= 15'b101111010111000;
		Coeff[8690] <= 15'b101111010111010;
		Coeff[8691] <= 15'b101111010111100;
		Coeff[8692] <= 15'b101111010111110;
		Coeff[8693] <= 15'b101111011000000;
		Coeff[8694] <= 15'b101111011000010;
		Coeff[8695] <= 15'b101111011000100;
		Coeff[8696] <= 15'b101111011000111;
		Coeff[8697] <= 15'b101111011001001;
		Coeff[8698] <= 15'b101111011001011;
		Coeff[8699] <= 15'b101111011001101;
		Coeff[8700] <= 15'b101111011001111;
		Coeff[8701] <= 15'b101111011010001;
		Coeff[8702] <= 15'b101111011010011;
		Coeff[8703] <= 15'b101111011010101;
		Coeff[8704] <= 15'b101111011010111;
		Coeff[8705] <= 15'b101111011011010;
		Coeff[8706] <= 15'b101111011011100;
		Coeff[8707] <= 15'b101111011011110;
		Coeff[8708] <= 15'b101111011100000;
		Coeff[8709] <= 15'b101111011100010;
		Coeff[8710] <= 15'b101111011100100;
		Coeff[8711] <= 15'b101111011100110;
		Coeff[8712] <= 15'b101111011101000;
		Coeff[8713] <= 15'b101111011101010;
		Coeff[8714] <= 15'b101111011101101;
		Coeff[8715] <= 15'b101111011101111;
		Coeff[8716] <= 15'b101111011110001;
		Coeff[8717] <= 15'b101111011110011;
		Coeff[8718] <= 15'b101111011110101;
		Coeff[8719] <= 15'b101111011110111;
		Coeff[8720] <= 15'b101111011111001;
		Coeff[8721] <= 15'b101111011111011;
		Coeff[8722] <= 15'b101111011111101;
		Coeff[8723] <= 15'b101111100000000;
		Coeff[8724] <= 15'b101111100000010;
		Coeff[8725] <= 15'b101111100000100;
		Coeff[8726] <= 15'b101111100000110;
		Coeff[8727] <= 15'b101111100001000;
		Coeff[8728] <= 15'b101111100001010;
		Coeff[8729] <= 15'b101111100001100;
		Coeff[8730] <= 15'b101111100001110;
		Coeff[8731] <= 15'b101111100010000;
		Coeff[8732] <= 15'b101111100010010;
		Coeff[8733] <= 15'b101111100010101;
		Coeff[8734] <= 15'b101111100010111;
		Coeff[8735] <= 15'b101111100011001;
		Coeff[8736] <= 15'b101111100011011;
		Coeff[8737] <= 15'b101111100011101;
		Coeff[8738] <= 15'b101111100011111;
		Coeff[8739] <= 15'b101111100100001;
		Coeff[8740] <= 15'b101111100100011;
		Coeff[8741] <= 15'b101111100100101;
		Coeff[8742] <= 15'b101111100100111;
		Coeff[8743] <= 15'b101111100101010;
		Coeff[8744] <= 15'b101111100101100;
		Coeff[8745] <= 15'b101111100101110;
		Coeff[8746] <= 15'b101111100110000;
		Coeff[8747] <= 15'b101111100110010;
		Coeff[8748] <= 15'b101111100110100;
		Coeff[8749] <= 15'b101111100110110;
		Coeff[8750] <= 15'b101111100111000;
		Coeff[8751] <= 15'b101111100111010;
		Coeff[8752] <= 15'b101111100111100;
		Coeff[8753] <= 15'b101111100111111;
		Coeff[8754] <= 15'b101111101000001;
		Coeff[8755] <= 15'b101111101000011;
		Coeff[8756] <= 15'b101111101000101;
		Coeff[8757] <= 15'b101111101000111;
		Coeff[8758] <= 15'b101111101001001;
		Coeff[8759] <= 15'b101111101001011;
		Coeff[8760] <= 15'b101111101001101;
		Coeff[8761] <= 15'b101111101001111;
		Coeff[8762] <= 15'b101111101010001;
		Coeff[8763] <= 15'b101111101010100;
		Coeff[8764] <= 15'b101111101010110;
		Coeff[8765] <= 15'b101111101011000;
		Coeff[8766] <= 15'b101111101011010;
		Coeff[8767] <= 15'b101111101011100;
		Coeff[8768] <= 15'b101111101011110;
		Coeff[8769] <= 15'b101111101100000;
		Coeff[8770] <= 15'b101111101100010;
		Coeff[8771] <= 15'b101111101100100;
		Coeff[8772] <= 15'b101111101100110;
		Coeff[8773] <= 15'b101111101101001;
		Coeff[8774] <= 15'b101111101101011;
		Coeff[8775] <= 15'b101111101101101;
		Coeff[8776] <= 15'b101111101101111;
		Coeff[8777] <= 15'b101111101110001;
		Coeff[8778] <= 15'b101111101110011;
		Coeff[8779] <= 15'b101111101110101;
		Coeff[8780] <= 15'b101111101110111;
		Coeff[8781] <= 15'b101111101111001;
		Coeff[8782] <= 15'b101111101111011;
		Coeff[8783] <= 15'b101111101111101;
		Coeff[8784] <= 15'b101111110000000;
		Coeff[8785] <= 15'b101111110000010;
		Coeff[8786] <= 15'b101111110000100;
		Coeff[8787] <= 15'b101111110000110;
		Coeff[8788] <= 15'b101111110001000;
		Coeff[8789] <= 15'b101111110001010;
		Coeff[8790] <= 15'b101111110001100;
		Coeff[8791] <= 15'b101111110001110;
		Coeff[8792] <= 15'b101111110010000;
		Coeff[8793] <= 15'b101111110010010;
		Coeff[8794] <= 15'b101111110010100;
		Coeff[8795] <= 15'b101111110010111;
		Coeff[8796] <= 15'b101111110011001;
		Coeff[8797] <= 15'b101111110011011;
		Coeff[8798] <= 15'b101111110011101;
		Coeff[8799] <= 15'b101111110011111;
		Coeff[8800] <= 15'b101111110100001;
		Coeff[8801] <= 15'b101111110100011;
		Coeff[8802] <= 15'b101111110100101;
		Coeff[8803] <= 15'b101111110100111;
		Coeff[8804] <= 15'b101111110101001;
		Coeff[8805] <= 15'b101111110101011;
		Coeff[8806] <= 15'b101111110101110;
		Coeff[8807] <= 15'b101111110110000;
		Coeff[8808] <= 15'b101111110110010;
		Coeff[8809] <= 15'b101111110110100;
		Coeff[8810] <= 15'b101111110110110;
		Coeff[8811] <= 15'b101111110111000;
		Coeff[8812] <= 15'b101111110111010;
		Coeff[8813] <= 15'b101111110111100;
		Coeff[8814] <= 15'b101111110111110;
		Coeff[8815] <= 15'b101111111000000;
		Coeff[8816] <= 15'b101111111000010;
		Coeff[8817] <= 15'b101111111000100;
		Coeff[8818] <= 15'b101111111000111;
		Coeff[8819] <= 15'b101111111001001;
		Coeff[8820] <= 15'b101111111001011;
		Coeff[8821] <= 15'b101111111001101;
		Coeff[8822] <= 15'b101111111001111;
		Coeff[8823] <= 15'b101111111010001;
		Coeff[8824] <= 15'b101111111010011;
		Coeff[8825] <= 15'b101111111010101;
		Coeff[8826] <= 15'b101111111010111;
		Coeff[8827] <= 15'b101111111011001;
		Coeff[8828] <= 15'b101111111011011;
		Coeff[8829] <= 15'b101111111011101;
		Coeff[8830] <= 15'b101111111100000;
		Coeff[8831] <= 15'b101111111100010;
		Coeff[8832] <= 15'b101111111100100;
		Coeff[8833] <= 15'b101111111100110;
		Coeff[8834] <= 15'b101111111101000;
		Coeff[8835] <= 15'b101111111101010;
		Coeff[8836] <= 15'b101111111101100;
		Coeff[8837] <= 15'b101111111101110;
		Coeff[8838] <= 15'b101111111110000;
		Coeff[8839] <= 15'b101111111110010;
		Coeff[8840] <= 15'b101111111110100;
		Coeff[8841] <= 15'b101111111110110;
		Coeff[8842] <= 15'b101111111111001;
		Coeff[8843] <= 15'b101111111111011;
		Coeff[8844] <= 15'b101111111111101;
		Coeff[8845] <= 15'b101111111111111;
		Coeff[8846] <= 15'b110000000000001;
		Coeff[8847] <= 15'b110000000000011;
		Coeff[8848] <= 15'b110000000000101;
		Coeff[8849] <= 15'b110000000000111;
		Coeff[8850] <= 15'b110000000001001;
		Coeff[8851] <= 15'b110000000001011;
		Coeff[8852] <= 15'b110000000001101;
		Coeff[8853] <= 15'b110000000001111;
		Coeff[8854] <= 15'b110000000010001;
		Coeff[8855] <= 15'b110000000010100;
		Coeff[8856] <= 15'b110000000010110;
		Coeff[8857] <= 15'b110000000011000;
		Coeff[8858] <= 15'b110000000011010;
		Coeff[8859] <= 15'b110000000011100;
		Coeff[8860] <= 15'b110000000011110;
		Coeff[8861] <= 15'b110000000100000;
		Coeff[8862] <= 15'b110000000100010;
		Coeff[8863] <= 15'b110000000100100;
		Coeff[8864] <= 15'b110000000100110;
		Coeff[8865] <= 15'b110000000101000;
		Coeff[8866] <= 15'b110000000101010;
		Coeff[8867] <= 15'b110000000101100;
		Coeff[8868] <= 15'b110000000101110;
		Coeff[8869] <= 15'b110000000110001;
		Coeff[8870] <= 15'b110000000110011;
		Coeff[8871] <= 15'b110000000110101;
		Coeff[8872] <= 15'b110000000110111;
		Coeff[8873] <= 15'b110000000111001;
		Coeff[8874] <= 15'b110000000111011;
		Coeff[8875] <= 15'b110000000111101;
		Coeff[8876] <= 15'b110000000111111;
		Coeff[8877] <= 15'b110000001000001;
		Coeff[8878] <= 15'b110000001000011;
		Coeff[8879] <= 15'b110000001000101;
		Coeff[8880] <= 15'b110000001000111;
		Coeff[8881] <= 15'b110000001001001;
		Coeff[8882] <= 15'b110000001001011;
		Coeff[8883] <= 15'b110000001001110;
		Coeff[8884] <= 15'b110000001010000;
		Coeff[8885] <= 15'b110000001010010;
		Coeff[8886] <= 15'b110000001010100;
		Coeff[8887] <= 15'b110000001010110;
		Coeff[8888] <= 15'b110000001011000;
		Coeff[8889] <= 15'b110000001011010;
		Coeff[8890] <= 15'b110000001011100;
		Coeff[8891] <= 15'b110000001011110;
		Coeff[8892] <= 15'b110000001100000;
		Coeff[8893] <= 15'b110000001100010;
		Coeff[8894] <= 15'b110000001100100;
		Coeff[8895] <= 15'b110000001100110;
		Coeff[8896] <= 15'b110000001101000;
		Coeff[8897] <= 15'b110000001101010;
		Coeff[8898] <= 15'b110000001101101;
		Coeff[8899] <= 15'b110000001101111;
		Coeff[8900] <= 15'b110000001110001;
		Coeff[8901] <= 15'b110000001110011;
		Coeff[8902] <= 15'b110000001110101;
		Coeff[8903] <= 15'b110000001110111;
		Coeff[8904] <= 15'b110000001111001;
		Coeff[8905] <= 15'b110000001111011;
		Coeff[8906] <= 15'b110000001111101;
		Coeff[8907] <= 15'b110000001111111;
		Coeff[8908] <= 15'b110000010000001;
		Coeff[8909] <= 15'b110000010000011;
		Coeff[8910] <= 15'b110000010000101;
		Coeff[8911] <= 15'b110000010000111;
		Coeff[8912] <= 15'b110000010001001;
		Coeff[8913] <= 15'b110000010001100;
		Coeff[8914] <= 15'b110000010001110;
		Coeff[8915] <= 15'b110000010010000;
		Coeff[8916] <= 15'b110000010010010;
		Coeff[8917] <= 15'b110000010010100;
		Coeff[8918] <= 15'b110000010010110;
		Coeff[8919] <= 15'b110000010011000;
		Coeff[8920] <= 15'b110000010011010;
		Coeff[8921] <= 15'b110000010011100;
		Coeff[8922] <= 15'b110000010011110;
		Coeff[8923] <= 15'b110000010100000;
		Coeff[8924] <= 15'b110000010100010;
		Coeff[8925] <= 15'b110000010100100;
		Coeff[8926] <= 15'b110000010100110;
		Coeff[8927] <= 15'b110000010101000;
		Coeff[8928] <= 15'b110000010101010;
		Coeff[8929] <= 15'b110000010101100;
		Coeff[8930] <= 15'b110000010101111;
		Coeff[8931] <= 15'b110000010110001;
		Coeff[8932] <= 15'b110000010110011;
		Coeff[8933] <= 15'b110000010110101;
		Coeff[8934] <= 15'b110000010110111;
		Coeff[8935] <= 15'b110000010111001;
		Coeff[8936] <= 15'b110000010111011;
		Coeff[8937] <= 15'b110000010111101;
		Coeff[8938] <= 15'b110000010111111;
		Coeff[8939] <= 15'b110000011000001;
		Coeff[8940] <= 15'b110000011000011;
		Coeff[8941] <= 15'b110000011000101;
		Coeff[8942] <= 15'b110000011000111;
		Coeff[8943] <= 15'b110000011001001;
		Coeff[8944] <= 15'b110000011001011;
		Coeff[8945] <= 15'b110000011001101;
		Coeff[8946] <= 15'b110000011001111;
		Coeff[8947] <= 15'b110000011010010;
		Coeff[8948] <= 15'b110000011010100;
		Coeff[8949] <= 15'b110000011010110;
		Coeff[8950] <= 15'b110000011011000;
		Coeff[8951] <= 15'b110000011011010;
		Coeff[8952] <= 15'b110000011011100;
		Coeff[8953] <= 15'b110000011011110;
		Coeff[8954] <= 15'b110000011100000;
		Coeff[8955] <= 15'b110000011100010;
		Coeff[8956] <= 15'b110000011100100;
		Coeff[8957] <= 15'b110000011100110;
		Coeff[8958] <= 15'b110000011101000;
		Coeff[8959] <= 15'b110000011101010;
		Coeff[8960] <= 15'b110000011101100;
		Coeff[8961] <= 15'b110000011101110;
		Coeff[8962] <= 15'b110000011110000;
		Coeff[8963] <= 15'b110000011110010;
		Coeff[8964] <= 15'b110000011110100;
		Coeff[8965] <= 15'b110000011110110;
		Coeff[8966] <= 15'b110000011111001;
		Coeff[8967] <= 15'b110000011111011;
		Coeff[8968] <= 15'b110000011111101;
		Coeff[8969] <= 15'b110000011111111;
		Coeff[8970] <= 15'b110000100000001;
		Coeff[8971] <= 15'b110000100000011;
		Coeff[8972] <= 15'b110000100000101;
		Coeff[8973] <= 15'b110000100000111;
		Coeff[8974] <= 15'b110000100001001;
		Coeff[8975] <= 15'b110000100001011;
		Coeff[8976] <= 15'b110000100001101;
		Coeff[8977] <= 15'b110000100001111;
		Coeff[8978] <= 15'b110000100010001;
		Coeff[8979] <= 15'b110000100010011;
		Coeff[8980] <= 15'b110000100010101;
		Coeff[8981] <= 15'b110000100010111;
		Coeff[8982] <= 15'b110000100011001;
		Coeff[8983] <= 15'b110000100011011;
		Coeff[8984] <= 15'b110000100011101;
		Coeff[8985] <= 15'b110000100011111;
		Coeff[8986] <= 15'b110000100100001;
		Coeff[8987] <= 15'b110000100100100;
		Coeff[8988] <= 15'b110000100100110;
		Coeff[8989] <= 15'b110000100101000;
		Coeff[8990] <= 15'b110000100101010;
		Coeff[8991] <= 15'b110000100101100;
		Coeff[8992] <= 15'b110000100101110;
		Coeff[8993] <= 15'b110000100110000;
		Coeff[8994] <= 15'b110000100110010;
		Coeff[8995] <= 15'b110000100110100;
		Coeff[8996] <= 15'b110000100110110;
		Coeff[8997] <= 15'b110000100111000;
		Coeff[8998] <= 15'b110000100111010;
		Coeff[8999] <= 15'b110000100111100;
		Coeff[9000] <= 15'b110000100111110;
		Coeff[9001] <= 15'b110000101000000;
		Coeff[9002] <= 15'b110000101000010;
		Coeff[9003] <= 15'b110000101000100;
		Coeff[9004] <= 15'b110000101000110;
		Coeff[9005] <= 15'b110000101001000;
		Coeff[9006] <= 15'b110000101001010;
		Coeff[9007] <= 15'b110000101001100;
		Coeff[9008] <= 15'b110000101001110;
		Coeff[9009] <= 15'b110000101010000;
		Coeff[9010] <= 15'b110000101010011;
		Coeff[9011] <= 15'b110000101010101;
		Coeff[9012] <= 15'b110000101010111;
		Coeff[9013] <= 15'b110000101011001;
		Coeff[9014] <= 15'b110000101011011;
		Coeff[9015] <= 15'b110000101011101;
		Coeff[9016] <= 15'b110000101011111;
		Coeff[9017] <= 15'b110000101100001;
		Coeff[9018] <= 15'b110000101100011;
		Coeff[9019] <= 15'b110000101100101;
		Coeff[9020] <= 15'b110000101100111;
		Coeff[9021] <= 15'b110000101101001;
		Coeff[9022] <= 15'b110000101101011;
		Coeff[9023] <= 15'b110000101101101;
		Coeff[9024] <= 15'b110000101101111;
		Coeff[9025] <= 15'b110000101110001;
		Coeff[9026] <= 15'b110000101110011;
		Coeff[9027] <= 15'b110000101110101;
		Coeff[9028] <= 15'b110000101110111;
		Coeff[9029] <= 15'b110000101111001;
		Coeff[9030] <= 15'b110000101111011;
		Coeff[9031] <= 15'b110000101111101;
		Coeff[9032] <= 15'b110000101111111;
		Coeff[9033] <= 15'b110000110000001;
		Coeff[9034] <= 15'b110000110000011;
		Coeff[9035] <= 15'b110000110000101;
		Coeff[9036] <= 15'b110000110001000;
		Coeff[9037] <= 15'b110000110001010;
		Coeff[9038] <= 15'b110000110001100;
		Coeff[9039] <= 15'b110000110001110;
		Coeff[9040] <= 15'b110000110010000;
		Coeff[9041] <= 15'b110000110010010;
		Coeff[9042] <= 15'b110000110010100;
		Coeff[9043] <= 15'b110000110010110;
		Coeff[9044] <= 15'b110000110011000;
		Coeff[9045] <= 15'b110000110011010;
		Coeff[9046] <= 15'b110000110011100;
		Coeff[9047] <= 15'b110000110011110;
		Coeff[9048] <= 15'b110000110100000;
		Coeff[9049] <= 15'b110000110100010;
		Coeff[9050] <= 15'b110000110100100;
		Coeff[9051] <= 15'b110000110100110;
		Coeff[9052] <= 15'b110000110101000;
		Coeff[9053] <= 15'b110000110101010;
		Coeff[9054] <= 15'b110000110101100;
		Coeff[9055] <= 15'b110000110101110;
		Coeff[9056] <= 15'b110000110110000;
		Coeff[9057] <= 15'b110000110110010;
		Coeff[9058] <= 15'b110000110110100;
		Coeff[9059] <= 15'b110000110110110;
		Coeff[9060] <= 15'b110000110111000;
		Coeff[9061] <= 15'b110000110111010;
		Coeff[9062] <= 15'b110000110111100;
		Coeff[9063] <= 15'b110000110111110;
		Coeff[9064] <= 15'b110000111000000;
		Coeff[9065] <= 15'b110000111000010;
		Coeff[9066] <= 15'b110000111000100;
		Coeff[9067] <= 15'b110000111000110;
		Coeff[9068] <= 15'b110000111001001;
		Coeff[9069] <= 15'b110000111001011;
		Coeff[9070] <= 15'b110000111001101;
		Coeff[9071] <= 15'b110000111001111;
		Coeff[9072] <= 15'b110000111010001;
		Coeff[9073] <= 15'b110000111010011;
		Coeff[9074] <= 15'b110000111010101;
		Coeff[9075] <= 15'b110000111010111;
		Coeff[9076] <= 15'b110000111011001;
		Coeff[9077] <= 15'b110000111011011;
		Coeff[9078] <= 15'b110000111011101;
		Coeff[9079] <= 15'b110000111011111;
		Coeff[9080] <= 15'b110000111100001;
		Coeff[9081] <= 15'b110000111100011;
		Coeff[9082] <= 15'b110000111100101;
		Coeff[9083] <= 15'b110000111100111;
		Coeff[9084] <= 15'b110000111101001;
		Coeff[9085] <= 15'b110000111101011;
		Coeff[9086] <= 15'b110000111101101;
		Coeff[9087] <= 15'b110000111101111;
		Coeff[9088] <= 15'b110000111110001;
		Coeff[9089] <= 15'b110000111110011;
		Coeff[9090] <= 15'b110000111110101;
		Coeff[9091] <= 15'b110000111110111;
		Coeff[9092] <= 15'b110000111111001;
		Coeff[9093] <= 15'b110000111111011;
		Coeff[9094] <= 15'b110000111111101;
		Coeff[9095] <= 15'b110000111111111;
		Coeff[9096] <= 15'b110001000000001;
		Coeff[9097] <= 15'b110001000000011;
		Coeff[9098] <= 15'b110001000000101;
		Coeff[9099] <= 15'b110001000000111;
		Coeff[9100] <= 15'b110001000001001;
		Coeff[9101] <= 15'b110001000001011;
		Coeff[9102] <= 15'b110001000001101;
		Coeff[9103] <= 15'b110001000001111;
		Coeff[9104] <= 15'b110001000010001;
		Coeff[9105] <= 15'b110001000010011;
		Coeff[9106] <= 15'b110001000010101;
		Coeff[9107] <= 15'b110001000010111;
		Coeff[9108] <= 15'b110001000011001;
		Coeff[9109] <= 15'b110001000011011;
		Coeff[9110] <= 15'b110001000011101;
		Coeff[9111] <= 15'b110001000011111;
		Coeff[9112] <= 15'b110001000100001;
		Coeff[9113] <= 15'b110001000100011;
		Coeff[9114] <= 15'b110001000100110;
		Coeff[9115] <= 15'b110001000101000;
		Coeff[9116] <= 15'b110001000101010;
		Coeff[9117] <= 15'b110001000101100;
		Coeff[9118] <= 15'b110001000101110;
		Coeff[9119] <= 15'b110001000110000;
		Coeff[9120] <= 15'b110001000110010;
		Coeff[9121] <= 15'b110001000110100;
		Coeff[9122] <= 15'b110001000110110;
		Coeff[9123] <= 15'b110001000111000;
		Coeff[9124] <= 15'b110001000111010;
		Coeff[9125] <= 15'b110001000111100;
		Coeff[9126] <= 15'b110001000111110;
		Coeff[9127] <= 15'b110001001000000;
		Coeff[9128] <= 15'b110001001000010;
		Coeff[9129] <= 15'b110001001000100;
		Coeff[9130] <= 15'b110001001000110;
		Coeff[9131] <= 15'b110001001001000;
		Coeff[9132] <= 15'b110001001001010;
		Coeff[9133] <= 15'b110001001001100;
		Coeff[9134] <= 15'b110001001001110;
		Coeff[9135] <= 15'b110001001010000;
		Coeff[9136] <= 15'b110001001010010;
		Coeff[9137] <= 15'b110001001010100;
		Coeff[9138] <= 15'b110001001010110;
		Coeff[9139] <= 15'b110001001011000;
		Coeff[9140] <= 15'b110001001011010;
		Coeff[9141] <= 15'b110001001011100;
		Coeff[9142] <= 15'b110001001011110;
		Coeff[9143] <= 15'b110001001100000;
		Coeff[9144] <= 15'b110001001100010;
		Coeff[9145] <= 15'b110001001100100;
		Coeff[9146] <= 15'b110001001100110;
		Coeff[9147] <= 15'b110001001101000;
		Coeff[9148] <= 15'b110001001101010;
		Coeff[9149] <= 15'b110001001101100;
		Coeff[9150] <= 15'b110001001101110;
		Coeff[9151] <= 15'b110001001110000;
		Coeff[9152] <= 15'b110001001110010;
		Coeff[9153] <= 15'b110001001110100;
		Coeff[9154] <= 15'b110001001110110;
		Coeff[9155] <= 15'b110001001111000;
		Coeff[9156] <= 15'b110001001111010;
		Coeff[9157] <= 15'b110001001111100;
		Coeff[9158] <= 15'b110001001111110;
		Coeff[9159] <= 15'b110001010000000;
		Coeff[9160] <= 15'b110001010000010;
		Coeff[9161] <= 15'b110001010000100;
		Coeff[9162] <= 15'b110001010000110;
		Coeff[9163] <= 15'b110001010001000;
		Coeff[9164] <= 15'b110001010001010;
		Coeff[9165] <= 15'b110001010001100;
		Coeff[9166] <= 15'b110001010001110;
		Coeff[9167] <= 15'b110001010010000;
		Coeff[9168] <= 15'b110001010010010;
		Coeff[9169] <= 15'b110001010010100;
		Coeff[9170] <= 15'b110001010010110;
		Coeff[9171] <= 15'b110001010011000;
		Coeff[9172] <= 15'b110001010011010;
		Coeff[9173] <= 15'b110001010011100;
		Coeff[9174] <= 15'b110001010011110;
		Coeff[9175] <= 15'b110001010100000;
		Coeff[9176] <= 15'b110001010100010;
		Coeff[9177] <= 15'b110001010100100;
		Coeff[9178] <= 15'b110001010100110;
		Coeff[9179] <= 15'b110001010101000;
		Coeff[9180] <= 15'b110001010101010;
		Coeff[9181] <= 15'b110001010101100;
		Coeff[9182] <= 15'b110001010101110;
		Coeff[9183] <= 15'b110001010110000;
		Coeff[9184] <= 15'b110001010110010;
		Coeff[9185] <= 15'b110001010110100;
		Coeff[9186] <= 15'b110001010110110;
		Coeff[9187] <= 15'b110001010111000;
		Coeff[9188] <= 15'b110001010111010;
		Coeff[9189] <= 15'b110001010111100;
		Coeff[9190] <= 15'b110001010111110;
		Coeff[9191] <= 15'b110001011000000;
		Coeff[9192] <= 15'b110001011000010;
		Coeff[9193] <= 15'b110001011000100;
		Coeff[9194] <= 15'b110001011000110;
		Coeff[9195] <= 15'b110001011001000;
		Coeff[9196] <= 15'b110001011001010;
		Coeff[9197] <= 15'b110001011001100;
		Coeff[9198] <= 15'b110001011001110;
		Coeff[9199] <= 15'b110001011010000;
		Coeff[9200] <= 15'b110001011010010;
		Coeff[9201] <= 15'b110001011010100;
		Coeff[9202] <= 15'b110001011010110;
		Coeff[9203] <= 15'b110001011011000;
		Coeff[9204] <= 15'b110001011011010;
		Coeff[9205] <= 15'b110001011011100;
		Coeff[9206] <= 15'b110001011011110;
		Coeff[9207] <= 15'b110001011100000;
		Coeff[9208] <= 15'b110001011100010;
		Coeff[9209] <= 15'b110001011100100;
		Coeff[9210] <= 15'b110001011100110;
		Coeff[9211] <= 15'b110001011101000;
		Coeff[9212] <= 15'b110001011101010;
		Coeff[9213] <= 15'b110001011101100;
		Coeff[9214] <= 15'b110001011101110;
		Coeff[9215] <= 15'b110001011110000;
		Coeff[9216] <= 15'b110001011110010;
		Coeff[9217] <= 15'b110001011110100;
		Coeff[9218] <= 15'b110001011110110;
		Coeff[9219] <= 15'b110001011111000;
		Coeff[9220] <= 15'b110001011111010;
		Coeff[9221] <= 15'b110001011111100;
		Coeff[9222] <= 15'b110001011111110;
		Coeff[9223] <= 15'b110001100000000;
		Coeff[9224] <= 15'b110001100000010;
		Coeff[9225] <= 15'b110001100000100;
		Coeff[9226] <= 15'b110001100000110;
		Coeff[9227] <= 15'b110001100001000;
		Coeff[9228] <= 15'b110001100001010;
		Coeff[9229] <= 15'b110001100001100;
		Coeff[9230] <= 15'b110001100001110;
		Coeff[9231] <= 15'b110001100010000;
		Coeff[9232] <= 15'b110001100010010;
		Coeff[9233] <= 15'b110001100010100;
		Coeff[9234] <= 15'b110001100010110;
		Coeff[9235] <= 15'b110001100011000;
		Coeff[9236] <= 15'b110001100011010;
		Coeff[9237] <= 15'b110001100011100;
		Coeff[9238] <= 15'b110001100011110;
		Coeff[9239] <= 15'b110001100100000;
		Coeff[9240] <= 15'b110001100100010;
		Coeff[9241] <= 15'b110001100100100;
		Coeff[9242] <= 15'b110001100100110;
		Coeff[9243] <= 15'b110001100101000;
		Coeff[9244] <= 15'b110001100101010;
		Coeff[9245] <= 15'b110001100101100;
		Coeff[9246] <= 15'b110001100101110;
		Coeff[9247] <= 15'b110001100110000;
		Coeff[9248] <= 15'b110001100110010;
		Coeff[9249] <= 15'b110001100110100;
		Coeff[9250] <= 15'b110001100110110;
		Coeff[9251] <= 15'b110001100111000;
		Coeff[9252] <= 15'b110001100111010;
		Coeff[9253] <= 15'b110001100111100;
		Coeff[9254] <= 15'b110001100111110;
		Coeff[9255] <= 15'b110001101000000;
		Coeff[9256] <= 15'b110001101000010;
		Coeff[9257] <= 15'b110001101000100;
		Coeff[9258] <= 15'b110001101000110;
		Coeff[9259] <= 15'b110001101000111;
		Coeff[9260] <= 15'b110001101001001;
		Coeff[9261] <= 15'b110001101001011;
		Coeff[9262] <= 15'b110001101001101;
		Coeff[9263] <= 15'b110001101001111;
		Coeff[9264] <= 15'b110001101010001;
		Coeff[9265] <= 15'b110001101010011;
		Coeff[9266] <= 15'b110001101010101;
		Coeff[9267] <= 15'b110001101010111;
		Coeff[9268] <= 15'b110001101011001;
		Coeff[9269] <= 15'b110001101011011;
		Coeff[9270] <= 15'b110001101011101;
		Coeff[9271] <= 15'b110001101011111;
		Coeff[9272] <= 15'b110001101100001;
		Coeff[9273] <= 15'b110001101100011;
		Coeff[9274] <= 15'b110001101100101;
		Coeff[9275] <= 15'b110001101100111;
		Coeff[9276] <= 15'b110001101101001;
		Coeff[9277] <= 15'b110001101101011;
		Coeff[9278] <= 15'b110001101101101;
		Coeff[9279] <= 15'b110001101101111;
		Coeff[9280] <= 15'b110001101110001;
		Coeff[9281] <= 15'b110001101110011;
		Coeff[9282] <= 15'b110001101110101;
		Coeff[9283] <= 15'b110001101110111;
		Coeff[9284] <= 15'b110001101111001;
		Coeff[9285] <= 15'b110001101111011;
		Coeff[9286] <= 15'b110001101111101;
		Coeff[9287] <= 15'b110001101111111;
		Coeff[9288] <= 15'b110001110000001;
		Coeff[9289] <= 15'b110001110000011;
		Coeff[9290] <= 15'b110001110000101;
		Coeff[9291] <= 15'b110001110000111;
		Coeff[9292] <= 15'b110001110001001;
		Coeff[9293] <= 15'b110001110001011;
		Coeff[9294] <= 15'b110001110001101;
		Coeff[9295] <= 15'b110001110001111;
		Coeff[9296] <= 15'b110001110010001;
		Coeff[9297] <= 15'b110001110010011;
		Coeff[9298] <= 15'b110001110010101;
		Coeff[9299] <= 15'b110001110010111;
		Coeff[9300] <= 15'b110001110011001;
		Coeff[9301] <= 15'b110001110011011;
		Coeff[9302] <= 15'b110001110011101;
		Coeff[9303] <= 15'b110001110011111;
		Coeff[9304] <= 15'b110001110100000;
		Coeff[9305] <= 15'b110001110100010;
		Coeff[9306] <= 15'b110001110100100;
		Coeff[9307] <= 15'b110001110100110;
		Coeff[9308] <= 15'b110001110101000;
		Coeff[9309] <= 15'b110001110101010;
		Coeff[9310] <= 15'b110001110101100;
		Coeff[9311] <= 15'b110001110101110;
		Coeff[9312] <= 15'b110001110110000;
		Coeff[9313] <= 15'b110001110110010;
		Coeff[9314] <= 15'b110001110110100;
		Coeff[9315] <= 15'b110001110110110;
		Coeff[9316] <= 15'b110001110111000;
		Coeff[9317] <= 15'b110001110111010;
		Coeff[9318] <= 15'b110001110111100;
		Coeff[9319] <= 15'b110001110111110;
		Coeff[9320] <= 15'b110001111000000;
		Coeff[9321] <= 15'b110001111000010;
		Coeff[9322] <= 15'b110001111000100;
		Coeff[9323] <= 15'b110001111000110;
		Coeff[9324] <= 15'b110001111001000;
		Coeff[9325] <= 15'b110001111001010;
		Coeff[9326] <= 15'b110001111001100;
		Coeff[9327] <= 15'b110001111001110;
		Coeff[9328] <= 15'b110001111010000;
		Coeff[9329] <= 15'b110001111010010;
		Coeff[9330] <= 15'b110001111010100;
		Coeff[9331] <= 15'b110001111010110;
		Coeff[9332] <= 15'b110001111011000;
		Coeff[9333] <= 15'b110001111011010;
		Coeff[9334] <= 15'b110001111011100;
		Coeff[9335] <= 15'b110001111011110;
		Coeff[9336] <= 15'b110001111011111;
		Coeff[9337] <= 15'b110001111100001;
		Coeff[9338] <= 15'b110001111100011;
		Coeff[9339] <= 15'b110001111100101;
		Coeff[9340] <= 15'b110001111100111;
		Coeff[9341] <= 15'b110001111101001;
		Coeff[9342] <= 15'b110001111101011;
		Coeff[9343] <= 15'b110001111101101;
		Coeff[9344] <= 15'b110001111101111;
		Coeff[9345] <= 15'b110001111110001;
		Coeff[9346] <= 15'b110001111110011;
		Coeff[9347] <= 15'b110001111110101;
		Coeff[9348] <= 15'b110001111110111;
		Coeff[9349] <= 15'b110001111111001;
		Coeff[9350] <= 15'b110001111111011;
		Coeff[9351] <= 15'b110001111111101;
		Coeff[9352] <= 15'b110001111111111;
		Coeff[9353] <= 15'b110010000000001;
		Coeff[9354] <= 15'b110010000000011;
		Coeff[9355] <= 15'b110010000000101;
		Coeff[9356] <= 15'b110010000000111;
		Coeff[9357] <= 15'b110010000001001;
		Coeff[9358] <= 15'b110010000001011;
		Coeff[9359] <= 15'b110010000001101;
		Coeff[9360] <= 15'b110010000001111;
		Coeff[9361] <= 15'b110010000010001;
		Coeff[9362] <= 15'b110010000010010;
		Coeff[9363] <= 15'b110010000010100;
		Coeff[9364] <= 15'b110010000010110;
		Coeff[9365] <= 15'b110010000011000;
		Coeff[9366] <= 15'b110010000011010;
		Coeff[9367] <= 15'b110010000011100;
		Coeff[9368] <= 15'b110010000011110;
		Coeff[9369] <= 15'b110010000100000;
		Coeff[9370] <= 15'b110010000100010;
		Coeff[9371] <= 15'b110010000100100;
		Coeff[9372] <= 15'b110010000100110;
		Coeff[9373] <= 15'b110010000101000;
		Coeff[9374] <= 15'b110010000101010;
		Coeff[9375] <= 15'b110010000101100;
		Coeff[9376] <= 15'b110010000101110;
		Coeff[9377] <= 15'b110010000110000;
		Coeff[9378] <= 15'b110010000110010;
		Coeff[9379] <= 15'b110010000110100;
		Coeff[9380] <= 15'b110010000110110;
		Coeff[9381] <= 15'b110010000111000;
		Coeff[9382] <= 15'b110010000111010;
		Coeff[9383] <= 15'b110010000111100;
		Coeff[9384] <= 15'b110010000111110;
		Coeff[9385] <= 15'b110010000111111;
		Coeff[9386] <= 15'b110010001000001;
		Coeff[9387] <= 15'b110010001000011;
		Coeff[9388] <= 15'b110010001000101;
		Coeff[9389] <= 15'b110010001000111;
		Coeff[9390] <= 15'b110010001001001;
		Coeff[9391] <= 15'b110010001001011;
		Coeff[9392] <= 15'b110010001001101;
		Coeff[9393] <= 15'b110010001001111;
		Coeff[9394] <= 15'b110010001010001;
		Coeff[9395] <= 15'b110010001010011;
		Coeff[9396] <= 15'b110010001010101;
		Coeff[9397] <= 15'b110010001010111;
		Coeff[9398] <= 15'b110010001011001;
		Coeff[9399] <= 15'b110010001011011;
		Coeff[9400] <= 15'b110010001011101;
		Coeff[9401] <= 15'b110010001011111;
		Coeff[9402] <= 15'b110010001100001;
		Coeff[9403] <= 15'b110010001100011;
		Coeff[9404] <= 15'b110010001100101;
		Coeff[9405] <= 15'b110010001100111;
		Coeff[9406] <= 15'b110010001101000;
		Coeff[9407] <= 15'b110010001101010;
		Coeff[9408] <= 15'b110010001101100;
		Coeff[9409] <= 15'b110010001101110;
		Coeff[9410] <= 15'b110010001110000;
		Coeff[9411] <= 15'b110010001110010;
		Coeff[9412] <= 15'b110010001110100;
		Coeff[9413] <= 15'b110010001110110;
		Coeff[9414] <= 15'b110010001111000;
		Coeff[9415] <= 15'b110010001111010;
		Coeff[9416] <= 15'b110010001111100;
		Coeff[9417] <= 15'b110010001111110;
		Coeff[9418] <= 15'b110010010000000;
		Coeff[9419] <= 15'b110010010000010;
		Coeff[9420] <= 15'b110010010000100;
		Coeff[9421] <= 15'b110010010000110;
		Coeff[9422] <= 15'b110010010001000;
		Coeff[9423] <= 15'b110010010001010;
		Coeff[9424] <= 15'b110010010001011;
		Coeff[9425] <= 15'b110010010001101;
		Coeff[9426] <= 15'b110010010001111;
		Coeff[9427] <= 15'b110010010010001;
		Coeff[9428] <= 15'b110010010010011;
		Coeff[9429] <= 15'b110010010010101;
		Coeff[9430] <= 15'b110010010010111;
		Coeff[9431] <= 15'b110010010011001;
		Coeff[9432] <= 15'b110010010011011;
		Coeff[9433] <= 15'b110010010011101;
		Coeff[9434] <= 15'b110010010011111;
		Coeff[9435] <= 15'b110010010100001;
		Coeff[9436] <= 15'b110010010100011;
		Coeff[9437] <= 15'b110010010100101;
		Coeff[9438] <= 15'b110010010100111;
		Coeff[9439] <= 15'b110010010101001;
		Coeff[9440] <= 15'b110010010101011;
		Coeff[9441] <= 15'b110010010101101;
		Coeff[9442] <= 15'b110010010101110;
		Coeff[9443] <= 15'b110010010110000;
		Coeff[9444] <= 15'b110010010110010;
		Coeff[9445] <= 15'b110010010110100;
		Coeff[9446] <= 15'b110010010110110;
		Coeff[9447] <= 15'b110010010111000;
		Coeff[9448] <= 15'b110010010111010;
		Coeff[9449] <= 15'b110010010111100;
		Coeff[9450] <= 15'b110010010111110;
		Coeff[9451] <= 15'b110010011000000;
		Coeff[9452] <= 15'b110010011000010;
		Coeff[9453] <= 15'b110010011000100;
		Coeff[9454] <= 15'b110010011000110;
		Coeff[9455] <= 15'b110010011001000;
		Coeff[9456] <= 15'b110010011001010;
		Coeff[9457] <= 15'b110010011001100;
		Coeff[9458] <= 15'b110010011001101;
		Coeff[9459] <= 15'b110010011001111;
		Coeff[9460] <= 15'b110010011010001;
		Coeff[9461] <= 15'b110010011010011;
		Coeff[9462] <= 15'b110010011010101;
		Coeff[9463] <= 15'b110010011010111;
		Coeff[9464] <= 15'b110010011011001;
		Coeff[9465] <= 15'b110010011011011;
		Coeff[9466] <= 15'b110010011011101;
		Coeff[9467] <= 15'b110010011011111;
		Coeff[9468] <= 15'b110010011100001;
		Coeff[9469] <= 15'b110010011100011;
		Coeff[9470] <= 15'b110010011100101;
		Coeff[9471] <= 15'b110010011100111;
		Coeff[9472] <= 15'b110010011101001;
		Coeff[9473] <= 15'b110010011101010;
		Coeff[9474] <= 15'b110010011101100;
		Coeff[9475] <= 15'b110010011101110;
		Coeff[9476] <= 15'b110010011110000;
		Coeff[9477] <= 15'b110010011110010;
		Coeff[9478] <= 15'b110010011110100;
		Coeff[9479] <= 15'b110010011110110;
		Coeff[9480] <= 15'b110010011111000;
		Coeff[9481] <= 15'b110010011111010;
		Coeff[9482] <= 15'b110010011111100;
		Coeff[9483] <= 15'b110010011111110;
		Coeff[9484] <= 15'b110010100000000;
		Coeff[9485] <= 15'b110010100000010;
		Coeff[9486] <= 15'b110010100000100;
		Coeff[9487] <= 15'b110010100000110;
		Coeff[9488] <= 15'b110010100000111;
		Coeff[9489] <= 15'b110010100001001;
		Coeff[9490] <= 15'b110010100001011;
		Coeff[9491] <= 15'b110010100001101;
		Coeff[9492] <= 15'b110010100001111;
		Coeff[9493] <= 15'b110010100010001;
		Coeff[9494] <= 15'b110010100010011;
		Coeff[9495] <= 15'b110010100010101;
		Coeff[9496] <= 15'b110010100010111;
		Coeff[9497] <= 15'b110010100011001;
		Coeff[9498] <= 15'b110010100011011;
		Coeff[9499] <= 15'b110010100011101;
		Coeff[9500] <= 15'b110010100011111;
		Coeff[9501] <= 15'b110010100100000;
		Coeff[9502] <= 15'b110010100100010;
		Coeff[9503] <= 15'b110010100100100;
		Coeff[9504] <= 15'b110010100100110;
		Coeff[9505] <= 15'b110010100101000;
		Coeff[9506] <= 15'b110010100101010;
		Coeff[9507] <= 15'b110010100101100;
		Coeff[9508] <= 15'b110010100101110;
		Coeff[9509] <= 15'b110010100110000;
		Coeff[9510] <= 15'b110010100110010;
		Coeff[9511] <= 15'b110010100110100;
		Coeff[9512] <= 15'b110010100110110;
		Coeff[9513] <= 15'b110010100111000;
		Coeff[9514] <= 15'b110010100111010;
		Coeff[9515] <= 15'b110010100111011;
		Coeff[9516] <= 15'b110010100111101;
		Coeff[9517] <= 15'b110010100111111;
		Coeff[9518] <= 15'b110010101000001;
		Coeff[9519] <= 15'b110010101000011;
		Coeff[9520] <= 15'b110010101000101;
		Coeff[9521] <= 15'b110010101000111;
		Coeff[9522] <= 15'b110010101001001;
		Coeff[9523] <= 15'b110010101001011;
		Coeff[9524] <= 15'b110010101001101;
		Coeff[9525] <= 15'b110010101001111;
		Coeff[9526] <= 15'b110010101010001;
		Coeff[9527] <= 15'b110010101010010;
		Coeff[9528] <= 15'b110010101010100;
		Coeff[9529] <= 15'b110010101010110;
		Coeff[9530] <= 15'b110010101011000;
		Coeff[9531] <= 15'b110010101011010;
		Coeff[9532] <= 15'b110010101011100;
		Coeff[9533] <= 15'b110010101011110;
		Coeff[9534] <= 15'b110010101100000;
		Coeff[9535] <= 15'b110010101100010;
		Coeff[9536] <= 15'b110010101100100;
		Coeff[9537] <= 15'b110010101100110;
		Coeff[9538] <= 15'b110010101101000;
		Coeff[9539] <= 15'b110010101101001;
		Coeff[9540] <= 15'b110010101101011;
		Coeff[9541] <= 15'b110010101101101;
		Coeff[9542] <= 15'b110010101101111;
		Coeff[9543] <= 15'b110010101110001;
		Coeff[9544] <= 15'b110010101110011;
		Coeff[9545] <= 15'b110010101110101;
		Coeff[9546] <= 15'b110010101110111;
		Coeff[9547] <= 15'b110010101111001;
		Coeff[9548] <= 15'b110010101111011;
		Coeff[9549] <= 15'b110010101111101;
		Coeff[9550] <= 15'b110010101111111;
		Coeff[9551] <= 15'b110010110000000;
		Coeff[9552] <= 15'b110010110000010;
		Coeff[9553] <= 15'b110010110000100;
		Coeff[9554] <= 15'b110010110000110;
		Coeff[9555] <= 15'b110010110001000;
		Coeff[9556] <= 15'b110010110001010;
		Coeff[9557] <= 15'b110010110001100;
		Coeff[9558] <= 15'b110010110001110;
		Coeff[9559] <= 15'b110010110010000;
		Coeff[9560] <= 15'b110010110010010;
		Coeff[9561] <= 15'b110010110010100;
		Coeff[9562] <= 15'b110010110010110;
		Coeff[9563] <= 15'b110010110010111;
		Coeff[9564] <= 15'b110010110011001;
		Coeff[9565] <= 15'b110010110011011;
		Coeff[9566] <= 15'b110010110011101;
		Coeff[9567] <= 15'b110010110011111;
		Coeff[9568] <= 15'b110010110100001;
		Coeff[9569] <= 15'b110010110100011;
		Coeff[9570] <= 15'b110010110100101;
		Coeff[9571] <= 15'b110010110100111;
		Coeff[9572] <= 15'b110010110101001;
		Coeff[9573] <= 15'b110010110101011;
		Coeff[9574] <= 15'b110010110101100;
		Coeff[9575] <= 15'b110010110101110;
		Coeff[9576] <= 15'b110010110110000;
		Coeff[9577] <= 15'b110010110110010;
		Coeff[9578] <= 15'b110010110110100;
		Coeff[9579] <= 15'b110010110110110;
		Coeff[9580] <= 15'b110010110111000;
		Coeff[9581] <= 15'b110010110111010;
		Coeff[9582] <= 15'b110010110111100;
		Coeff[9583] <= 15'b110010110111110;
		Coeff[9584] <= 15'b110010111000000;
		Coeff[9585] <= 15'b110010111000001;
		Coeff[9586] <= 15'b110010111000011;
		Coeff[9587] <= 15'b110010111000101;
		Coeff[9588] <= 15'b110010111000111;
		Coeff[9589] <= 15'b110010111001001;
		Coeff[9590] <= 15'b110010111001011;
		Coeff[9591] <= 15'b110010111001101;
		Coeff[9592] <= 15'b110010111001111;
		Coeff[9593] <= 15'b110010111010001;
		Coeff[9594] <= 15'b110010111010011;
		Coeff[9595] <= 15'b110010111010100;
		Coeff[9596] <= 15'b110010111010110;
		Coeff[9597] <= 15'b110010111011000;
		Coeff[9598] <= 15'b110010111011010;
		Coeff[9599] <= 15'b110010111011100;
		Coeff[9600] <= 15'b110010111011110;
		Coeff[9601] <= 15'b110010111100000;
		Coeff[9602] <= 15'b110010111100010;
		Coeff[9603] <= 15'b110010111100100;
		Coeff[9604] <= 15'b110010111100110;
		Coeff[9605] <= 15'b110010111100111;
		Coeff[9606] <= 15'b110010111101001;
		Coeff[9607] <= 15'b110010111101011;
		Coeff[9608] <= 15'b110010111101101;
		Coeff[9609] <= 15'b110010111101111;
		Coeff[9610] <= 15'b110010111110001;
		Coeff[9611] <= 15'b110010111110011;
		Coeff[9612] <= 15'b110010111110101;
		Coeff[9613] <= 15'b110010111110111;
		Coeff[9614] <= 15'b110010111111001;
		Coeff[9615] <= 15'b110010111111010;
		Coeff[9616] <= 15'b110010111111100;
		Coeff[9617] <= 15'b110010111111110;
		Coeff[9618] <= 15'b110011000000000;
		Coeff[9619] <= 15'b110011000000010;
		Coeff[9620] <= 15'b110011000000100;
		Coeff[9621] <= 15'b110011000000110;
		Coeff[9622] <= 15'b110011000001000;
		Coeff[9623] <= 15'b110011000001010;
		Coeff[9624] <= 15'b110011000001100;
		Coeff[9625] <= 15'b110011000001101;
		Coeff[9626] <= 15'b110011000001111;
		Coeff[9627] <= 15'b110011000010001;
		Coeff[9628] <= 15'b110011000010011;
		Coeff[9629] <= 15'b110011000010101;
		Coeff[9630] <= 15'b110011000010111;
		Coeff[9631] <= 15'b110011000011001;
		Coeff[9632] <= 15'b110011000011011;
		Coeff[9633] <= 15'b110011000011101;
		Coeff[9634] <= 15'b110011000011111;
		Coeff[9635] <= 15'b110011000100000;
		Coeff[9636] <= 15'b110011000100010;
		Coeff[9637] <= 15'b110011000100100;
		Coeff[9638] <= 15'b110011000100110;
		Coeff[9639] <= 15'b110011000101000;
		Coeff[9640] <= 15'b110011000101010;
		Coeff[9641] <= 15'b110011000101100;
		Coeff[9642] <= 15'b110011000101110;
		Coeff[9643] <= 15'b110011000110000;
		Coeff[9644] <= 15'b110011000110001;
		Coeff[9645] <= 15'b110011000110011;
		Coeff[9646] <= 15'b110011000110101;
		Coeff[9647] <= 15'b110011000110111;
		Coeff[9648] <= 15'b110011000111001;
		Coeff[9649] <= 15'b110011000111011;
		Coeff[9650] <= 15'b110011000111101;
		Coeff[9651] <= 15'b110011000111111;
		Coeff[9652] <= 15'b110011001000001;
		Coeff[9653] <= 15'b110011001000010;
		Coeff[9654] <= 15'b110011001000100;
		Coeff[9655] <= 15'b110011001000110;
		Coeff[9656] <= 15'b110011001001000;
		Coeff[9657] <= 15'b110011001001010;
		Coeff[9658] <= 15'b110011001001100;
		Coeff[9659] <= 15'b110011001001110;
		Coeff[9660] <= 15'b110011001010000;
		Coeff[9661] <= 15'b110011001010010;
		Coeff[9662] <= 15'b110011001010011;
		Coeff[9663] <= 15'b110011001010101;
		Coeff[9664] <= 15'b110011001010111;
		Coeff[9665] <= 15'b110011001011001;
		Coeff[9666] <= 15'b110011001011011;
		Coeff[9667] <= 15'b110011001011101;
		Coeff[9668] <= 15'b110011001011111;
		Coeff[9669] <= 15'b110011001100001;
		Coeff[9670] <= 15'b110011001100011;
		Coeff[9671] <= 15'b110011001100100;
		Coeff[9672] <= 15'b110011001100110;
		Coeff[9673] <= 15'b110011001101000;
		Coeff[9674] <= 15'b110011001101010;
		Coeff[9675] <= 15'b110011001101100;
		Coeff[9676] <= 15'b110011001101110;
		Coeff[9677] <= 15'b110011001110000;
		Coeff[9678] <= 15'b110011001110010;
		Coeff[9679] <= 15'b110011001110100;
		Coeff[9680] <= 15'b110011001110101;
		Coeff[9681] <= 15'b110011001110111;
		Coeff[9682] <= 15'b110011001111001;
		Coeff[9683] <= 15'b110011001111011;
		Coeff[9684] <= 15'b110011001111101;
		Coeff[9685] <= 15'b110011001111111;
		Coeff[9686] <= 15'b110011010000001;
		Coeff[9687] <= 15'b110011010000011;
		Coeff[9688] <= 15'b110011010000100;
		Coeff[9689] <= 15'b110011010000110;
		Coeff[9690] <= 15'b110011010001000;
		Coeff[9691] <= 15'b110011010001010;
		Coeff[9692] <= 15'b110011010001100;
		Coeff[9693] <= 15'b110011010001110;
		Coeff[9694] <= 15'b110011010010000;
		Coeff[9695] <= 15'b110011010010010;
		Coeff[9696] <= 15'b110011010010011;
		Coeff[9697] <= 15'b110011010010101;
		Coeff[9698] <= 15'b110011010010111;
		Coeff[9699] <= 15'b110011010011001;
		Coeff[9700] <= 15'b110011010011011;
		Coeff[9701] <= 15'b110011010011101;
		Coeff[9702] <= 15'b110011010011111;
		Coeff[9703] <= 15'b110011010100001;
		Coeff[9704] <= 15'b110011010100011;
		Coeff[9705] <= 15'b110011010100100;
		Coeff[9706] <= 15'b110011010100110;
		Coeff[9707] <= 15'b110011010101000;
		Coeff[9708] <= 15'b110011010101010;
		Coeff[9709] <= 15'b110011010101100;
		Coeff[9710] <= 15'b110011010101110;
		Coeff[9711] <= 15'b110011010110000;
		Coeff[9712] <= 15'b110011010110010;
		Coeff[9713] <= 15'b110011010110011;
		Coeff[9714] <= 15'b110011010110101;
		Coeff[9715] <= 15'b110011010110111;
		Coeff[9716] <= 15'b110011010111001;
		Coeff[9717] <= 15'b110011010111011;
		Coeff[9718] <= 15'b110011010111101;
		Coeff[9719] <= 15'b110011010111111;
		Coeff[9720] <= 15'b110011011000001;
		Coeff[9721] <= 15'b110011011000010;
		Coeff[9722] <= 15'b110011011000100;
		Coeff[9723] <= 15'b110011011000110;
		Coeff[9724] <= 15'b110011011001000;
		Coeff[9725] <= 15'b110011011001010;
		Coeff[9726] <= 15'b110011011001100;
		Coeff[9727] <= 15'b110011011001110;
		Coeff[9728] <= 15'b110011011010000;
		Coeff[9729] <= 15'b110011011010001;
		Coeff[9730] <= 15'b110011011010011;
		Coeff[9731] <= 15'b110011011010101;
		Coeff[9732] <= 15'b110011011010111;
		Coeff[9733] <= 15'b110011011011001;
		Coeff[9734] <= 15'b110011011011011;
		Coeff[9735] <= 15'b110011011011101;
		Coeff[9736] <= 15'b110011011011110;
		Coeff[9737] <= 15'b110011011100000;
		Coeff[9738] <= 15'b110011011100010;
		Coeff[9739] <= 15'b110011011100100;
		Coeff[9740] <= 15'b110011011100110;
		Coeff[9741] <= 15'b110011011101000;
		Coeff[9742] <= 15'b110011011101010;
		Coeff[9743] <= 15'b110011011101100;
		Coeff[9744] <= 15'b110011011101101;
		Coeff[9745] <= 15'b110011011101111;
		Coeff[9746] <= 15'b110011011110001;
		Coeff[9747] <= 15'b110011011110011;
		Coeff[9748] <= 15'b110011011110101;
		Coeff[9749] <= 15'b110011011110111;
		Coeff[9750] <= 15'b110011011111001;
		Coeff[9751] <= 15'b110011011111010;
		Coeff[9752] <= 15'b110011011111100;
		Coeff[9753] <= 15'b110011011111110;
		Coeff[9754] <= 15'b110011100000000;
		Coeff[9755] <= 15'b110011100000010;
		Coeff[9756] <= 15'b110011100000100;
		Coeff[9757] <= 15'b110011100000110;
		Coeff[9758] <= 15'b110011100001000;
		Coeff[9759] <= 15'b110011100001001;
		Coeff[9760] <= 15'b110011100001011;
		Coeff[9761] <= 15'b110011100001101;
		Coeff[9762] <= 15'b110011100001111;
		Coeff[9763] <= 15'b110011100010001;
		Coeff[9764] <= 15'b110011100010011;
		Coeff[9765] <= 15'b110011100010101;
		Coeff[9766] <= 15'b110011100010110;
		Coeff[9767] <= 15'b110011100011000;
		Coeff[9768] <= 15'b110011100011010;
		Coeff[9769] <= 15'b110011100011100;
		Coeff[9770] <= 15'b110011100011110;
		Coeff[9771] <= 15'b110011100100000;
		Coeff[9772] <= 15'b110011100100010;
		Coeff[9773] <= 15'b110011100100011;
		Coeff[9774] <= 15'b110011100100101;
		Coeff[9775] <= 15'b110011100100111;
		Coeff[9776] <= 15'b110011100101001;
		Coeff[9777] <= 15'b110011100101011;
		Coeff[9778] <= 15'b110011100101101;
		Coeff[9779] <= 15'b110011100101111;
		Coeff[9780] <= 15'b110011100110000;
		Coeff[9781] <= 15'b110011100110010;
		Coeff[9782] <= 15'b110011100110100;
		Coeff[9783] <= 15'b110011100110110;
		Coeff[9784] <= 15'b110011100111000;
		Coeff[9785] <= 15'b110011100111010;
		Coeff[9786] <= 15'b110011100111100;
		Coeff[9787] <= 15'b110011100111101;
		Coeff[9788] <= 15'b110011100111111;
		Coeff[9789] <= 15'b110011101000001;
		Coeff[9790] <= 15'b110011101000011;
		Coeff[9791] <= 15'b110011101000101;
		Coeff[9792] <= 15'b110011101000111;
		Coeff[9793] <= 15'b110011101001001;
		Coeff[9794] <= 15'b110011101001010;
		Coeff[9795] <= 15'b110011101001100;
		Coeff[9796] <= 15'b110011101001110;
		Coeff[9797] <= 15'b110011101010000;
		Coeff[9798] <= 15'b110011101010010;
		Coeff[9799] <= 15'b110011101010100;
		Coeff[9800] <= 15'b110011101010110;
		Coeff[9801] <= 15'b110011101010111;
		Coeff[9802] <= 15'b110011101011001;
		Coeff[9803] <= 15'b110011101011011;
		Coeff[9804] <= 15'b110011101011101;
		Coeff[9805] <= 15'b110011101011111;
		Coeff[9806] <= 15'b110011101100001;
		Coeff[9807] <= 15'b110011101100011;
		Coeff[9808] <= 15'b110011101100100;
		Coeff[9809] <= 15'b110011101100110;
		Coeff[9810] <= 15'b110011101101000;
		Coeff[9811] <= 15'b110011101101010;
		Coeff[9812] <= 15'b110011101101100;
		Coeff[9813] <= 15'b110011101101110;
		Coeff[9814] <= 15'b110011101110000;
		Coeff[9815] <= 15'b110011101110001;
		Coeff[9816] <= 15'b110011101110011;
		Coeff[9817] <= 15'b110011101110101;
		Coeff[9818] <= 15'b110011101110111;
		Coeff[9819] <= 15'b110011101111001;
		Coeff[9820] <= 15'b110011101111011;
		Coeff[9821] <= 15'b110011101111101;
		Coeff[9822] <= 15'b110011101111110;
		Coeff[9823] <= 15'b110011110000000;
		Coeff[9824] <= 15'b110011110000010;
		Coeff[9825] <= 15'b110011110000100;
		Coeff[9826] <= 15'b110011110000110;
		Coeff[9827] <= 15'b110011110001000;
		Coeff[9828] <= 15'b110011110001001;
		Coeff[9829] <= 15'b110011110001011;
		Coeff[9830] <= 15'b110011110001101;
		Coeff[9831] <= 15'b110011110001111;
		Coeff[9832] <= 15'b110011110010001;
		Coeff[9833] <= 15'b110011110010011;
		Coeff[9834] <= 15'b110011110010101;
		Coeff[9835] <= 15'b110011110010110;
		Coeff[9836] <= 15'b110011110011000;
		Coeff[9837] <= 15'b110011110011010;
		Coeff[9838] <= 15'b110011110011100;
		Coeff[9839] <= 15'b110011110011110;
		Coeff[9840] <= 15'b110011110100000;
		Coeff[9841] <= 15'b110011110100001;
		Coeff[9842] <= 15'b110011110100011;
		Coeff[9843] <= 15'b110011110100101;
		Coeff[9844] <= 15'b110011110100111;
		Coeff[9845] <= 15'b110011110101001;
		Coeff[9846] <= 15'b110011110101011;
		Coeff[9847] <= 15'b110011110101100;
		Coeff[9848] <= 15'b110011110101110;
		Coeff[9849] <= 15'b110011110110000;
		Coeff[9850] <= 15'b110011110110010;
		Coeff[9851] <= 15'b110011110110100;
		Coeff[9852] <= 15'b110011110110110;
		Coeff[9853] <= 15'b110011110111000;
		Coeff[9854] <= 15'b110011110111001;
		Coeff[9855] <= 15'b110011110111011;
		Coeff[9856] <= 15'b110011110111101;
		Coeff[9857] <= 15'b110011110111111;
		Coeff[9858] <= 15'b110011111000001;
		Coeff[9859] <= 15'b110011111000011;
		Coeff[9860] <= 15'b110011111000100;
		Coeff[9861] <= 15'b110011111000110;
		Coeff[9862] <= 15'b110011111001000;
		Coeff[9863] <= 15'b110011111001010;
		Coeff[9864] <= 15'b110011111001100;
		Coeff[9865] <= 15'b110011111001110;
		Coeff[9866] <= 15'b110011111001111;
		Coeff[9867] <= 15'b110011111010001;
		Coeff[9868] <= 15'b110011111010011;
		Coeff[9869] <= 15'b110011111010101;
		Coeff[9870] <= 15'b110011111010111;
		Coeff[9871] <= 15'b110011111011001;
		Coeff[9872] <= 15'b110011111011010;
		Coeff[9873] <= 15'b110011111011100;
		Coeff[9874] <= 15'b110011111011110;
		Coeff[9875] <= 15'b110011111100000;
		Coeff[9876] <= 15'b110011111100010;
		Coeff[9877] <= 15'b110011111100100;
		Coeff[9878] <= 15'b110011111100101;
		Coeff[9879] <= 15'b110011111100111;
		Coeff[9880] <= 15'b110011111101001;
		Coeff[9881] <= 15'b110011111101011;
		Coeff[9882] <= 15'b110011111101101;
		Coeff[9883] <= 15'b110011111101111;
		Coeff[9884] <= 15'b110011111110000;
		Coeff[9885] <= 15'b110011111110010;
		Coeff[9886] <= 15'b110011111110100;
		Coeff[9887] <= 15'b110011111110110;
		Coeff[9888] <= 15'b110011111111000;
		Coeff[9889] <= 15'b110011111111010;
		Coeff[9890] <= 15'b110011111111011;
		Coeff[9891] <= 15'b110011111111101;
		Coeff[9892] <= 15'b110011111111111;
		Coeff[9893] <= 15'b110100000000001;
		Coeff[9894] <= 15'b110100000000011;
		Coeff[9895] <= 15'b110100000000101;
		Coeff[9896] <= 15'b110100000000110;
		Coeff[9897] <= 15'b110100000001000;
		Coeff[9898] <= 15'b110100000001010;
		Coeff[9899] <= 15'b110100000001100;
		Coeff[9900] <= 15'b110100000001110;
		Coeff[9901] <= 15'b110100000010000;
		Coeff[9902] <= 15'b110100000010001;
		Coeff[9903] <= 15'b110100000010011;
		Coeff[9904] <= 15'b110100000010101;
		Coeff[9905] <= 15'b110100000010111;
		Coeff[9906] <= 15'b110100000011001;
		Coeff[9907] <= 15'b110100000011011;
		Coeff[9908] <= 15'b110100000011100;
		Coeff[9909] <= 15'b110100000011110;
		Coeff[9910] <= 15'b110100000100000;
		Coeff[9911] <= 15'b110100000100010;
		Coeff[9912] <= 15'b110100000100100;
		Coeff[9913] <= 15'b110100000100110;
		Coeff[9914] <= 15'b110100000100111;
		Coeff[9915] <= 15'b110100000101001;
		Coeff[9916] <= 15'b110100000101011;
		Coeff[9917] <= 15'b110100000101101;
		Coeff[9918] <= 15'b110100000101111;
		Coeff[9919] <= 15'b110100000110001;
		Coeff[9920] <= 15'b110100000110010;
		Coeff[9921] <= 15'b110100000110100;
		Coeff[9922] <= 15'b110100000110110;
		Coeff[9923] <= 15'b110100000111000;
		Coeff[9924] <= 15'b110100000111010;
		Coeff[9925] <= 15'b110100000111011;
		Coeff[9926] <= 15'b110100000111101;
		Coeff[9927] <= 15'b110100000111111;
		Coeff[9928] <= 15'b110100001000001;
		Coeff[9929] <= 15'b110100001000011;
		Coeff[9930] <= 15'b110100001000101;
		Coeff[9931] <= 15'b110100001000110;
		Coeff[9932] <= 15'b110100001001000;
		Coeff[9933] <= 15'b110100001001010;
		Coeff[9934] <= 15'b110100001001100;
		Coeff[9935] <= 15'b110100001001110;
		Coeff[9936] <= 15'b110100001010000;
		Coeff[9937] <= 15'b110100001010001;
		Coeff[9938] <= 15'b110100001010011;
		Coeff[9939] <= 15'b110100001010101;
		Coeff[9940] <= 15'b110100001010111;
		Coeff[9941] <= 15'b110100001011001;
		Coeff[9942] <= 15'b110100001011010;
		Coeff[9943] <= 15'b110100001011100;
		Coeff[9944] <= 15'b110100001011110;
		Coeff[9945] <= 15'b110100001100000;
		Coeff[9946] <= 15'b110100001100010;
		Coeff[9947] <= 15'b110100001100100;
		Coeff[9948] <= 15'b110100001100101;
		Coeff[9949] <= 15'b110100001100111;
		Coeff[9950] <= 15'b110100001101001;
		Coeff[9951] <= 15'b110100001101011;
		Coeff[9952] <= 15'b110100001101101;
		Coeff[9953] <= 15'b110100001101110;
		Coeff[9954] <= 15'b110100001110000;
		Coeff[9955] <= 15'b110100001110010;
		Coeff[9956] <= 15'b110100001110100;
		Coeff[9957] <= 15'b110100001110110;
		Coeff[9958] <= 15'b110100001111000;
		Coeff[9959] <= 15'b110100001111001;
		Coeff[9960] <= 15'b110100001111011;
		Coeff[9961] <= 15'b110100001111101;
		Coeff[9962] <= 15'b110100001111111;
		Coeff[9963] <= 15'b110100010000001;
		Coeff[9964] <= 15'b110100010000010;
		Coeff[9965] <= 15'b110100010000100;
		Coeff[9966] <= 15'b110100010000110;
		Coeff[9967] <= 15'b110100010001000;
		Coeff[9968] <= 15'b110100010001010;
		Coeff[9969] <= 15'b110100010001011;
		Coeff[9970] <= 15'b110100010001101;
		Coeff[9971] <= 15'b110100010001111;
		Coeff[9972] <= 15'b110100010010001;
		Coeff[9973] <= 15'b110100010010011;
		Coeff[9974] <= 15'b110100010010101;
		Coeff[9975] <= 15'b110100010010110;
		Coeff[9976] <= 15'b110100010011000;
		Coeff[9977] <= 15'b110100010011010;
		Coeff[9978] <= 15'b110100010011100;
		Coeff[9979] <= 15'b110100010011110;
		Coeff[9980] <= 15'b110100010011111;
		Coeff[9981] <= 15'b110100010100001;
		Coeff[9982] <= 15'b110100010100011;
		Coeff[9983] <= 15'b110100010100101;
		Coeff[9984] <= 15'b110100010100111;
		Coeff[9985] <= 15'b110100010101000;
		Coeff[9986] <= 15'b110100010101010;
		Coeff[9987] <= 15'b110100010101100;
		Coeff[9988] <= 15'b110100010101110;
		Coeff[9989] <= 15'b110100010110000;
		Coeff[9990] <= 15'b110100010110001;
		Coeff[9991] <= 15'b110100010110011;
		Coeff[9992] <= 15'b110100010110101;
		Coeff[9993] <= 15'b110100010110111;
		Coeff[9994] <= 15'b110100010111001;
		Coeff[9995] <= 15'b110100010111011;
		Coeff[9996] <= 15'b110100010111100;
		Coeff[9997] <= 15'b110100010111110;
		Coeff[9998] <= 15'b110100011000000;
		Coeff[9999] <= 15'b110100011000010;
		Coeff[10000] <= 15'b110100011000100;
		Coeff[10001] <= 15'b110100011000101;
		Coeff[10002] <= 15'b110100011000111;
		Coeff[10003] <= 15'b110100011001001;
		Coeff[10004] <= 15'b110100011001011;
		Coeff[10005] <= 15'b110100011001101;
		Coeff[10006] <= 15'b110100011001110;
		Coeff[10007] <= 15'b110100011010000;
		Coeff[10008] <= 15'b110100011010010;
		Coeff[10009] <= 15'b110100011010100;
		Coeff[10010] <= 15'b110100011010110;
		Coeff[10011] <= 15'b110100011010111;
		Coeff[10012] <= 15'b110100011011001;
		Coeff[10013] <= 15'b110100011011011;
		Coeff[10014] <= 15'b110100011011101;
		Coeff[10015] <= 15'b110100011011111;
		Coeff[10016] <= 15'b110100011100000;
		Coeff[10017] <= 15'b110100011100010;
		Coeff[10018] <= 15'b110100011100100;
		Coeff[10019] <= 15'b110100011100110;
		Coeff[10020] <= 15'b110100011101000;
		Coeff[10021] <= 15'b110100011101001;
		Coeff[10022] <= 15'b110100011101011;
		Coeff[10023] <= 15'b110100011101101;
		Coeff[10024] <= 15'b110100011101111;
		Coeff[10025] <= 15'b110100011110001;
		Coeff[10026] <= 15'b110100011110010;
		Coeff[10027] <= 15'b110100011110100;
		Coeff[10028] <= 15'b110100011110110;
		Coeff[10029] <= 15'b110100011111000;
		Coeff[10030] <= 15'b110100011111010;
		Coeff[10031] <= 15'b110100011111011;
		Coeff[10032] <= 15'b110100011111101;
		Coeff[10033] <= 15'b110100011111111;
		Coeff[10034] <= 15'b110100100000001;
		Coeff[10035] <= 15'b110100100000011;
		Coeff[10036] <= 15'b110100100000100;
		Coeff[10037] <= 15'b110100100000110;
		Coeff[10038] <= 15'b110100100001000;
		Coeff[10039] <= 15'b110100100001010;
		Coeff[10040] <= 15'b110100100001100;
		Coeff[10041] <= 15'b110100100001101;
		Coeff[10042] <= 15'b110100100001111;
		Coeff[10043] <= 15'b110100100010001;
		Coeff[10044] <= 15'b110100100010011;
		Coeff[10045] <= 15'b110100100010101;
		Coeff[10046] <= 15'b110100100010110;
		Coeff[10047] <= 15'b110100100011000;
		Coeff[10048] <= 15'b110100100011010;
		Coeff[10049] <= 15'b110100100011100;
		Coeff[10050] <= 15'b110100100011101;
		Coeff[10051] <= 15'b110100100011111;
		Coeff[10052] <= 15'b110100100100001;
		Coeff[10053] <= 15'b110100100100011;
		Coeff[10054] <= 15'b110100100100101;
		Coeff[10055] <= 15'b110100100100110;
		Coeff[10056] <= 15'b110100100101000;
		Coeff[10057] <= 15'b110100100101010;
		Coeff[10058] <= 15'b110100100101100;
		Coeff[10059] <= 15'b110100100101110;
		Coeff[10060] <= 15'b110100100101111;
		Coeff[10061] <= 15'b110100100110001;
		Coeff[10062] <= 15'b110100100110011;
		Coeff[10063] <= 15'b110100100110101;
		Coeff[10064] <= 15'b110100100110111;
		Coeff[10065] <= 15'b110100100111000;
		Coeff[10066] <= 15'b110100100111010;
		Coeff[10067] <= 15'b110100100111100;
		Coeff[10068] <= 15'b110100100111110;
		Coeff[10069] <= 15'b110100100111111;
		Coeff[10070] <= 15'b110100101000001;
		Coeff[10071] <= 15'b110100101000011;
		Coeff[10072] <= 15'b110100101000101;
		Coeff[10073] <= 15'b110100101000111;
		Coeff[10074] <= 15'b110100101001000;
		Coeff[10075] <= 15'b110100101001010;
		Coeff[10076] <= 15'b110100101001100;
		Coeff[10077] <= 15'b110100101001110;
		Coeff[10078] <= 15'b110100101010000;
		Coeff[10079] <= 15'b110100101010001;
		Coeff[10080] <= 15'b110100101010011;
		Coeff[10081] <= 15'b110100101010101;
		Coeff[10082] <= 15'b110100101010111;
		Coeff[10083] <= 15'b110100101011000;
		Coeff[10084] <= 15'b110100101011010;
		Coeff[10085] <= 15'b110100101011100;
		Coeff[10086] <= 15'b110100101011110;
		Coeff[10087] <= 15'b110100101100000;
		Coeff[10088] <= 15'b110100101100001;
		Coeff[10089] <= 15'b110100101100011;
		Coeff[10090] <= 15'b110100101100101;
		Coeff[10091] <= 15'b110100101100111;
		Coeff[10092] <= 15'b110100101101001;
		Coeff[10093] <= 15'b110100101101010;
		Coeff[10094] <= 15'b110100101101100;
		Coeff[10095] <= 15'b110100101101110;
		Coeff[10096] <= 15'b110100101110000;
		Coeff[10097] <= 15'b110100101110001;
		Coeff[10098] <= 15'b110100101110011;
		Coeff[10099] <= 15'b110100101110101;
		Coeff[10100] <= 15'b110100101110111;
		Coeff[10101] <= 15'b110100101111001;
		Coeff[10102] <= 15'b110100101111010;
		Coeff[10103] <= 15'b110100101111100;
		Coeff[10104] <= 15'b110100101111110;
		Coeff[10105] <= 15'b110100110000000;
		Coeff[10106] <= 15'b110100110000001;
		Coeff[10107] <= 15'b110100110000011;
		Coeff[10108] <= 15'b110100110000101;
		Coeff[10109] <= 15'b110100110000111;
		Coeff[10110] <= 15'b110100110001001;
		Coeff[10111] <= 15'b110100110001010;
		Coeff[10112] <= 15'b110100110001100;
		Coeff[10113] <= 15'b110100110001110;
		Coeff[10114] <= 15'b110100110010000;
		Coeff[10115] <= 15'b110100110010001;
		Coeff[10116] <= 15'b110100110010011;
		Coeff[10117] <= 15'b110100110010101;
		Coeff[10118] <= 15'b110100110010111;
		Coeff[10119] <= 15'b110100110011001;
		Coeff[10120] <= 15'b110100110011010;
		Coeff[10121] <= 15'b110100110011100;
		Coeff[10122] <= 15'b110100110011110;
		Coeff[10123] <= 15'b110100110100000;
		Coeff[10124] <= 15'b110100110100001;
		Coeff[10125] <= 15'b110100110100011;
		Coeff[10126] <= 15'b110100110100101;
		Coeff[10127] <= 15'b110100110100111;
		Coeff[10128] <= 15'b110100110101001;
		Coeff[10129] <= 15'b110100110101010;
		Coeff[10130] <= 15'b110100110101100;
		Coeff[10131] <= 15'b110100110101110;
		Coeff[10132] <= 15'b110100110110000;
		Coeff[10133] <= 15'b110100110110001;
		Coeff[10134] <= 15'b110100110110011;
		Coeff[10135] <= 15'b110100110110101;
		Coeff[10136] <= 15'b110100110110111;
		Coeff[10137] <= 15'b110100110111000;
		Coeff[10138] <= 15'b110100110111010;
		Coeff[10139] <= 15'b110100110111100;
		Coeff[10140] <= 15'b110100110111110;
		Coeff[10141] <= 15'b110100111000000;
		Coeff[10142] <= 15'b110100111000001;
		Coeff[10143] <= 15'b110100111000011;
		Coeff[10144] <= 15'b110100111000101;
		Coeff[10145] <= 15'b110100111000111;
		Coeff[10146] <= 15'b110100111001000;
		Coeff[10147] <= 15'b110100111001010;
		Coeff[10148] <= 15'b110100111001100;
		Coeff[10149] <= 15'b110100111001110;
		Coeff[10150] <= 15'b110100111010000;
		Coeff[10151] <= 15'b110100111010001;
		Coeff[10152] <= 15'b110100111010011;
		Coeff[10153] <= 15'b110100111010101;
		Coeff[10154] <= 15'b110100111010111;
		Coeff[10155] <= 15'b110100111011000;
		Coeff[10156] <= 15'b110100111011010;
		Coeff[10157] <= 15'b110100111011100;
		Coeff[10158] <= 15'b110100111011110;
		Coeff[10159] <= 15'b110100111011111;
		Coeff[10160] <= 15'b110100111100001;
		Coeff[10161] <= 15'b110100111100011;
		Coeff[10162] <= 15'b110100111100101;
		Coeff[10163] <= 15'b110100111100110;
		Coeff[10164] <= 15'b110100111101000;
		Coeff[10165] <= 15'b110100111101010;
		Coeff[10166] <= 15'b110100111101100;
		Coeff[10167] <= 15'b110100111101110;
		Coeff[10168] <= 15'b110100111101111;
		Coeff[10169] <= 15'b110100111110001;
		Coeff[10170] <= 15'b110100111110011;
		Coeff[10171] <= 15'b110100111110101;
		Coeff[10172] <= 15'b110100111110110;
		Coeff[10173] <= 15'b110100111111000;
		Coeff[10174] <= 15'b110100111111010;
		Coeff[10175] <= 15'b110100111111100;
		Coeff[10176] <= 15'b110100111111101;
		Coeff[10177] <= 15'b110100111111111;
		Coeff[10178] <= 15'b110101000000001;
		Coeff[10179] <= 15'b110101000000011;
		Coeff[10180] <= 15'b110101000000100;
		Coeff[10181] <= 15'b110101000000110;
		Coeff[10182] <= 15'b110101000001000;
		Coeff[10183] <= 15'b110101000001010;
		Coeff[10184] <= 15'b110101000001011;
		Coeff[10185] <= 15'b110101000001101;
		Coeff[10186] <= 15'b110101000001111;
		Coeff[10187] <= 15'b110101000010001;
		Coeff[10188] <= 15'b110101000010010;
		Coeff[10189] <= 15'b110101000010100;
		Coeff[10190] <= 15'b110101000010110;
		Coeff[10191] <= 15'b110101000011000;
		Coeff[10192] <= 15'b110101000011010;
		Coeff[10193] <= 15'b110101000011011;
		Coeff[10194] <= 15'b110101000011101;
		Coeff[10195] <= 15'b110101000011111;
		Coeff[10196] <= 15'b110101000100001;
		Coeff[10197] <= 15'b110101000100010;
		Coeff[10198] <= 15'b110101000100100;
		Coeff[10199] <= 15'b110101000100110;
		Coeff[10200] <= 15'b110101000101000;
		Coeff[10201] <= 15'b110101000101001;
		Coeff[10202] <= 15'b110101000101011;
		Coeff[10203] <= 15'b110101000101101;
		Coeff[10204] <= 15'b110101000101111;
		Coeff[10205] <= 15'b110101000110000;
		Coeff[10206] <= 15'b110101000110010;
		Coeff[10207] <= 15'b110101000110100;
		Coeff[10208] <= 15'b110101000110110;
		Coeff[10209] <= 15'b110101000110111;
		Coeff[10210] <= 15'b110101000111001;
		Coeff[10211] <= 15'b110101000111011;
		Coeff[10212] <= 15'b110101000111101;
		Coeff[10213] <= 15'b110101000111110;
		Coeff[10214] <= 15'b110101001000000;
		Coeff[10215] <= 15'b110101001000010;
		Coeff[10216] <= 15'b110101001000100;
		Coeff[10217] <= 15'b110101001000101;
		Coeff[10218] <= 15'b110101001000111;
		Coeff[10219] <= 15'b110101001001001;
		Coeff[10220] <= 15'b110101001001011;
		Coeff[10221] <= 15'b110101001001100;
		Coeff[10222] <= 15'b110101001001110;
		Coeff[10223] <= 15'b110101001010000;
		Coeff[10224] <= 15'b110101001010010;
		Coeff[10225] <= 15'b110101001010011;
		Coeff[10226] <= 15'b110101001010101;
		Coeff[10227] <= 15'b110101001010111;
		Coeff[10228] <= 15'b110101001011001;
		Coeff[10229] <= 15'b110101001011010;
		Coeff[10230] <= 15'b110101001011100;
		Coeff[10231] <= 15'b110101001011110;
		Coeff[10232] <= 15'b110101001100000;
		Coeff[10233] <= 15'b110101001100001;
		Coeff[10234] <= 15'b110101001100011;
		Coeff[10235] <= 15'b110101001100101;
		Coeff[10236] <= 15'b110101001100111;
		Coeff[10237] <= 15'b110101001101000;
		Coeff[10238] <= 15'b110101001101010;
		Coeff[10239] <= 15'b110101001101100;
		Coeff[10240] <= 15'b110101001101110;
		Coeff[10241] <= 15'b110101001101111;
		Coeff[10242] <= 15'b110101001110001;
		Coeff[10243] <= 15'b110101001110011;
		Coeff[10244] <= 15'b110101001110101;
		Coeff[10245] <= 15'b110101001110110;
		Coeff[10246] <= 15'b110101001111000;
		Coeff[10247] <= 15'b110101001111010;
		Coeff[10248] <= 15'b110101001111100;
		Coeff[10249] <= 15'b110101001111101;
		Coeff[10250] <= 15'b110101001111111;
		Coeff[10251] <= 15'b110101010000001;
		Coeff[10252] <= 15'b110101010000011;
		Coeff[10253] <= 15'b110101010000100;
		Coeff[10254] <= 15'b110101010000110;
		Coeff[10255] <= 15'b110101010001000;
		Coeff[10256] <= 15'b110101010001001;
		Coeff[10257] <= 15'b110101010001011;
		Coeff[10258] <= 15'b110101010001101;
		Coeff[10259] <= 15'b110101010001111;
		Coeff[10260] <= 15'b110101010010000;
		Coeff[10261] <= 15'b110101010010010;
		Coeff[10262] <= 15'b110101010010100;
		Coeff[10263] <= 15'b110101010010110;
		Coeff[10264] <= 15'b110101010010111;
		Coeff[10265] <= 15'b110101010011001;
		Coeff[10266] <= 15'b110101010011011;
		Coeff[10267] <= 15'b110101010011101;
		Coeff[10268] <= 15'b110101010011110;
		Coeff[10269] <= 15'b110101010100000;
		Coeff[10270] <= 15'b110101010100010;
		Coeff[10271] <= 15'b110101010100100;
		Coeff[10272] <= 15'b110101010100101;
		Coeff[10273] <= 15'b110101010100111;
		Coeff[10274] <= 15'b110101010101001;
		Coeff[10275] <= 15'b110101010101011;
		Coeff[10276] <= 15'b110101010101100;
		Coeff[10277] <= 15'b110101010101110;
		Coeff[10278] <= 15'b110101010110000;
		Coeff[10279] <= 15'b110101010110001;
		Coeff[10280] <= 15'b110101010110011;
		Coeff[10281] <= 15'b110101010110101;
		Coeff[10282] <= 15'b110101010110111;
		Coeff[10283] <= 15'b110101010111000;
		Coeff[10284] <= 15'b110101010111010;
		Coeff[10285] <= 15'b110101010111100;
		Coeff[10286] <= 15'b110101010111110;
		Coeff[10287] <= 15'b110101010111111;
		Coeff[10288] <= 15'b110101011000001;
		Coeff[10289] <= 15'b110101011000011;
		Coeff[10290] <= 15'b110101011000101;
		Coeff[10291] <= 15'b110101011000110;
		Coeff[10292] <= 15'b110101011001000;
		Coeff[10293] <= 15'b110101011001010;
		Coeff[10294] <= 15'b110101011001011;
		Coeff[10295] <= 15'b110101011001101;
		Coeff[10296] <= 15'b110101011001111;
		Coeff[10297] <= 15'b110101011010001;
		Coeff[10298] <= 15'b110101011010010;
		Coeff[10299] <= 15'b110101011010100;
		Coeff[10300] <= 15'b110101011010110;
		Coeff[10301] <= 15'b110101011011000;
		Coeff[10302] <= 15'b110101011011001;
		Coeff[10303] <= 15'b110101011011011;
		Coeff[10304] <= 15'b110101011011101;
		Coeff[10305] <= 15'b110101011011111;
		Coeff[10306] <= 15'b110101011100000;
		Coeff[10307] <= 15'b110101011100010;
		Coeff[10308] <= 15'b110101011100100;
		Coeff[10309] <= 15'b110101011100101;
		Coeff[10310] <= 15'b110101011100111;
		Coeff[10311] <= 15'b110101011101001;
		Coeff[10312] <= 15'b110101011101011;
		Coeff[10313] <= 15'b110101011101100;
		Coeff[10314] <= 15'b110101011101110;
		Coeff[10315] <= 15'b110101011110000;
		Coeff[10316] <= 15'b110101011110010;
		Coeff[10317] <= 15'b110101011110011;
		Coeff[10318] <= 15'b110101011110101;
		Coeff[10319] <= 15'b110101011110111;
		Coeff[10320] <= 15'b110101011111000;
		Coeff[10321] <= 15'b110101011111010;
		Coeff[10322] <= 15'b110101011111100;
		Coeff[10323] <= 15'b110101011111110;
		Coeff[10324] <= 15'b110101011111111;
		Coeff[10325] <= 15'b110101100000001;
		Coeff[10326] <= 15'b110101100000011;
		Coeff[10327] <= 15'b110101100000100;
		Coeff[10328] <= 15'b110101100000110;
		Coeff[10329] <= 15'b110101100001000;
		Coeff[10330] <= 15'b110101100001010;
		Coeff[10331] <= 15'b110101100001011;
		Coeff[10332] <= 15'b110101100001101;
		Coeff[10333] <= 15'b110101100001111;
		Coeff[10334] <= 15'b110101100010001;
		Coeff[10335] <= 15'b110101100010010;
		Coeff[10336] <= 15'b110101100010100;
		Coeff[10337] <= 15'b110101100010110;
		Coeff[10338] <= 15'b110101100010111;
		Coeff[10339] <= 15'b110101100011001;
		Coeff[10340] <= 15'b110101100011011;
		Coeff[10341] <= 15'b110101100011101;
		Coeff[10342] <= 15'b110101100011110;
		Coeff[10343] <= 15'b110101100100000;
		Coeff[10344] <= 15'b110101100100010;
		Coeff[10345] <= 15'b110101100100011;
		Coeff[10346] <= 15'b110101100100101;
		Coeff[10347] <= 15'b110101100100111;
		Coeff[10348] <= 15'b110101100101001;
		Coeff[10349] <= 15'b110101100101010;
		Coeff[10350] <= 15'b110101100101100;
		Coeff[10351] <= 15'b110101100101110;
		Coeff[10352] <= 15'b110101100110000;
		Coeff[10353] <= 15'b110101100110001;
		Coeff[10354] <= 15'b110101100110011;
		Coeff[10355] <= 15'b110101100110101;
		Coeff[10356] <= 15'b110101100110110;
		Coeff[10357] <= 15'b110101100111000;
		Coeff[10358] <= 15'b110101100111010;
		Coeff[10359] <= 15'b110101100111100;
		Coeff[10360] <= 15'b110101100111101;
		Coeff[10361] <= 15'b110101100111111;
		Coeff[10362] <= 15'b110101101000001;
		Coeff[10363] <= 15'b110101101000010;
		Coeff[10364] <= 15'b110101101000100;
		Coeff[10365] <= 15'b110101101000110;
		Coeff[10366] <= 15'b110101101001000;
		Coeff[10367] <= 15'b110101101001001;
		Coeff[10368] <= 15'b110101101001011;
		Coeff[10369] <= 15'b110101101001101;
		Coeff[10370] <= 15'b110101101001110;
		Coeff[10371] <= 15'b110101101010000;
		Coeff[10372] <= 15'b110101101010010;
		Coeff[10373] <= 15'b110101101010100;
		Coeff[10374] <= 15'b110101101010101;
		Coeff[10375] <= 15'b110101101010111;
		Coeff[10376] <= 15'b110101101011001;
		Coeff[10377] <= 15'b110101101011010;
		Coeff[10378] <= 15'b110101101011100;
		Coeff[10379] <= 15'b110101101011110;
		Coeff[10380] <= 15'b110101101011111;
		Coeff[10381] <= 15'b110101101100001;
		Coeff[10382] <= 15'b110101101100011;
		Coeff[10383] <= 15'b110101101100101;
		Coeff[10384] <= 15'b110101101100110;
		Coeff[10385] <= 15'b110101101101000;
		Coeff[10386] <= 15'b110101101101010;
		Coeff[10387] <= 15'b110101101101011;
		Coeff[10388] <= 15'b110101101101101;
		Coeff[10389] <= 15'b110101101101111;
		Coeff[10390] <= 15'b110101101110001;
		Coeff[10391] <= 15'b110101101110010;
		Coeff[10392] <= 15'b110101101110100;
		Coeff[10393] <= 15'b110101101110110;
		Coeff[10394] <= 15'b110101101110111;
		Coeff[10395] <= 15'b110101101111001;
		Coeff[10396] <= 15'b110101101111011;
		Coeff[10397] <= 15'b110101101111101;
		Coeff[10398] <= 15'b110101101111110;
		Coeff[10399] <= 15'b110101110000000;
		Coeff[10400] <= 15'b110101110000010;
		Coeff[10401] <= 15'b110101110000011;
		Coeff[10402] <= 15'b110101110000101;
		Coeff[10403] <= 15'b110101110000111;
		Coeff[10404] <= 15'b110101110001000;
		Coeff[10405] <= 15'b110101110001010;
		Coeff[10406] <= 15'b110101110001100;
		Coeff[10407] <= 15'b110101110001110;
		Coeff[10408] <= 15'b110101110001111;
		Coeff[10409] <= 15'b110101110010001;
		Coeff[10410] <= 15'b110101110010011;
		Coeff[10411] <= 15'b110101110010100;
		Coeff[10412] <= 15'b110101110010110;
		Coeff[10413] <= 15'b110101110011000;
		Coeff[10414] <= 15'b110101110011001;
		Coeff[10415] <= 15'b110101110011011;
		Coeff[10416] <= 15'b110101110011101;
		Coeff[10417] <= 15'b110101110011111;
		Coeff[10418] <= 15'b110101110100000;
		Coeff[10419] <= 15'b110101110100010;
		Coeff[10420] <= 15'b110101110100100;
		Coeff[10421] <= 15'b110101110100101;
		Coeff[10422] <= 15'b110101110100111;
		Coeff[10423] <= 15'b110101110101001;
		Coeff[10424] <= 15'b110101110101010;
		Coeff[10425] <= 15'b110101110101100;
		Coeff[10426] <= 15'b110101110101110;
		Coeff[10427] <= 15'b110101110110000;
		Coeff[10428] <= 15'b110101110110001;
		Coeff[10429] <= 15'b110101110110011;
		Coeff[10430] <= 15'b110101110110101;
		Coeff[10431] <= 15'b110101110110110;
		Coeff[10432] <= 15'b110101110111000;
		Coeff[10433] <= 15'b110101110111010;
		Coeff[10434] <= 15'b110101110111011;
		Coeff[10435] <= 15'b110101110111101;
		Coeff[10436] <= 15'b110101110111111;
		Coeff[10437] <= 15'b110101111000001;
		Coeff[10438] <= 15'b110101111000010;
		Coeff[10439] <= 15'b110101111000100;
		Coeff[10440] <= 15'b110101111000110;
		Coeff[10441] <= 15'b110101111000111;
		Coeff[10442] <= 15'b110101111001001;
		Coeff[10443] <= 15'b110101111001011;
		Coeff[10444] <= 15'b110101111001100;
		Coeff[10445] <= 15'b110101111001110;
		Coeff[10446] <= 15'b110101111010000;
		Coeff[10447] <= 15'b110101111010001;
		Coeff[10448] <= 15'b110101111010011;
		Coeff[10449] <= 15'b110101111010101;
		Coeff[10450] <= 15'b110101111010111;
		Coeff[10451] <= 15'b110101111011000;
		Coeff[10452] <= 15'b110101111011010;
		Coeff[10453] <= 15'b110101111011100;
		Coeff[10454] <= 15'b110101111011101;
		Coeff[10455] <= 15'b110101111011111;
		Coeff[10456] <= 15'b110101111100001;
		Coeff[10457] <= 15'b110101111100010;
		Coeff[10458] <= 15'b110101111100100;
		Coeff[10459] <= 15'b110101111100110;
		Coeff[10460] <= 15'b110101111100111;
		Coeff[10461] <= 15'b110101111101001;
		Coeff[10462] <= 15'b110101111101011;
		Coeff[10463] <= 15'b110101111101101;
		Coeff[10464] <= 15'b110101111101110;
		Coeff[10465] <= 15'b110101111110000;
		Coeff[10466] <= 15'b110101111110010;
		Coeff[10467] <= 15'b110101111110011;
		Coeff[10468] <= 15'b110101111110101;
		Coeff[10469] <= 15'b110101111110111;
		Coeff[10470] <= 15'b110101111111000;
		Coeff[10471] <= 15'b110101111111010;
		Coeff[10472] <= 15'b110101111111100;
		Coeff[10473] <= 15'b110101111111101;
		Coeff[10474] <= 15'b110101111111111;
		Coeff[10475] <= 15'b110110000000001;
		Coeff[10476] <= 15'b110110000000010;
		Coeff[10477] <= 15'b110110000000100;
		Coeff[10478] <= 15'b110110000000110;
		Coeff[10479] <= 15'b110110000001000;
		Coeff[10480] <= 15'b110110000001001;
		Coeff[10481] <= 15'b110110000001011;
		Coeff[10482] <= 15'b110110000001101;
		Coeff[10483] <= 15'b110110000001110;
		Coeff[10484] <= 15'b110110000010000;
		Coeff[10485] <= 15'b110110000010010;
		Coeff[10486] <= 15'b110110000010011;
		Coeff[10487] <= 15'b110110000010101;
		Coeff[10488] <= 15'b110110000010111;
		Coeff[10489] <= 15'b110110000011000;
		Coeff[10490] <= 15'b110110000011010;
		Coeff[10491] <= 15'b110110000011100;
		Coeff[10492] <= 15'b110110000011101;
		Coeff[10493] <= 15'b110110000011111;
		Coeff[10494] <= 15'b110110000100001;
		Coeff[10495] <= 15'b110110000100010;
		Coeff[10496] <= 15'b110110000100100;
		Coeff[10497] <= 15'b110110000100110;
		Coeff[10498] <= 15'b110110000101000;
		Coeff[10499] <= 15'b110110000101001;
		Coeff[10500] <= 15'b110110000101011;
		Coeff[10501] <= 15'b110110000101101;
		Coeff[10502] <= 15'b110110000101110;
		Coeff[10503] <= 15'b110110000110000;
		Coeff[10504] <= 15'b110110000110010;
		Coeff[10505] <= 15'b110110000110011;
		Coeff[10506] <= 15'b110110000110101;
		Coeff[10507] <= 15'b110110000110111;
		Coeff[10508] <= 15'b110110000111000;
		Coeff[10509] <= 15'b110110000111010;
		Coeff[10510] <= 15'b110110000111100;
		Coeff[10511] <= 15'b110110000111101;
		Coeff[10512] <= 15'b110110000111111;
		Coeff[10513] <= 15'b110110001000001;
		Coeff[10514] <= 15'b110110001000010;
		Coeff[10515] <= 15'b110110001000100;
		Coeff[10516] <= 15'b110110001000110;
		Coeff[10517] <= 15'b110110001000111;
		Coeff[10518] <= 15'b110110001001001;
		Coeff[10519] <= 15'b110110001001011;
		Coeff[10520] <= 15'b110110001001100;
		Coeff[10521] <= 15'b110110001001110;
		Coeff[10522] <= 15'b110110001010000;
		Coeff[10523] <= 15'b110110001010001;
		Coeff[10524] <= 15'b110110001010011;
		Coeff[10525] <= 15'b110110001010101;
		Coeff[10526] <= 15'b110110001010110;
		Coeff[10527] <= 15'b110110001011000;
		Coeff[10528] <= 15'b110110001011010;
		Coeff[10529] <= 15'b110110001011011;
		Coeff[10530] <= 15'b110110001011101;
		Coeff[10531] <= 15'b110110001011111;
		Coeff[10532] <= 15'b110110001100001;
		Coeff[10533] <= 15'b110110001100010;
		Coeff[10534] <= 15'b110110001100100;
		Coeff[10535] <= 15'b110110001100110;
		Coeff[10536] <= 15'b110110001100111;
		Coeff[10537] <= 15'b110110001101001;
		Coeff[10538] <= 15'b110110001101011;
		Coeff[10539] <= 15'b110110001101100;
		Coeff[10540] <= 15'b110110001101110;
		Coeff[10541] <= 15'b110110001110000;
		Coeff[10542] <= 15'b110110001110001;
		Coeff[10543] <= 15'b110110001110011;
		Coeff[10544] <= 15'b110110001110101;
		Coeff[10545] <= 15'b110110001110110;
		Coeff[10546] <= 15'b110110001111000;
		Coeff[10547] <= 15'b110110001111010;
		Coeff[10548] <= 15'b110110001111011;
		Coeff[10549] <= 15'b110110001111101;
		Coeff[10550] <= 15'b110110001111111;
		Coeff[10551] <= 15'b110110010000000;
		Coeff[10552] <= 15'b110110010000010;
		Coeff[10553] <= 15'b110110010000100;
		Coeff[10554] <= 15'b110110010000101;
		Coeff[10555] <= 15'b110110010000111;
		Coeff[10556] <= 15'b110110010001001;
		Coeff[10557] <= 15'b110110010001010;
		Coeff[10558] <= 15'b110110010001100;
		Coeff[10559] <= 15'b110110010001110;
		Coeff[10560] <= 15'b110110010001111;
		Coeff[10561] <= 15'b110110010010001;
		Coeff[10562] <= 15'b110110010010011;
		Coeff[10563] <= 15'b110110010010100;
		Coeff[10564] <= 15'b110110010010110;
		Coeff[10565] <= 15'b110110010011000;
		Coeff[10566] <= 15'b110110010011001;
		Coeff[10567] <= 15'b110110010011011;
		Coeff[10568] <= 15'b110110010011101;
		Coeff[10569] <= 15'b110110010011110;
		Coeff[10570] <= 15'b110110010100000;
		Coeff[10571] <= 15'b110110010100010;
		Coeff[10572] <= 15'b110110010100011;
		Coeff[10573] <= 15'b110110010100101;
		Coeff[10574] <= 15'b110110010100110;
		Coeff[10575] <= 15'b110110010101000;
		Coeff[10576] <= 15'b110110010101010;
		Coeff[10577] <= 15'b110110010101011;
		Coeff[10578] <= 15'b110110010101101;
		Coeff[10579] <= 15'b110110010101111;
		Coeff[10580] <= 15'b110110010110000;
		Coeff[10581] <= 15'b110110010110010;
		Coeff[10582] <= 15'b110110010110100;
		Coeff[10583] <= 15'b110110010110101;
		Coeff[10584] <= 15'b110110010110111;
		Coeff[10585] <= 15'b110110010111001;
		Coeff[10586] <= 15'b110110010111010;
		Coeff[10587] <= 15'b110110010111100;
		Coeff[10588] <= 15'b110110010111110;
		Coeff[10589] <= 15'b110110010111111;
		Coeff[10590] <= 15'b110110011000001;
		Coeff[10591] <= 15'b110110011000011;
		Coeff[10592] <= 15'b110110011000100;
		Coeff[10593] <= 15'b110110011000110;
		Coeff[10594] <= 15'b110110011001000;
		Coeff[10595] <= 15'b110110011001001;
		Coeff[10596] <= 15'b110110011001011;
		Coeff[10597] <= 15'b110110011001101;
		Coeff[10598] <= 15'b110110011001110;
		Coeff[10599] <= 15'b110110011010000;
		Coeff[10600] <= 15'b110110011010010;
		Coeff[10601] <= 15'b110110011010011;
		Coeff[10602] <= 15'b110110011010101;
		Coeff[10603] <= 15'b110110011010111;
		Coeff[10604] <= 15'b110110011011000;
		Coeff[10605] <= 15'b110110011011010;
		Coeff[10606] <= 15'b110110011011100;
		Coeff[10607] <= 15'b110110011011101;
		Coeff[10608] <= 15'b110110011011111;
		Coeff[10609] <= 15'b110110011100000;
		Coeff[10610] <= 15'b110110011100010;
		Coeff[10611] <= 15'b110110011100100;
		Coeff[10612] <= 15'b110110011100101;
		Coeff[10613] <= 15'b110110011100111;
		Coeff[10614] <= 15'b110110011101001;
		Coeff[10615] <= 15'b110110011101010;
		Coeff[10616] <= 15'b110110011101100;
		Coeff[10617] <= 15'b110110011101110;
		Coeff[10618] <= 15'b110110011101111;
		Coeff[10619] <= 15'b110110011110001;
		Coeff[10620] <= 15'b110110011110011;
		Coeff[10621] <= 15'b110110011110100;
		Coeff[10622] <= 15'b110110011110110;
		Coeff[10623] <= 15'b110110011111000;
		Coeff[10624] <= 15'b110110011111001;
		Coeff[10625] <= 15'b110110011111011;
		Coeff[10626] <= 15'b110110011111101;
		Coeff[10627] <= 15'b110110011111110;
		Coeff[10628] <= 15'b110110100000000;
		Coeff[10629] <= 15'b110110100000001;
		Coeff[10630] <= 15'b110110100000011;
		Coeff[10631] <= 15'b110110100000101;
		Coeff[10632] <= 15'b110110100000110;
		Coeff[10633] <= 15'b110110100001000;
		Coeff[10634] <= 15'b110110100001010;
		Coeff[10635] <= 15'b110110100001011;
		Coeff[10636] <= 15'b110110100001101;
		Coeff[10637] <= 15'b110110100001111;
		Coeff[10638] <= 15'b110110100010000;
		Coeff[10639] <= 15'b110110100010010;
		Coeff[10640] <= 15'b110110100010100;
		Coeff[10641] <= 15'b110110100010101;
		Coeff[10642] <= 15'b110110100010111;
		Coeff[10643] <= 15'b110110100011000;
		Coeff[10644] <= 15'b110110100011010;
		Coeff[10645] <= 15'b110110100011100;
		Coeff[10646] <= 15'b110110100011101;
		Coeff[10647] <= 15'b110110100011111;
		Coeff[10648] <= 15'b110110100100001;
		Coeff[10649] <= 15'b110110100100010;
		Coeff[10650] <= 15'b110110100100100;
		Coeff[10651] <= 15'b110110100100110;
		Coeff[10652] <= 15'b110110100100111;
		Coeff[10653] <= 15'b110110100101001;
		Coeff[10654] <= 15'b110110100101011;
		Coeff[10655] <= 15'b110110100101100;
		Coeff[10656] <= 15'b110110100101110;
		Coeff[10657] <= 15'b110110100101111;
		Coeff[10658] <= 15'b110110100110001;
		Coeff[10659] <= 15'b110110100110011;
		Coeff[10660] <= 15'b110110100110100;
		Coeff[10661] <= 15'b110110100110110;
		Coeff[10662] <= 15'b110110100111000;
		Coeff[10663] <= 15'b110110100111001;
		Coeff[10664] <= 15'b110110100111011;
		Coeff[10665] <= 15'b110110100111101;
		Coeff[10666] <= 15'b110110100111110;
		Coeff[10667] <= 15'b110110101000000;
		Coeff[10668] <= 15'b110110101000001;
		Coeff[10669] <= 15'b110110101000011;
		Coeff[10670] <= 15'b110110101000101;
		Coeff[10671] <= 15'b110110101000110;
		Coeff[10672] <= 15'b110110101001000;
		Coeff[10673] <= 15'b110110101001010;
		Coeff[10674] <= 15'b110110101001011;
		Coeff[10675] <= 15'b110110101001101;
		Coeff[10676] <= 15'b110110101001111;
		Coeff[10677] <= 15'b110110101010000;
		Coeff[10678] <= 15'b110110101010010;
		Coeff[10679] <= 15'b110110101010011;
		Coeff[10680] <= 15'b110110101010101;
		Coeff[10681] <= 15'b110110101010111;
		Coeff[10682] <= 15'b110110101011000;
		Coeff[10683] <= 15'b110110101011010;
		Coeff[10684] <= 15'b110110101011100;
		Coeff[10685] <= 15'b110110101011101;
		Coeff[10686] <= 15'b110110101011111;
		Coeff[10687] <= 15'b110110101100001;
		Coeff[10688] <= 15'b110110101100010;
		Coeff[10689] <= 15'b110110101100100;
		Coeff[10690] <= 15'b110110101100101;
		Coeff[10691] <= 15'b110110101100111;
		Coeff[10692] <= 15'b110110101101001;
		Coeff[10693] <= 15'b110110101101010;
		Coeff[10694] <= 15'b110110101101100;
		Coeff[10695] <= 15'b110110101101110;
		Coeff[10696] <= 15'b110110101101111;
		Coeff[10697] <= 15'b110110101110001;
		Coeff[10698] <= 15'b110110101110010;
		Coeff[10699] <= 15'b110110101110100;
		Coeff[10700] <= 15'b110110101110110;
		Coeff[10701] <= 15'b110110101110111;
		Coeff[10702] <= 15'b110110101111001;
		Coeff[10703] <= 15'b110110101111011;
		Coeff[10704] <= 15'b110110101111100;
		Coeff[10705] <= 15'b110110101111110;
		Coeff[10706] <= 15'b110110101111111;
		Coeff[10707] <= 15'b110110110000001;
		Coeff[10708] <= 15'b110110110000011;
		Coeff[10709] <= 15'b110110110000100;
		Coeff[10710] <= 15'b110110110000110;
		Coeff[10711] <= 15'b110110110001000;
		Coeff[10712] <= 15'b110110110001001;
		Coeff[10713] <= 15'b110110110001011;
		Coeff[10714] <= 15'b110110110001100;
		Coeff[10715] <= 15'b110110110001110;
		Coeff[10716] <= 15'b110110110010000;
		Coeff[10717] <= 15'b110110110010001;
		Coeff[10718] <= 15'b110110110010011;
		Coeff[10719] <= 15'b110110110010101;
		Coeff[10720] <= 15'b110110110010110;
		Coeff[10721] <= 15'b110110110011000;
		Coeff[10722] <= 15'b110110110011001;
		Coeff[10723] <= 15'b110110110011011;
		Coeff[10724] <= 15'b110110110011101;
		Coeff[10725] <= 15'b110110110011110;
		Coeff[10726] <= 15'b110110110100000;
		Coeff[10727] <= 15'b110110110100010;
		Coeff[10728] <= 15'b110110110100011;
		Coeff[10729] <= 15'b110110110100101;
		Coeff[10730] <= 15'b110110110100110;
		Coeff[10731] <= 15'b110110110101000;
		Coeff[10732] <= 15'b110110110101010;
		Coeff[10733] <= 15'b110110110101011;
		Coeff[10734] <= 15'b110110110101101;
		Coeff[10735] <= 15'b110110110101111;
		Coeff[10736] <= 15'b110110110110000;
		Coeff[10737] <= 15'b110110110110010;
		Coeff[10738] <= 15'b110110110110011;
		Coeff[10739] <= 15'b110110110110101;
		Coeff[10740] <= 15'b110110110110111;
		Coeff[10741] <= 15'b110110110111000;
		Coeff[10742] <= 15'b110110110111010;
		Coeff[10743] <= 15'b110110110111100;
		Coeff[10744] <= 15'b110110110111101;
		Coeff[10745] <= 15'b110110110111111;
		Coeff[10746] <= 15'b110110111000000;
		Coeff[10747] <= 15'b110110111000010;
		Coeff[10748] <= 15'b110110111000100;
		Coeff[10749] <= 15'b110110111000101;
		Coeff[10750] <= 15'b110110111000111;
		Coeff[10751] <= 15'b110110111001000;
		Coeff[10752] <= 15'b110110111001010;
		Coeff[10753] <= 15'b110110111001100;
		Coeff[10754] <= 15'b110110111001101;
		Coeff[10755] <= 15'b110110111001111;
		Coeff[10756] <= 15'b110110111010001;
		Coeff[10757] <= 15'b110110111010010;
		Coeff[10758] <= 15'b110110111010100;
		Coeff[10759] <= 15'b110110111010101;
		Coeff[10760] <= 15'b110110111010111;
		Coeff[10761] <= 15'b110110111011001;
		Coeff[10762] <= 15'b110110111011010;
		Coeff[10763] <= 15'b110110111011100;
		Coeff[10764] <= 15'b110110111011101;
		Coeff[10765] <= 15'b110110111011111;
		Coeff[10766] <= 15'b110110111100001;
		Coeff[10767] <= 15'b110110111100010;
		Coeff[10768] <= 15'b110110111100100;
		Coeff[10769] <= 15'b110110111100101;
		Coeff[10770] <= 15'b110110111100111;
		Coeff[10771] <= 15'b110110111101001;
		Coeff[10772] <= 15'b110110111101010;
		Coeff[10773] <= 15'b110110111101100;
		Coeff[10774] <= 15'b110110111101110;
		Coeff[10775] <= 15'b110110111101111;
		Coeff[10776] <= 15'b110110111110001;
		Coeff[10777] <= 15'b110110111110010;
		Coeff[10778] <= 15'b110110111110100;
		Coeff[10779] <= 15'b110110111110110;
		Coeff[10780] <= 15'b110110111110111;
		Coeff[10781] <= 15'b110110111111001;
		Coeff[10782] <= 15'b110110111111010;
		Coeff[10783] <= 15'b110110111111100;
		Coeff[10784] <= 15'b110110111111110;
		Coeff[10785] <= 15'b110110111111111;
		Coeff[10786] <= 15'b110111000000001;
		Coeff[10787] <= 15'b110111000000010;
		Coeff[10788] <= 15'b110111000000100;
		Coeff[10789] <= 15'b110111000000110;
		Coeff[10790] <= 15'b110111000000111;
		Coeff[10791] <= 15'b110111000001001;
		Coeff[10792] <= 15'b110111000001010;
		Coeff[10793] <= 15'b110111000001100;
		Coeff[10794] <= 15'b110111000001110;
		Coeff[10795] <= 15'b110111000001111;
		Coeff[10796] <= 15'b110111000010001;
		Coeff[10797] <= 15'b110111000010010;
		Coeff[10798] <= 15'b110111000010100;
		Coeff[10799] <= 15'b110111000010110;
		Coeff[10800] <= 15'b110111000010111;
		Coeff[10801] <= 15'b110111000011001;
		Coeff[10802] <= 15'b110111000011010;
		Coeff[10803] <= 15'b110111000011100;
		Coeff[10804] <= 15'b110111000011110;
		Coeff[10805] <= 15'b110111000011111;
		Coeff[10806] <= 15'b110111000100001;
		Coeff[10807] <= 15'b110111000100010;
		Coeff[10808] <= 15'b110111000100100;
		Coeff[10809] <= 15'b110111000100110;
		Coeff[10810] <= 15'b110111000100111;
		Coeff[10811] <= 15'b110111000101001;
		Coeff[10812] <= 15'b110111000101010;
		Coeff[10813] <= 15'b110111000101100;
		Coeff[10814] <= 15'b110111000101110;
		Coeff[10815] <= 15'b110111000101111;
		Coeff[10816] <= 15'b110111000110001;
		Coeff[10817] <= 15'b110111000110010;
		Coeff[10818] <= 15'b110111000110100;
		Coeff[10819] <= 15'b110111000110110;
		Coeff[10820] <= 15'b110111000110111;
		Coeff[10821] <= 15'b110111000111001;
		Coeff[10822] <= 15'b110111000111010;
		Coeff[10823] <= 15'b110111000111100;
		Coeff[10824] <= 15'b110111000111110;
		Coeff[10825] <= 15'b110111000111111;
		Coeff[10826] <= 15'b110111001000001;
		Coeff[10827] <= 15'b110111001000010;
		Coeff[10828] <= 15'b110111001000100;
		Coeff[10829] <= 15'b110111001000110;
		Coeff[10830] <= 15'b110111001000111;
		Coeff[10831] <= 15'b110111001001001;
		Coeff[10832] <= 15'b110111001001010;
		Coeff[10833] <= 15'b110111001001100;
		Coeff[10834] <= 15'b110111001001110;
		Coeff[10835] <= 15'b110111001001111;
		Coeff[10836] <= 15'b110111001010001;
		Coeff[10837] <= 15'b110111001010010;
		Coeff[10838] <= 15'b110111001010100;
		Coeff[10839] <= 15'b110111001010110;
		Coeff[10840] <= 15'b110111001010111;
		Coeff[10841] <= 15'b110111001011001;
		Coeff[10842] <= 15'b110111001011010;
		Coeff[10843] <= 15'b110111001011100;
		Coeff[10844] <= 15'b110111001011110;
		Coeff[10845] <= 15'b110111001011111;
		Coeff[10846] <= 15'b110111001100001;
		Coeff[10847] <= 15'b110111001100010;
		Coeff[10848] <= 15'b110111001100100;
		Coeff[10849] <= 15'b110111001100101;
		Coeff[10850] <= 15'b110111001100111;
		Coeff[10851] <= 15'b110111001101001;
		Coeff[10852] <= 15'b110111001101010;
		Coeff[10853] <= 15'b110111001101100;
		Coeff[10854] <= 15'b110111001101101;
		Coeff[10855] <= 15'b110111001101111;
		Coeff[10856] <= 15'b110111001110001;
		Coeff[10857] <= 15'b110111001110010;
		Coeff[10858] <= 15'b110111001110100;
		Coeff[10859] <= 15'b110111001110101;
		Coeff[10860] <= 15'b110111001110111;
		Coeff[10861] <= 15'b110111001111001;
		Coeff[10862] <= 15'b110111001111010;
		Coeff[10863] <= 15'b110111001111100;
		Coeff[10864] <= 15'b110111001111101;
		Coeff[10865] <= 15'b110111001111111;
		Coeff[10866] <= 15'b110111010000000;
		Coeff[10867] <= 15'b110111010000010;
		Coeff[10868] <= 15'b110111010000100;
		Coeff[10869] <= 15'b110111010000101;
		Coeff[10870] <= 15'b110111010000111;
		Coeff[10871] <= 15'b110111010001000;
		Coeff[10872] <= 15'b110111010001010;
		Coeff[10873] <= 15'b110111010001100;
		Coeff[10874] <= 15'b110111010001101;
		Coeff[10875] <= 15'b110111010001111;
		Coeff[10876] <= 15'b110111010010000;
		Coeff[10877] <= 15'b110111010010010;
		Coeff[10878] <= 15'b110111010010011;
		Coeff[10879] <= 15'b110111010010101;
		Coeff[10880] <= 15'b110111010010111;
		Coeff[10881] <= 15'b110111010011000;
		Coeff[10882] <= 15'b110111010011010;
		Coeff[10883] <= 15'b110111010011011;
		Coeff[10884] <= 15'b110111010011101;
		Coeff[10885] <= 15'b110111010011111;
		Coeff[10886] <= 15'b110111010100000;
		Coeff[10887] <= 15'b110111010100010;
		Coeff[10888] <= 15'b110111010100011;
		Coeff[10889] <= 15'b110111010100101;
		Coeff[10890] <= 15'b110111010100110;
		Coeff[10891] <= 15'b110111010101000;
		Coeff[10892] <= 15'b110111010101010;
		Coeff[10893] <= 15'b110111010101011;
		Coeff[10894] <= 15'b110111010101101;
		Coeff[10895] <= 15'b110111010101110;
		Coeff[10896] <= 15'b110111010110000;
		Coeff[10897] <= 15'b110111010110010;
		Coeff[10898] <= 15'b110111010110011;
		Coeff[10899] <= 15'b110111010110101;
		Coeff[10900] <= 15'b110111010110110;
		Coeff[10901] <= 15'b110111010111000;
		Coeff[10902] <= 15'b110111010111001;
		Coeff[10903] <= 15'b110111010111011;
		Coeff[10904] <= 15'b110111010111101;
		Coeff[10905] <= 15'b110111010111110;
		Coeff[10906] <= 15'b110111011000000;
		Coeff[10907] <= 15'b110111011000001;
		Coeff[10908] <= 15'b110111011000011;
		Coeff[10909] <= 15'b110111011000100;
		Coeff[10910] <= 15'b110111011000110;
		Coeff[10911] <= 15'b110111011001000;
		Coeff[10912] <= 15'b110111011001001;
		Coeff[10913] <= 15'b110111011001011;
		Coeff[10914] <= 15'b110111011001100;
		Coeff[10915] <= 15'b110111011001110;
		Coeff[10916] <= 15'b110111011001111;
		Coeff[10917] <= 15'b110111011010001;
		Coeff[10918] <= 15'b110111011010011;
		Coeff[10919] <= 15'b110111011010100;
		Coeff[10920] <= 15'b110111011010110;
		Coeff[10921] <= 15'b110111011010111;
		Coeff[10922] <= 15'b110111011011001;
		Coeff[10923] <= 15'b110111011011010;
		Coeff[10924] <= 15'b110111011011100;
		Coeff[10925] <= 15'b110111011011110;
		Coeff[10926] <= 15'b110111011011111;
		Coeff[10927] <= 15'b110111011100001;
		Coeff[10928] <= 15'b110111011100010;
		Coeff[10929] <= 15'b110111011100100;
		Coeff[10930] <= 15'b110111011100101;
		Coeff[10931] <= 15'b110111011100111;
		Coeff[10932] <= 15'b110111011101001;
		Coeff[10933] <= 15'b110111011101010;
		Coeff[10934] <= 15'b110111011101100;
		Coeff[10935] <= 15'b110111011101101;
		Coeff[10936] <= 15'b110111011101111;
		Coeff[10937] <= 15'b110111011110000;
		Coeff[10938] <= 15'b110111011110010;
		Coeff[10939] <= 15'b110111011110100;
		Coeff[10940] <= 15'b110111011110101;
		Coeff[10941] <= 15'b110111011110111;
		Coeff[10942] <= 15'b110111011111000;
		Coeff[10943] <= 15'b110111011111010;
		Coeff[10944] <= 15'b110111011111011;
		Coeff[10945] <= 15'b110111011111101;
		Coeff[10946] <= 15'b110111011111111;
		Coeff[10947] <= 15'b110111100000000;
		Coeff[10948] <= 15'b110111100000010;
		Coeff[10949] <= 15'b110111100000011;
		Coeff[10950] <= 15'b110111100000101;
		Coeff[10951] <= 15'b110111100000110;
		Coeff[10952] <= 15'b110111100001000;
		Coeff[10953] <= 15'b110111100001001;
		Coeff[10954] <= 15'b110111100001011;
		Coeff[10955] <= 15'b110111100001101;
		Coeff[10956] <= 15'b110111100001110;
		Coeff[10957] <= 15'b110111100010000;
		Coeff[10958] <= 15'b110111100010001;
		Coeff[10959] <= 15'b110111100010011;
		Coeff[10960] <= 15'b110111100010100;
		Coeff[10961] <= 15'b110111100010110;
		Coeff[10962] <= 15'b110111100011000;
		Coeff[10963] <= 15'b110111100011001;
		Coeff[10964] <= 15'b110111100011011;
		Coeff[10965] <= 15'b110111100011100;
		Coeff[10966] <= 15'b110111100011110;
		Coeff[10967] <= 15'b110111100011111;
		Coeff[10968] <= 15'b110111100100001;
		Coeff[10969] <= 15'b110111100100010;
		Coeff[10970] <= 15'b110111100100100;
		Coeff[10971] <= 15'b110111100100110;
		Coeff[10972] <= 15'b110111100100111;
		Coeff[10973] <= 15'b110111100101001;
		Coeff[10974] <= 15'b110111100101010;
		Coeff[10975] <= 15'b110111100101100;
		Coeff[10976] <= 15'b110111100101101;
		Coeff[10977] <= 15'b110111100101111;
		Coeff[10978] <= 15'b110111100110000;
		Coeff[10979] <= 15'b110111100110010;
		Coeff[10980] <= 15'b110111100110100;
		Coeff[10981] <= 15'b110111100110101;
		Coeff[10982] <= 15'b110111100110111;
		Coeff[10983] <= 15'b110111100111000;
		Coeff[10984] <= 15'b110111100111010;
		Coeff[10985] <= 15'b110111100111011;
		Coeff[10986] <= 15'b110111100111101;
		Coeff[10987] <= 15'b110111100111110;
		Coeff[10988] <= 15'b110111101000000;
		Coeff[10989] <= 15'b110111101000010;
		Coeff[10990] <= 15'b110111101000011;
		Coeff[10991] <= 15'b110111101000101;
		Coeff[10992] <= 15'b110111101000110;
		Coeff[10993] <= 15'b110111101001000;
		Coeff[10994] <= 15'b110111101001001;
		Coeff[10995] <= 15'b110111101001011;
		Coeff[10996] <= 15'b110111101001100;
		Coeff[10997] <= 15'b110111101001110;
		Coeff[10998] <= 15'b110111101010000;
		Coeff[10999] <= 15'b110111101010001;
		Coeff[11000] <= 15'b110111101010011;
		Coeff[11001] <= 15'b110111101010100;
		Coeff[11002] <= 15'b110111101010110;
		Coeff[11003] <= 15'b110111101010111;
		Coeff[11004] <= 15'b110111101011001;
		Coeff[11005] <= 15'b110111101011010;
		Coeff[11006] <= 15'b110111101011100;
		Coeff[11007] <= 15'b110111101011101;
		Coeff[11008] <= 15'b110111101011111;
		Coeff[11009] <= 15'b110111101100001;
		Coeff[11010] <= 15'b110111101100010;
		Coeff[11011] <= 15'b110111101100100;
		Coeff[11012] <= 15'b110111101100101;
		Coeff[11013] <= 15'b110111101100111;
		Coeff[11014] <= 15'b110111101101000;
		Coeff[11015] <= 15'b110111101101010;
		Coeff[11016] <= 15'b110111101101011;
		Coeff[11017] <= 15'b110111101101101;
		Coeff[11018] <= 15'b110111101101110;
		Coeff[11019] <= 15'b110111101110000;
		Coeff[11020] <= 15'b110111101110010;
		Coeff[11021] <= 15'b110111101110011;
		Coeff[11022] <= 15'b110111101110101;
		Coeff[11023] <= 15'b110111101110110;
		Coeff[11024] <= 15'b110111101111000;
		Coeff[11025] <= 15'b110111101111001;
		Coeff[11026] <= 15'b110111101111011;
		Coeff[11027] <= 15'b110111101111100;
		Coeff[11028] <= 15'b110111101111110;
		Coeff[11029] <= 15'b110111101111111;
		Coeff[11030] <= 15'b110111110000001;
		Coeff[11031] <= 15'b110111110000011;
		Coeff[11032] <= 15'b110111110000100;
		Coeff[11033] <= 15'b110111110000110;
		Coeff[11034] <= 15'b110111110000111;
		Coeff[11035] <= 15'b110111110001001;
		Coeff[11036] <= 15'b110111110001010;
		Coeff[11037] <= 15'b110111110001100;
		Coeff[11038] <= 15'b110111110001101;
		Coeff[11039] <= 15'b110111110001111;
		Coeff[11040] <= 15'b110111110010000;
		Coeff[11041] <= 15'b110111110010010;
		Coeff[11042] <= 15'b110111110010100;
		Coeff[11043] <= 15'b110111110010101;
		Coeff[11044] <= 15'b110111110010111;
		Coeff[11045] <= 15'b110111110011000;
		Coeff[11046] <= 15'b110111110011010;
		Coeff[11047] <= 15'b110111110011011;
		Coeff[11048] <= 15'b110111110011101;
		Coeff[11049] <= 15'b110111110011110;
		Coeff[11050] <= 15'b110111110100000;
		Coeff[11051] <= 15'b110111110100001;
		Coeff[11052] <= 15'b110111110100011;
		Coeff[11053] <= 15'b110111110100100;
		Coeff[11054] <= 15'b110111110100110;
		Coeff[11055] <= 15'b110111110100111;
		Coeff[11056] <= 15'b110111110101001;
		Coeff[11057] <= 15'b110111110101011;
		Coeff[11058] <= 15'b110111110101100;
		Coeff[11059] <= 15'b110111110101110;
		Coeff[11060] <= 15'b110111110101111;
		Coeff[11061] <= 15'b110111110110001;
		Coeff[11062] <= 15'b110111110110010;
		Coeff[11063] <= 15'b110111110110100;
		Coeff[11064] <= 15'b110111110110101;
		Coeff[11065] <= 15'b110111110110111;
		Coeff[11066] <= 15'b110111110111000;
		Coeff[11067] <= 15'b110111110111010;
		Coeff[11068] <= 15'b110111110111011;
		Coeff[11069] <= 15'b110111110111101;
		Coeff[11070] <= 15'b110111110111111;
		Coeff[11071] <= 15'b110111111000000;
		Coeff[11072] <= 15'b110111111000010;
		Coeff[11073] <= 15'b110111111000011;
		Coeff[11074] <= 15'b110111111000101;
		Coeff[11075] <= 15'b110111111000110;
		Coeff[11076] <= 15'b110111111001000;
		Coeff[11077] <= 15'b110111111001001;
		Coeff[11078] <= 15'b110111111001011;
		Coeff[11079] <= 15'b110111111001100;
		Coeff[11080] <= 15'b110111111001110;
		Coeff[11081] <= 15'b110111111001111;
		Coeff[11082] <= 15'b110111111010001;
		Coeff[11083] <= 15'b110111111010010;
		Coeff[11084] <= 15'b110111111010100;
		Coeff[11085] <= 15'b110111111010101;
		Coeff[11086] <= 15'b110111111010111;
		Coeff[11087] <= 15'b110111111011001;
		Coeff[11088] <= 15'b110111111011010;
		Coeff[11089] <= 15'b110111111011100;
		Coeff[11090] <= 15'b110111111011101;
		Coeff[11091] <= 15'b110111111011111;
		Coeff[11092] <= 15'b110111111100000;
		Coeff[11093] <= 15'b110111111100010;
		Coeff[11094] <= 15'b110111111100011;
		Coeff[11095] <= 15'b110111111100101;
		Coeff[11096] <= 15'b110111111100110;
		Coeff[11097] <= 15'b110111111101000;
		Coeff[11098] <= 15'b110111111101001;
		Coeff[11099] <= 15'b110111111101011;
		Coeff[11100] <= 15'b110111111101100;
		Coeff[11101] <= 15'b110111111101110;
		Coeff[11102] <= 15'b110111111101111;
		Coeff[11103] <= 15'b110111111110001;
		Coeff[11104] <= 15'b110111111110010;
		Coeff[11105] <= 15'b110111111110100;
		Coeff[11106] <= 15'b110111111110110;
		Coeff[11107] <= 15'b110111111110111;
		Coeff[11108] <= 15'b110111111111001;
		Coeff[11109] <= 15'b110111111111010;
		Coeff[11110] <= 15'b110111111111100;
		Coeff[11111] <= 15'b110111111111101;
		Coeff[11112] <= 15'b110111111111111;
		Coeff[11113] <= 15'b111000000000000;
		Coeff[11114] <= 15'b111000000000010;
		Coeff[11115] <= 15'b111000000000011;
		Coeff[11116] <= 15'b111000000000101;
		Coeff[11117] <= 15'b111000000000110;
		Coeff[11118] <= 15'b111000000001000;
		Coeff[11119] <= 15'b111000000001001;
		Coeff[11120] <= 15'b111000000001011;
		Coeff[11121] <= 15'b111000000001100;
		Coeff[11122] <= 15'b111000000001110;
		Coeff[11123] <= 15'b111000000001111;
		Coeff[11124] <= 15'b111000000010001;
		Coeff[11125] <= 15'b111000000010010;
		Coeff[11126] <= 15'b111000000010100;
		Coeff[11127] <= 15'b111000000010101;
		Coeff[11128] <= 15'b111000000010111;
		Coeff[11129] <= 15'b111000000011000;
		Coeff[11130] <= 15'b111000000011010;
		Coeff[11131] <= 15'b111000000011011;
		Coeff[11132] <= 15'b111000000011101;
		Coeff[11133] <= 15'b111000000011111;
		Coeff[11134] <= 15'b111000000100000;
		Coeff[11135] <= 15'b111000000100010;
		Coeff[11136] <= 15'b111000000100011;
		Coeff[11137] <= 15'b111000000100101;
		Coeff[11138] <= 15'b111000000100110;
		Coeff[11139] <= 15'b111000000101000;
		Coeff[11140] <= 15'b111000000101001;
		Coeff[11141] <= 15'b111000000101011;
		Coeff[11142] <= 15'b111000000101100;
		Coeff[11143] <= 15'b111000000101110;
		Coeff[11144] <= 15'b111000000101111;
		Coeff[11145] <= 15'b111000000110001;
		Coeff[11146] <= 15'b111000000110010;
		Coeff[11147] <= 15'b111000000110100;
		Coeff[11148] <= 15'b111000000110101;
		Coeff[11149] <= 15'b111000000110111;
		Coeff[11150] <= 15'b111000000111000;
		Coeff[11151] <= 15'b111000000111010;
		Coeff[11152] <= 15'b111000000111011;
		Coeff[11153] <= 15'b111000000111101;
		Coeff[11154] <= 15'b111000000111110;
		Coeff[11155] <= 15'b111000001000000;
		Coeff[11156] <= 15'b111000001000001;
		Coeff[11157] <= 15'b111000001000011;
		Coeff[11158] <= 15'b111000001000100;
		Coeff[11159] <= 15'b111000001000110;
		Coeff[11160] <= 15'b111000001000111;
		Coeff[11161] <= 15'b111000001001001;
		Coeff[11162] <= 15'b111000001001010;
		Coeff[11163] <= 15'b111000001001100;
		Coeff[11164] <= 15'b111000001001101;
		Coeff[11165] <= 15'b111000001001111;
		Coeff[11166] <= 15'b111000001010000;
		Coeff[11167] <= 15'b111000001010010;
		Coeff[11168] <= 15'b111000001010011;
		Coeff[11169] <= 15'b111000001010101;
		Coeff[11170] <= 15'b111000001010110;
		Coeff[11171] <= 15'b111000001011000;
		Coeff[11172] <= 15'b111000001011001;
		Coeff[11173] <= 15'b111000001011011;
		Coeff[11174] <= 15'b111000001011100;
		Coeff[11175] <= 15'b111000001011110;
		Coeff[11176] <= 15'b111000001011111;
		Coeff[11177] <= 15'b111000001100001;
		Coeff[11178] <= 15'b111000001100010;
		Coeff[11179] <= 15'b111000001100100;
		Coeff[11180] <= 15'b111000001100101;
		Coeff[11181] <= 15'b111000001100111;
		Coeff[11182] <= 15'b111000001101000;
		Coeff[11183] <= 15'b111000001101010;
		Coeff[11184] <= 15'b111000001101011;
		Coeff[11185] <= 15'b111000001101101;
		Coeff[11186] <= 15'b111000001101110;
		Coeff[11187] <= 15'b111000001110000;
		Coeff[11188] <= 15'b111000001110001;
		Coeff[11189] <= 15'b111000001110011;
		Coeff[11190] <= 15'b111000001110100;
		Coeff[11191] <= 15'b111000001110110;
		Coeff[11192] <= 15'b111000001110111;
		Coeff[11193] <= 15'b111000001111001;
		Coeff[11194] <= 15'b111000001111010;
		Coeff[11195] <= 15'b111000001111100;
		Coeff[11196] <= 15'b111000001111101;
		Coeff[11197] <= 15'b111000001111111;
		Coeff[11198] <= 15'b111000010000000;
		Coeff[11199] <= 15'b111000010000010;
		Coeff[11200] <= 15'b111000010000011;
		Coeff[11201] <= 15'b111000010000101;
		Coeff[11202] <= 15'b111000010000110;
		Coeff[11203] <= 15'b111000010001000;
		Coeff[11204] <= 15'b111000010001001;
		Coeff[11205] <= 15'b111000010001011;
		Coeff[11206] <= 15'b111000010001100;
		Coeff[11207] <= 15'b111000010001110;
		Coeff[11208] <= 15'b111000010001111;
		Coeff[11209] <= 15'b111000010010001;
		Coeff[11210] <= 15'b111000010010010;
		Coeff[11211] <= 15'b111000010010100;
		Coeff[11212] <= 15'b111000010010101;
		Coeff[11213] <= 15'b111000010010111;
		Coeff[11214] <= 15'b111000010011000;
		Coeff[11215] <= 15'b111000010011010;
		Coeff[11216] <= 15'b111000010011011;
		Coeff[11217] <= 15'b111000010011101;
		Coeff[11218] <= 15'b111000010011110;
		Coeff[11219] <= 15'b111000010100000;
		Coeff[11220] <= 15'b111000010100001;
		Coeff[11221] <= 15'b111000010100011;
		Coeff[11222] <= 15'b111000010100100;
		Coeff[11223] <= 15'b111000010100110;
		Coeff[11224] <= 15'b111000010100111;
		Coeff[11225] <= 15'b111000010101001;
		Coeff[11226] <= 15'b111000010101010;
		Coeff[11227] <= 15'b111000010101100;
		Coeff[11228] <= 15'b111000010101101;
		Coeff[11229] <= 15'b111000010101111;
		Coeff[11230] <= 15'b111000010110000;
		Coeff[11231] <= 15'b111000010110010;
		Coeff[11232] <= 15'b111000010110011;
		Coeff[11233] <= 15'b111000010110101;
		Coeff[11234] <= 15'b111000010110110;
		Coeff[11235] <= 15'b111000010111000;
		Coeff[11236] <= 15'b111000010111001;
		Coeff[11237] <= 15'b111000010111011;
		Coeff[11238] <= 15'b111000010111100;
		Coeff[11239] <= 15'b111000010111110;
		Coeff[11240] <= 15'b111000010111111;
		Coeff[11241] <= 15'b111000011000001;
		Coeff[11242] <= 15'b111000011000010;
		Coeff[11243] <= 15'b111000011000100;
		Coeff[11244] <= 15'b111000011000101;
		Coeff[11245] <= 15'b111000011000111;
		Coeff[11246] <= 15'b111000011001000;
		Coeff[11247] <= 15'b111000011001010;
		Coeff[11248] <= 15'b111000011001011;
		Coeff[11249] <= 15'b111000011001101;
		Coeff[11250] <= 15'b111000011001110;
		Coeff[11251] <= 15'b111000011010000;
		Coeff[11252] <= 15'b111000011010001;
		Coeff[11253] <= 15'b111000011010010;
		Coeff[11254] <= 15'b111000011010100;
		Coeff[11255] <= 15'b111000011010101;
		Coeff[11256] <= 15'b111000011010111;
		Coeff[11257] <= 15'b111000011011000;
		Coeff[11258] <= 15'b111000011011010;
		Coeff[11259] <= 15'b111000011011011;
		Coeff[11260] <= 15'b111000011011101;
		Coeff[11261] <= 15'b111000011011110;
		Coeff[11262] <= 15'b111000011100000;
		Coeff[11263] <= 15'b111000011100001;
		Coeff[11264] <= 15'b111000011100011;
		Coeff[11265] <= 15'b111000011100100;
		Coeff[11266] <= 15'b111000011100110;
		Coeff[11267] <= 15'b111000011100111;
		Coeff[11268] <= 15'b111000011101001;
		Coeff[11269] <= 15'b111000011101010;
		Coeff[11270] <= 15'b111000011101100;
		Coeff[11271] <= 15'b111000011101101;
		Coeff[11272] <= 15'b111000011101111;
		Coeff[11273] <= 15'b111000011110000;
		Coeff[11274] <= 15'b111000011110010;
		Coeff[11275] <= 15'b111000011110011;
		Coeff[11276] <= 15'b111000011110101;
		Coeff[11277] <= 15'b111000011110110;
		Coeff[11278] <= 15'b111000011111000;
		Coeff[11279] <= 15'b111000011111001;
		Coeff[11280] <= 15'b111000011111010;
		Coeff[11281] <= 15'b111000011111100;
		Coeff[11282] <= 15'b111000011111101;
		Coeff[11283] <= 15'b111000011111111;
		Coeff[11284] <= 15'b111000100000000;
		Coeff[11285] <= 15'b111000100000010;
		Coeff[11286] <= 15'b111000100000011;
		Coeff[11287] <= 15'b111000100000101;
		Coeff[11288] <= 15'b111000100000110;
		Coeff[11289] <= 15'b111000100001000;
		Coeff[11290] <= 15'b111000100001001;
		Coeff[11291] <= 15'b111000100001011;
		Coeff[11292] <= 15'b111000100001100;
		Coeff[11293] <= 15'b111000100001110;
		Coeff[11294] <= 15'b111000100001111;
		Coeff[11295] <= 15'b111000100010001;
		Coeff[11296] <= 15'b111000100010010;
		Coeff[11297] <= 15'b111000100010100;
		Coeff[11298] <= 15'b111000100010101;
		Coeff[11299] <= 15'b111000100010110;
		Coeff[11300] <= 15'b111000100011000;
		Coeff[11301] <= 15'b111000100011001;
		Coeff[11302] <= 15'b111000100011011;
		Coeff[11303] <= 15'b111000100011100;
		Coeff[11304] <= 15'b111000100011110;
		Coeff[11305] <= 15'b111000100011111;
		Coeff[11306] <= 15'b111000100100001;
		Coeff[11307] <= 15'b111000100100010;
		Coeff[11308] <= 15'b111000100100100;
		Coeff[11309] <= 15'b111000100100101;
		Coeff[11310] <= 15'b111000100100111;
		Coeff[11311] <= 15'b111000100101000;
		Coeff[11312] <= 15'b111000100101010;
		Coeff[11313] <= 15'b111000100101011;
		Coeff[11314] <= 15'b111000100101101;
		Coeff[11315] <= 15'b111000100101110;
		Coeff[11316] <= 15'b111000100101111;
		Coeff[11317] <= 15'b111000100110001;
		Coeff[11318] <= 15'b111000100110010;
		Coeff[11319] <= 15'b111000100110100;
		Coeff[11320] <= 15'b111000100110101;
		Coeff[11321] <= 15'b111000100110111;
		Coeff[11322] <= 15'b111000100111000;
		Coeff[11323] <= 15'b111000100111010;
		Coeff[11324] <= 15'b111000100111011;
		Coeff[11325] <= 15'b111000100111101;
		Coeff[11326] <= 15'b111000100111110;
		Coeff[11327] <= 15'b111000101000000;
		Coeff[11328] <= 15'b111000101000001;
		Coeff[11329] <= 15'b111000101000010;
		Coeff[11330] <= 15'b111000101000100;
		Coeff[11331] <= 15'b111000101000101;
		Coeff[11332] <= 15'b111000101000111;
		Coeff[11333] <= 15'b111000101001000;
		Coeff[11334] <= 15'b111000101001010;
		Coeff[11335] <= 15'b111000101001011;
		Coeff[11336] <= 15'b111000101001101;
		Coeff[11337] <= 15'b111000101001110;
		Coeff[11338] <= 15'b111000101010000;
		Coeff[11339] <= 15'b111000101010001;
		Coeff[11340] <= 15'b111000101010011;
		Coeff[11341] <= 15'b111000101010100;
		Coeff[11342] <= 15'b111000101010101;
		Coeff[11343] <= 15'b111000101010111;
		Coeff[11344] <= 15'b111000101011000;
		Coeff[11345] <= 15'b111000101011010;
		Coeff[11346] <= 15'b111000101011011;
		Coeff[11347] <= 15'b111000101011101;
		Coeff[11348] <= 15'b111000101011110;
		Coeff[11349] <= 15'b111000101100000;
		Coeff[11350] <= 15'b111000101100001;
		Coeff[11351] <= 15'b111000101100011;
		Coeff[11352] <= 15'b111000101100100;
		Coeff[11353] <= 15'b111000101100110;
		Coeff[11354] <= 15'b111000101100111;
		Coeff[11355] <= 15'b111000101101000;
		Coeff[11356] <= 15'b111000101101010;
		Coeff[11357] <= 15'b111000101101011;
		Coeff[11358] <= 15'b111000101101101;
		Coeff[11359] <= 15'b111000101101110;
		Coeff[11360] <= 15'b111000101110000;
		Coeff[11361] <= 15'b111000101110001;
		Coeff[11362] <= 15'b111000101110011;
		Coeff[11363] <= 15'b111000101110100;
		Coeff[11364] <= 15'b111000101110110;
		Coeff[11365] <= 15'b111000101110111;
		Coeff[11366] <= 15'b111000101111000;
		Coeff[11367] <= 15'b111000101111010;
		Coeff[11368] <= 15'b111000101111011;
		Coeff[11369] <= 15'b111000101111101;
		Coeff[11370] <= 15'b111000101111110;
		Coeff[11371] <= 15'b111000110000000;
		Coeff[11372] <= 15'b111000110000001;
		Coeff[11373] <= 15'b111000110000011;
		Coeff[11374] <= 15'b111000110000100;
		Coeff[11375] <= 15'b111000110000110;
		Coeff[11376] <= 15'b111000110000111;
		Coeff[11377] <= 15'b111000110001000;
		Coeff[11378] <= 15'b111000110001010;
		Coeff[11379] <= 15'b111000110001011;
		Coeff[11380] <= 15'b111000110001101;
		Coeff[11381] <= 15'b111000110001110;
		Coeff[11382] <= 15'b111000110010000;
		Coeff[11383] <= 15'b111000110010001;
		Coeff[11384] <= 15'b111000110010011;
		Coeff[11385] <= 15'b111000110010100;
		Coeff[11386] <= 15'b111000110010101;
		Coeff[11387] <= 15'b111000110010111;
		Coeff[11388] <= 15'b111000110011000;
		Coeff[11389] <= 15'b111000110011010;
		Coeff[11390] <= 15'b111000110011011;
		Coeff[11391] <= 15'b111000110011101;
		Coeff[11392] <= 15'b111000110011110;
		Coeff[11393] <= 15'b111000110100000;
		Coeff[11394] <= 15'b111000110100001;
		Coeff[11395] <= 15'b111000110100011;
		Coeff[11396] <= 15'b111000110100100;
		Coeff[11397] <= 15'b111000110100101;
		Coeff[11398] <= 15'b111000110100111;
		Coeff[11399] <= 15'b111000110101000;
		Coeff[11400] <= 15'b111000110101010;
		Coeff[11401] <= 15'b111000110101011;
		Coeff[11402] <= 15'b111000110101101;
		Coeff[11403] <= 15'b111000110101110;
		Coeff[11404] <= 15'b111000110110000;
		Coeff[11405] <= 15'b111000110110001;
		Coeff[11406] <= 15'b111000110110010;
		Coeff[11407] <= 15'b111000110110100;
		Coeff[11408] <= 15'b111000110110101;
		Coeff[11409] <= 15'b111000110110111;
		Coeff[11410] <= 15'b111000110111000;
		Coeff[11411] <= 15'b111000110111010;
		Coeff[11412] <= 15'b111000110111011;
		Coeff[11413] <= 15'b111000110111100;
		Coeff[11414] <= 15'b111000110111110;
		Coeff[11415] <= 15'b111000110111111;
		Coeff[11416] <= 15'b111000111000001;
		Coeff[11417] <= 15'b111000111000010;
		Coeff[11418] <= 15'b111000111000100;
		Coeff[11419] <= 15'b111000111000101;
		Coeff[11420] <= 15'b111000111000111;
		Coeff[11421] <= 15'b111000111001000;
		Coeff[11422] <= 15'b111000111001001;
		Coeff[11423] <= 15'b111000111001011;
		Coeff[11424] <= 15'b111000111001100;
		Coeff[11425] <= 15'b111000111001110;
		Coeff[11426] <= 15'b111000111001111;
		Coeff[11427] <= 15'b111000111010001;
		Coeff[11428] <= 15'b111000111010010;
		Coeff[11429] <= 15'b111000111010100;
		Coeff[11430] <= 15'b111000111010101;
		Coeff[11431] <= 15'b111000111010110;
		Coeff[11432] <= 15'b111000111011000;
		Coeff[11433] <= 15'b111000111011001;
		Coeff[11434] <= 15'b111000111011011;
		Coeff[11435] <= 15'b111000111011100;
		Coeff[11436] <= 15'b111000111011110;
		Coeff[11437] <= 15'b111000111011111;
		Coeff[11438] <= 15'b111000111100000;
		Coeff[11439] <= 15'b111000111100010;
		Coeff[11440] <= 15'b111000111100011;
		Coeff[11441] <= 15'b111000111100101;
		Coeff[11442] <= 15'b111000111100110;
		Coeff[11443] <= 15'b111000111101000;
		Coeff[11444] <= 15'b111000111101001;
		Coeff[11445] <= 15'b111000111101010;
		Coeff[11446] <= 15'b111000111101100;
		Coeff[11447] <= 15'b111000111101101;
		Coeff[11448] <= 15'b111000111101111;
		Coeff[11449] <= 15'b111000111110000;
		Coeff[11450] <= 15'b111000111110010;
		Coeff[11451] <= 15'b111000111110011;
		Coeff[11452] <= 15'b111000111110101;
		Coeff[11453] <= 15'b111000111110110;
		Coeff[11454] <= 15'b111000111110111;
		Coeff[11455] <= 15'b111000111111001;
		Coeff[11456] <= 15'b111000111111010;
		Coeff[11457] <= 15'b111000111111100;
		Coeff[11458] <= 15'b111000111111101;
		Coeff[11459] <= 15'b111000111111111;
		Coeff[11460] <= 15'b111001000000000;
		Coeff[11461] <= 15'b111001000000001;
		Coeff[11462] <= 15'b111001000000011;
		Coeff[11463] <= 15'b111001000000100;
		Coeff[11464] <= 15'b111001000000110;
		Coeff[11465] <= 15'b111001000000111;
		Coeff[11466] <= 15'b111001000001001;
		Coeff[11467] <= 15'b111001000001010;
		Coeff[11468] <= 15'b111001000001011;
		Coeff[11469] <= 15'b111001000001101;
		Coeff[11470] <= 15'b111001000001110;
		Coeff[11471] <= 15'b111001000010000;
		Coeff[11472] <= 15'b111001000010001;
		Coeff[11473] <= 15'b111001000010010;
		Coeff[11474] <= 15'b111001000010100;
		Coeff[11475] <= 15'b111001000010101;
		Coeff[11476] <= 15'b111001000010111;
		Coeff[11477] <= 15'b111001000011000;
		Coeff[11478] <= 15'b111001000011010;
		Coeff[11479] <= 15'b111001000011011;
		Coeff[11480] <= 15'b111001000011100;
		Coeff[11481] <= 15'b111001000011110;
		Coeff[11482] <= 15'b111001000011111;
		Coeff[11483] <= 15'b111001000100001;
		Coeff[11484] <= 15'b111001000100010;
		Coeff[11485] <= 15'b111001000100100;
		Coeff[11486] <= 15'b111001000100101;
		Coeff[11487] <= 15'b111001000100110;
		Coeff[11488] <= 15'b111001000101000;
		Coeff[11489] <= 15'b111001000101001;
		Coeff[11490] <= 15'b111001000101011;
		Coeff[11491] <= 15'b111001000101100;
		Coeff[11492] <= 15'b111001000101110;
		Coeff[11493] <= 15'b111001000101111;
		Coeff[11494] <= 15'b111001000110000;
		Coeff[11495] <= 15'b111001000110010;
		Coeff[11496] <= 15'b111001000110011;
		Coeff[11497] <= 15'b111001000110101;
		Coeff[11498] <= 15'b111001000110110;
		Coeff[11499] <= 15'b111001000110111;
		Coeff[11500] <= 15'b111001000111001;
		Coeff[11501] <= 15'b111001000111010;
		Coeff[11502] <= 15'b111001000111100;
		Coeff[11503] <= 15'b111001000111101;
		Coeff[11504] <= 15'b111001000111111;
		Coeff[11505] <= 15'b111001001000000;
		Coeff[11506] <= 15'b111001001000001;
		Coeff[11507] <= 15'b111001001000011;
		Coeff[11508] <= 15'b111001001000100;
		Coeff[11509] <= 15'b111001001000110;
		Coeff[11510] <= 15'b111001001000111;
		Coeff[11511] <= 15'b111001001001000;
		Coeff[11512] <= 15'b111001001001010;
		Coeff[11513] <= 15'b111001001001011;
		Coeff[11514] <= 15'b111001001001101;
		Coeff[11515] <= 15'b111001001001110;
		Coeff[11516] <= 15'b111001001010000;
		Coeff[11517] <= 15'b111001001010001;
		Coeff[11518] <= 15'b111001001010010;
		Coeff[11519] <= 15'b111001001010100;
		Coeff[11520] <= 15'b111001001010101;
		Coeff[11521] <= 15'b111001001010111;
		Coeff[11522] <= 15'b111001001011000;
		Coeff[11523] <= 15'b111001001011001;
		Coeff[11524] <= 15'b111001001011011;
		Coeff[11525] <= 15'b111001001011100;
		Coeff[11526] <= 15'b111001001011110;
		Coeff[11527] <= 15'b111001001011111;
		Coeff[11528] <= 15'b111001001100000;
		Coeff[11529] <= 15'b111001001100010;
		Coeff[11530] <= 15'b111001001100011;
		Coeff[11531] <= 15'b111001001100101;
		Coeff[11532] <= 15'b111001001100110;
		Coeff[11533] <= 15'b111001001101000;
		Coeff[11534] <= 15'b111001001101001;
		Coeff[11535] <= 15'b111001001101010;
		Coeff[11536] <= 15'b111001001101100;
		Coeff[11537] <= 15'b111001001101101;
		Coeff[11538] <= 15'b111001001101111;
		Coeff[11539] <= 15'b111001001110000;
		Coeff[11540] <= 15'b111001001110001;
		Coeff[11541] <= 15'b111001001110011;
		Coeff[11542] <= 15'b111001001110100;
		Coeff[11543] <= 15'b111001001110110;
		Coeff[11544] <= 15'b111001001110111;
		Coeff[11545] <= 15'b111001001111000;
		Coeff[11546] <= 15'b111001001111010;
		Coeff[11547] <= 15'b111001001111011;
		Coeff[11548] <= 15'b111001001111101;
		Coeff[11549] <= 15'b111001001111110;
		Coeff[11550] <= 15'b111001001111111;
		Coeff[11551] <= 15'b111001010000001;
		Coeff[11552] <= 15'b111001010000010;
		Coeff[11553] <= 15'b111001010000100;
		Coeff[11554] <= 15'b111001010000101;
		Coeff[11555] <= 15'b111001010000110;
		Coeff[11556] <= 15'b111001010001000;
		Coeff[11557] <= 15'b111001010001001;
		Coeff[11558] <= 15'b111001010001011;
		Coeff[11559] <= 15'b111001010001100;
		Coeff[11560] <= 15'b111001010001101;
		Coeff[11561] <= 15'b111001010001111;
		Coeff[11562] <= 15'b111001010010000;
		Coeff[11563] <= 15'b111001010010010;
		Coeff[11564] <= 15'b111001010010011;
		Coeff[11565] <= 15'b111001010010100;
		Coeff[11566] <= 15'b111001010010110;
		Coeff[11567] <= 15'b111001010010111;
		Coeff[11568] <= 15'b111001010011001;
		Coeff[11569] <= 15'b111001010011010;
		Coeff[11570] <= 15'b111001010011011;
		Coeff[11571] <= 15'b111001010011101;
		Coeff[11572] <= 15'b111001010011110;
		Coeff[11573] <= 15'b111001010100000;
		Coeff[11574] <= 15'b111001010100001;
		Coeff[11575] <= 15'b111001010100010;
		Coeff[11576] <= 15'b111001010100100;
		Coeff[11577] <= 15'b111001010100101;
		Coeff[11578] <= 15'b111001010100111;
		Coeff[11579] <= 15'b111001010101000;
		Coeff[11580] <= 15'b111001010101001;
		Coeff[11581] <= 15'b111001010101011;
		Coeff[11582] <= 15'b111001010101100;
		Coeff[11583] <= 15'b111001010101110;
		Coeff[11584] <= 15'b111001010101111;
		Coeff[11585] <= 15'b111001010110000;
		Coeff[11586] <= 15'b111001010110010;
		Coeff[11587] <= 15'b111001010110011;
		Coeff[11588] <= 15'b111001010110101;
		Coeff[11589] <= 15'b111001010110110;
		Coeff[11590] <= 15'b111001010110111;
		Coeff[11591] <= 15'b111001010111001;
		Coeff[11592] <= 15'b111001010111010;
		Coeff[11593] <= 15'b111001010111100;
		Coeff[11594] <= 15'b111001010111101;
		Coeff[11595] <= 15'b111001010111110;
		Coeff[11596] <= 15'b111001011000000;
		Coeff[11597] <= 15'b111001011000001;
		Coeff[11598] <= 15'b111001011000011;
		Coeff[11599] <= 15'b111001011000100;
		Coeff[11600] <= 15'b111001011000101;
		Coeff[11601] <= 15'b111001011000111;
		Coeff[11602] <= 15'b111001011001000;
		Coeff[11603] <= 15'b111001011001001;
		Coeff[11604] <= 15'b111001011001011;
		Coeff[11605] <= 15'b111001011001100;
		Coeff[11606] <= 15'b111001011001110;
		Coeff[11607] <= 15'b111001011001111;
		Coeff[11608] <= 15'b111001011010000;
		Coeff[11609] <= 15'b111001011010010;
		Coeff[11610] <= 15'b111001011010011;
		Coeff[11611] <= 15'b111001011010101;
		Coeff[11612] <= 15'b111001011010110;
		Coeff[11613] <= 15'b111001011010111;
		Coeff[11614] <= 15'b111001011011001;
		Coeff[11615] <= 15'b111001011011010;
		Coeff[11616] <= 15'b111001011011100;
		Coeff[11617] <= 15'b111001011011101;
		Coeff[11618] <= 15'b111001011011110;
		Coeff[11619] <= 15'b111001011100000;
		Coeff[11620] <= 15'b111001011100001;
		Coeff[11621] <= 15'b111001011100010;
		Coeff[11622] <= 15'b111001011100100;
		Coeff[11623] <= 15'b111001011100101;
		Coeff[11624] <= 15'b111001011100111;
		Coeff[11625] <= 15'b111001011101000;
		Coeff[11626] <= 15'b111001011101001;
		Coeff[11627] <= 15'b111001011101011;
		Coeff[11628] <= 15'b111001011101100;
		Coeff[11629] <= 15'b111001011101110;
		Coeff[11630] <= 15'b111001011101111;
		Coeff[11631] <= 15'b111001011110000;
		Coeff[11632] <= 15'b111001011110010;
		Coeff[11633] <= 15'b111001011110011;
		Coeff[11634] <= 15'b111001011110100;
		Coeff[11635] <= 15'b111001011110110;
		Coeff[11636] <= 15'b111001011110111;
		Coeff[11637] <= 15'b111001011111001;
		Coeff[11638] <= 15'b111001011111010;
		Coeff[11639] <= 15'b111001011111011;
		Coeff[11640] <= 15'b111001011111101;
		Coeff[11641] <= 15'b111001011111110;
		Coeff[11642] <= 15'b111001011111111;
		Coeff[11643] <= 15'b111001100000001;
		Coeff[11644] <= 15'b111001100000010;
		Coeff[11645] <= 15'b111001100000100;
		Coeff[11646] <= 15'b111001100000101;
		Coeff[11647] <= 15'b111001100000110;
		Coeff[11648] <= 15'b111001100001000;
		Coeff[11649] <= 15'b111001100001001;
		Coeff[11650] <= 15'b111001100001011;
		Coeff[11651] <= 15'b111001100001100;
		Coeff[11652] <= 15'b111001100001101;
		Coeff[11653] <= 15'b111001100001111;
		Coeff[11654] <= 15'b111001100010000;
		Coeff[11655] <= 15'b111001100010001;
		Coeff[11656] <= 15'b111001100010011;
		Coeff[11657] <= 15'b111001100010100;
		Coeff[11658] <= 15'b111001100010110;
		Coeff[11659] <= 15'b111001100010111;
		Coeff[11660] <= 15'b111001100011000;
		Coeff[11661] <= 15'b111001100011010;
		Coeff[11662] <= 15'b111001100011011;
		Coeff[11663] <= 15'b111001100011100;
		Coeff[11664] <= 15'b111001100011110;
		Coeff[11665] <= 15'b111001100011111;
		Coeff[11666] <= 15'b111001100100001;
		Coeff[11667] <= 15'b111001100100010;
		Coeff[11668] <= 15'b111001100100011;
		Coeff[11669] <= 15'b111001100100101;
		Coeff[11670] <= 15'b111001100100110;
		Coeff[11671] <= 15'b111001100100111;
		Coeff[11672] <= 15'b111001100101001;
		Coeff[11673] <= 15'b111001100101010;
		Coeff[11674] <= 15'b111001100101100;
		Coeff[11675] <= 15'b111001100101101;
		Coeff[11676] <= 15'b111001100101110;
		Coeff[11677] <= 15'b111001100110000;
		Coeff[11678] <= 15'b111001100110001;
		Coeff[11679] <= 15'b111001100110010;
		Coeff[11680] <= 15'b111001100110100;
		Coeff[11681] <= 15'b111001100110101;
		Coeff[11682] <= 15'b111001100110110;
		Coeff[11683] <= 15'b111001100111000;
		Coeff[11684] <= 15'b111001100111001;
		Coeff[11685] <= 15'b111001100111011;
		Coeff[11686] <= 15'b111001100111100;
		Coeff[11687] <= 15'b111001100111101;
		Coeff[11688] <= 15'b111001100111111;
		Coeff[11689] <= 15'b111001101000000;
		Coeff[11690] <= 15'b111001101000001;
		Coeff[11691] <= 15'b111001101000011;
		Coeff[11692] <= 15'b111001101000100;
		Coeff[11693] <= 15'b111001101000101;
		Coeff[11694] <= 15'b111001101000111;
		Coeff[11695] <= 15'b111001101001000;
		Coeff[11696] <= 15'b111001101001010;
		Coeff[11697] <= 15'b111001101001011;
		Coeff[11698] <= 15'b111001101001100;
		Coeff[11699] <= 15'b111001101001110;
		Coeff[11700] <= 15'b111001101001111;
		Coeff[11701] <= 15'b111001101010000;
		Coeff[11702] <= 15'b111001101010010;
		Coeff[11703] <= 15'b111001101010011;
		Coeff[11704] <= 15'b111001101010101;
		Coeff[11705] <= 15'b111001101010110;
		Coeff[11706] <= 15'b111001101010111;
		Coeff[11707] <= 15'b111001101011001;
		Coeff[11708] <= 15'b111001101011010;
		Coeff[11709] <= 15'b111001101011011;
		Coeff[11710] <= 15'b111001101011101;
		Coeff[11711] <= 15'b111001101011110;
		Coeff[11712] <= 15'b111001101011111;
		Coeff[11713] <= 15'b111001101100001;
		Coeff[11714] <= 15'b111001101100010;
		Coeff[11715] <= 15'b111001101100011;
		Coeff[11716] <= 15'b111001101100101;
		Coeff[11717] <= 15'b111001101100110;
		Coeff[11718] <= 15'b111001101101000;
		Coeff[11719] <= 15'b111001101101001;
		Coeff[11720] <= 15'b111001101101010;
		Coeff[11721] <= 15'b111001101101100;
		Coeff[11722] <= 15'b111001101101101;
		Coeff[11723] <= 15'b111001101101110;
		Coeff[11724] <= 15'b111001101110000;
		Coeff[11725] <= 15'b111001101110001;
		Coeff[11726] <= 15'b111001101110010;
		Coeff[11727] <= 15'b111001101110100;
		Coeff[11728] <= 15'b111001101110101;
		Coeff[11729] <= 15'b111001101110110;
		Coeff[11730] <= 15'b111001101111000;
		Coeff[11731] <= 15'b111001101111001;
		Coeff[11732] <= 15'b111001101111011;
		Coeff[11733] <= 15'b111001101111100;
		Coeff[11734] <= 15'b111001101111101;
		Coeff[11735] <= 15'b111001101111111;
		Coeff[11736] <= 15'b111001110000000;
		Coeff[11737] <= 15'b111001110000001;
		Coeff[11738] <= 15'b111001110000011;
		Coeff[11739] <= 15'b111001110000100;
		Coeff[11740] <= 15'b111001110000101;
		Coeff[11741] <= 15'b111001110000111;
		Coeff[11742] <= 15'b111001110001000;
		Coeff[11743] <= 15'b111001110001001;
		Coeff[11744] <= 15'b111001110001011;
		Coeff[11745] <= 15'b111001110001100;
		Coeff[11746] <= 15'b111001110001110;
		Coeff[11747] <= 15'b111001110001111;
		Coeff[11748] <= 15'b111001110010000;
		Coeff[11749] <= 15'b111001110010010;
		Coeff[11750] <= 15'b111001110010011;
		Coeff[11751] <= 15'b111001110010100;
		Coeff[11752] <= 15'b111001110010110;
		Coeff[11753] <= 15'b111001110010111;
		Coeff[11754] <= 15'b111001110011000;
		Coeff[11755] <= 15'b111001110011010;
		Coeff[11756] <= 15'b111001110011011;
		Coeff[11757] <= 15'b111001110011100;
		Coeff[11758] <= 15'b111001110011110;
		Coeff[11759] <= 15'b111001110011111;
		Coeff[11760] <= 15'b111001110100000;
		Coeff[11761] <= 15'b111001110100010;
		Coeff[11762] <= 15'b111001110100011;
		Coeff[11763] <= 15'b111001110100100;
		Coeff[11764] <= 15'b111001110100110;
		Coeff[11765] <= 15'b111001110100111;
		Coeff[11766] <= 15'b111001110101000;
		Coeff[11767] <= 15'b111001110101010;
		Coeff[11768] <= 15'b111001110101011;
		Coeff[11769] <= 15'b111001110101101;
		Coeff[11770] <= 15'b111001110101110;
		Coeff[11771] <= 15'b111001110101111;
		Coeff[11772] <= 15'b111001110110001;
		Coeff[11773] <= 15'b111001110110010;
		Coeff[11774] <= 15'b111001110110011;
		Coeff[11775] <= 15'b111001110110101;
		Coeff[11776] <= 15'b111001110110110;
		Coeff[11777] <= 15'b111001110110111;
		Coeff[11778] <= 15'b111001110111001;
		Coeff[11779] <= 15'b111001110111010;
		Coeff[11780] <= 15'b111001110111011;
		Coeff[11781] <= 15'b111001110111101;
		Coeff[11782] <= 15'b111001110111110;
		Coeff[11783] <= 15'b111001110111111;
		Coeff[11784] <= 15'b111001111000001;
		Coeff[11785] <= 15'b111001111000010;
		Coeff[11786] <= 15'b111001111000011;
		Coeff[11787] <= 15'b111001111000101;
		Coeff[11788] <= 15'b111001111000110;
		Coeff[11789] <= 15'b111001111000111;
		Coeff[11790] <= 15'b111001111001001;
		Coeff[11791] <= 15'b111001111001010;
		Coeff[11792] <= 15'b111001111001011;
		Coeff[11793] <= 15'b111001111001101;
		Coeff[11794] <= 15'b111001111001110;
		Coeff[11795] <= 15'b111001111001111;
		Coeff[11796] <= 15'b111001111010001;
		Coeff[11797] <= 15'b111001111010010;
		Coeff[11798] <= 15'b111001111010011;
		Coeff[11799] <= 15'b111001111010101;
		Coeff[11800] <= 15'b111001111010110;
		Coeff[11801] <= 15'b111001111010111;
		Coeff[11802] <= 15'b111001111011001;
		Coeff[11803] <= 15'b111001111011010;
		Coeff[11804] <= 15'b111001111011011;
		Coeff[11805] <= 15'b111001111011101;
		Coeff[11806] <= 15'b111001111011110;
		Coeff[11807] <= 15'b111001111011111;
		Coeff[11808] <= 15'b111001111100001;
		Coeff[11809] <= 15'b111001111100010;
		Coeff[11810] <= 15'b111001111100011;
		Coeff[11811] <= 15'b111001111100101;
		Coeff[11812] <= 15'b111001111100110;
		Coeff[11813] <= 15'b111001111100111;
		Coeff[11814] <= 15'b111001111101001;
		Coeff[11815] <= 15'b111001111101010;
		Coeff[11816] <= 15'b111001111101011;
		Coeff[11817] <= 15'b111001111101101;
		Coeff[11818] <= 15'b111001111101110;
		Coeff[11819] <= 15'b111001111101111;
		Coeff[11820] <= 15'b111001111110001;
		Coeff[11821] <= 15'b111001111110010;
		Coeff[11822] <= 15'b111001111110011;
		Coeff[11823] <= 15'b111001111110101;
		Coeff[11824] <= 15'b111001111110110;
		Coeff[11825] <= 15'b111001111110111;
		Coeff[11826] <= 15'b111001111111001;
		Coeff[11827] <= 15'b111001111111010;
		Coeff[11828] <= 15'b111001111111011;
		Coeff[11829] <= 15'b111001111111101;
		Coeff[11830] <= 15'b111001111111110;
		Coeff[11831] <= 15'b111001111111111;
		Coeff[11832] <= 15'b111010000000001;
		Coeff[11833] <= 15'b111010000000010;
		Coeff[11834] <= 15'b111010000000011;
		Coeff[11835] <= 15'b111010000000101;
		Coeff[11836] <= 15'b111010000000110;
		Coeff[11837] <= 15'b111010000000111;
		Coeff[11838] <= 15'b111010000001001;
		Coeff[11839] <= 15'b111010000001010;
		Coeff[11840] <= 15'b111010000001011;
		Coeff[11841] <= 15'b111010000001101;
		Coeff[11842] <= 15'b111010000001110;
		Coeff[11843] <= 15'b111010000001111;
		Coeff[11844] <= 15'b111010000010001;
		Coeff[11845] <= 15'b111010000010010;
		Coeff[11846] <= 15'b111010000010011;
		Coeff[11847] <= 15'b111010000010101;
		Coeff[11848] <= 15'b111010000010110;
		Coeff[11849] <= 15'b111010000010111;
		Coeff[11850] <= 15'b111010000011001;
		Coeff[11851] <= 15'b111010000011010;
		Coeff[11852] <= 15'b111010000011011;
		Coeff[11853] <= 15'b111010000011101;
		Coeff[11854] <= 15'b111010000011110;
		Coeff[11855] <= 15'b111010000011111;
		Coeff[11856] <= 15'b111010000100001;
		Coeff[11857] <= 15'b111010000100010;
		Coeff[11858] <= 15'b111010000100011;
		Coeff[11859] <= 15'b111010000100100;
		Coeff[11860] <= 15'b111010000100110;
		Coeff[11861] <= 15'b111010000100111;
		Coeff[11862] <= 15'b111010000101000;
		Coeff[11863] <= 15'b111010000101010;
		Coeff[11864] <= 15'b111010000101011;
		Coeff[11865] <= 15'b111010000101100;
		Coeff[11866] <= 15'b111010000101110;
		Coeff[11867] <= 15'b111010000101111;
		Coeff[11868] <= 15'b111010000110000;
		Coeff[11869] <= 15'b111010000110010;
		Coeff[11870] <= 15'b111010000110011;
		Coeff[11871] <= 15'b111010000110100;
		Coeff[11872] <= 15'b111010000110110;
		Coeff[11873] <= 15'b111010000110111;
		Coeff[11874] <= 15'b111010000111000;
		Coeff[11875] <= 15'b111010000111010;
		Coeff[11876] <= 15'b111010000111011;
		Coeff[11877] <= 15'b111010000111100;
		Coeff[11878] <= 15'b111010000111110;
		Coeff[11879] <= 15'b111010000111111;
		Coeff[11880] <= 15'b111010001000000;
		Coeff[11881] <= 15'b111010001000001;
		Coeff[11882] <= 15'b111010001000011;
		Coeff[11883] <= 15'b111010001000100;
		Coeff[11884] <= 15'b111010001000101;
		Coeff[11885] <= 15'b111010001000111;
		Coeff[11886] <= 15'b111010001001000;
		Coeff[11887] <= 15'b111010001001001;
		Coeff[11888] <= 15'b111010001001011;
		Coeff[11889] <= 15'b111010001001100;
		Coeff[11890] <= 15'b111010001001101;
		Coeff[11891] <= 15'b111010001001111;
		Coeff[11892] <= 15'b111010001010000;
		Coeff[11893] <= 15'b111010001010001;
		Coeff[11894] <= 15'b111010001010011;
		Coeff[11895] <= 15'b111010001010100;
		Coeff[11896] <= 15'b111010001010101;
		Coeff[11897] <= 15'b111010001010110;
		Coeff[11898] <= 15'b111010001011000;
		Coeff[11899] <= 15'b111010001011001;
		Coeff[11900] <= 15'b111010001011010;
		Coeff[11901] <= 15'b111010001011100;
		Coeff[11902] <= 15'b111010001011101;
		Coeff[11903] <= 15'b111010001011110;
		Coeff[11904] <= 15'b111010001100000;
		Coeff[11905] <= 15'b111010001100001;
		Coeff[11906] <= 15'b111010001100010;
		Coeff[11907] <= 15'b111010001100100;
		Coeff[11908] <= 15'b111010001100101;
		Coeff[11909] <= 15'b111010001100110;
		Coeff[11910] <= 15'b111010001100111;
		Coeff[11911] <= 15'b111010001101001;
		Coeff[11912] <= 15'b111010001101010;
		Coeff[11913] <= 15'b111010001101011;
		Coeff[11914] <= 15'b111010001101101;
		Coeff[11915] <= 15'b111010001101110;
		Coeff[11916] <= 15'b111010001101111;
		Coeff[11917] <= 15'b111010001110001;
		Coeff[11918] <= 15'b111010001110010;
		Coeff[11919] <= 15'b111010001110011;
		Coeff[11920] <= 15'b111010001110101;
		Coeff[11921] <= 15'b111010001110110;
		Coeff[11922] <= 15'b111010001110111;
		Coeff[11923] <= 15'b111010001111000;
		Coeff[11924] <= 15'b111010001111010;
		Coeff[11925] <= 15'b111010001111011;
		Coeff[11926] <= 15'b111010001111100;
		Coeff[11927] <= 15'b111010001111110;
		Coeff[11928] <= 15'b111010001111111;
		Coeff[11929] <= 15'b111010010000000;
		Coeff[11930] <= 15'b111010010000010;
		Coeff[11931] <= 15'b111010010000011;
		Coeff[11932] <= 15'b111010010000100;
		Coeff[11933] <= 15'b111010010000101;
		Coeff[11934] <= 15'b111010010000111;
		Coeff[11935] <= 15'b111010010001000;
		Coeff[11936] <= 15'b111010010001001;
		Coeff[11937] <= 15'b111010010001011;
		Coeff[11938] <= 15'b111010010001100;
		Coeff[11939] <= 15'b111010010001101;
		Coeff[11940] <= 15'b111010010001111;
		Coeff[11941] <= 15'b111010010010000;
		Coeff[11942] <= 15'b111010010010001;
		Coeff[11943] <= 15'b111010010010010;
		Coeff[11944] <= 15'b111010010010100;
		Coeff[11945] <= 15'b111010010010101;
		Coeff[11946] <= 15'b111010010010110;
		Coeff[11947] <= 15'b111010010011000;
		Coeff[11948] <= 15'b111010010011001;
		Coeff[11949] <= 15'b111010010011010;
		Coeff[11950] <= 15'b111010010011100;
		Coeff[11951] <= 15'b111010010011101;
		Coeff[11952] <= 15'b111010010011110;
		Coeff[11953] <= 15'b111010010011111;
		Coeff[11954] <= 15'b111010010100001;
		Coeff[11955] <= 15'b111010010100010;
		Coeff[11956] <= 15'b111010010100011;
		Coeff[11957] <= 15'b111010010100101;
		Coeff[11958] <= 15'b111010010100110;
		Coeff[11959] <= 15'b111010010100111;
		Coeff[11960] <= 15'b111010010101000;
		Coeff[11961] <= 15'b111010010101010;
		Coeff[11962] <= 15'b111010010101011;
		Coeff[11963] <= 15'b111010010101100;
		Coeff[11964] <= 15'b111010010101110;
		Coeff[11965] <= 15'b111010010101111;
		Coeff[11966] <= 15'b111010010110000;
		Coeff[11967] <= 15'b111010010110001;
		Coeff[11968] <= 15'b111010010110011;
		Coeff[11969] <= 15'b111010010110100;
		Coeff[11970] <= 15'b111010010110101;
		Coeff[11971] <= 15'b111010010110111;
		Coeff[11972] <= 15'b111010010111000;
		Coeff[11973] <= 15'b111010010111001;
		Coeff[11974] <= 15'b111010010111011;
		Coeff[11975] <= 15'b111010010111100;
		Coeff[11976] <= 15'b111010010111101;
		Coeff[11977] <= 15'b111010010111110;
		Coeff[11978] <= 15'b111010011000000;
		Coeff[11979] <= 15'b111010011000001;
		Coeff[11980] <= 15'b111010011000010;
		Coeff[11981] <= 15'b111010011000100;
		Coeff[11982] <= 15'b111010011000101;
		Coeff[11983] <= 15'b111010011000110;
		Coeff[11984] <= 15'b111010011000111;
		Coeff[11985] <= 15'b111010011001001;
		Coeff[11986] <= 15'b111010011001010;
		Coeff[11987] <= 15'b111010011001011;
		Coeff[11988] <= 15'b111010011001101;
		Coeff[11989] <= 15'b111010011001110;
		Coeff[11990] <= 15'b111010011001111;
		Coeff[11991] <= 15'b111010011010000;
		Coeff[11992] <= 15'b111010011010010;
		Coeff[11993] <= 15'b111010011010011;
		Coeff[11994] <= 15'b111010011010100;
		Coeff[11995] <= 15'b111010011010110;
		Coeff[11996] <= 15'b111010011010111;
		Coeff[11997] <= 15'b111010011011000;
		Coeff[11998] <= 15'b111010011011001;
		Coeff[11999] <= 15'b111010011011011;
		Coeff[12000] <= 15'b111010011011100;
		Coeff[12001] <= 15'b111010011011101;
		Coeff[12002] <= 15'b111010011011111;
		Coeff[12003] <= 15'b111010011100000;
		Coeff[12004] <= 15'b111010011100001;
		Coeff[12005] <= 15'b111010011100010;
		Coeff[12006] <= 15'b111010011100100;
		Coeff[12007] <= 15'b111010011100101;
		Coeff[12008] <= 15'b111010011100110;
		Coeff[12009] <= 15'b111010011100111;
		Coeff[12010] <= 15'b111010011101001;
		Coeff[12011] <= 15'b111010011101010;
		Coeff[12012] <= 15'b111010011101011;
		Coeff[12013] <= 15'b111010011101101;
		Coeff[12014] <= 15'b111010011101110;
		Coeff[12015] <= 15'b111010011101111;
		Coeff[12016] <= 15'b111010011110000;
		Coeff[12017] <= 15'b111010011110010;
		Coeff[12018] <= 15'b111010011110011;
		Coeff[12019] <= 15'b111010011110100;
		Coeff[12020] <= 15'b111010011110110;
		Coeff[12021] <= 15'b111010011110111;
		Coeff[12022] <= 15'b111010011111000;
		Coeff[12023] <= 15'b111010011111001;
		Coeff[12024] <= 15'b111010011111011;
		Coeff[12025] <= 15'b111010011111100;
		Coeff[12026] <= 15'b111010011111101;
		Coeff[12027] <= 15'b111010011111110;
		Coeff[12028] <= 15'b111010100000000;
		Coeff[12029] <= 15'b111010100000001;
		Coeff[12030] <= 15'b111010100000010;
		Coeff[12031] <= 15'b111010100000100;
		Coeff[12032] <= 15'b111010100000101;
		Coeff[12033] <= 15'b111010100000110;
		Coeff[12034] <= 15'b111010100000111;
		Coeff[12035] <= 15'b111010100001001;
		Coeff[12036] <= 15'b111010100001010;
		Coeff[12037] <= 15'b111010100001011;
		Coeff[12038] <= 15'b111010100001100;
		Coeff[12039] <= 15'b111010100001110;
		Coeff[12040] <= 15'b111010100001111;
		Coeff[12041] <= 15'b111010100010000;
		Coeff[12042] <= 15'b111010100010010;
		Coeff[12043] <= 15'b111010100010011;
		Coeff[12044] <= 15'b111010100010100;
		Coeff[12045] <= 15'b111010100010101;
		Coeff[12046] <= 15'b111010100010111;
		Coeff[12047] <= 15'b111010100011000;
		Coeff[12048] <= 15'b111010100011001;
		Coeff[12049] <= 15'b111010100011010;
		Coeff[12050] <= 15'b111010100011100;
		Coeff[12051] <= 15'b111010100011101;
		Coeff[12052] <= 15'b111010100011110;
		Coeff[12053] <= 15'b111010100011111;
		Coeff[12054] <= 15'b111010100100001;
		Coeff[12055] <= 15'b111010100100010;
		Coeff[12056] <= 15'b111010100100011;
		Coeff[12057] <= 15'b111010100100101;
		Coeff[12058] <= 15'b111010100100110;
		Coeff[12059] <= 15'b111010100100111;
		Coeff[12060] <= 15'b111010100101000;
		Coeff[12061] <= 15'b111010100101010;
		Coeff[12062] <= 15'b111010100101011;
		Coeff[12063] <= 15'b111010100101100;
		Coeff[12064] <= 15'b111010100101101;
		Coeff[12065] <= 15'b111010100101111;
		Coeff[12066] <= 15'b111010100110000;
		Coeff[12067] <= 15'b111010100110001;
		Coeff[12068] <= 15'b111010100110010;
		Coeff[12069] <= 15'b111010100110100;
		Coeff[12070] <= 15'b111010100110101;
		Coeff[12071] <= 15'b111010100110110;
		Coeff[12072] <= 15'b111010100111000;
		Coeff[12073] <= 15'b111010100111001;
		Coeff[12074] <= 15'b111010100111010;
		Coeff[12075] <= 15'b111010100111011;
		Coeff[12076] <= 15'b111010100111101;
		Coeff[12077] <= 15'b111010100111110;
		Coeff[12078] <= 15'b111010100111111;
		Coeff[12079] <= 15'b111010101000000;
		Coeff[12080] <= 15'b111010101000010;
		Coeff[12081] <= 15'b111010101000011;
		Coeff[12082] <= 15'b111010101000100;
		Coeff[12083] <= 15'b111010101000101;
		Coeff[12084] <= 15'b111010101000111;
		Coeff[12085] <= 15'b111010101001000;
		Coeff[12086] <= 15'b111010101001001;
		Coeff[12087] <= 15'b111010101001010;
		Coeff[12088] <= 15'b111010101001100;
		Coeff[12089] <= 15'b111010101001101;
		Coeff[12090] <= 15'b111010101001110;
		Coeff[12091] <= 15'b111010101001111;
		Coeff[12092] <= 15'b111010101010001;
		Coeff[12093] <= 15'b111010101010010;
		Coeff[12094] <= 15'b111010101010011;
		Coeff[12095] <= 15'b111010101010100;
		Coeff[12096] <= 15'b111010101010110;
		Coeff[12097] <= 15'b111010101010111;
		Coeff[12098] <= 15'b111010101011000;
		Coeff[12099] <= 15'b111010101011010;
		Coeff[12100] <= 15'b111010101011011;
		Coeff[12101] <= 15'b111010101011100;
		Coeff[12102] <= 15'b111010101011101;
		Coeff[12103] <= 15'b111010101011111;
		Coeff[12104] <= 15'b111010101100000;
		Coeff[12105] <= 15'b111010101100001;
		Coeff[12106] <= 15'b111010101100010;
		Coeff[12107] <= 15'b111010101100100;
		Coeff[12108] <= 15'b111010101100101;
		Coeff[12109] <= 15'b111010101100110;
		Coeff[12110] <= 15'b111010101100111;
		Coeff[12111] <= 15'b111010101101001;
		Coeff[12112] <= 15'b111010101101010;
		Coeff[12113] <= 15'b111010101101011;
		Coeff[12114] <= 15'b111010101101100;
		Coeff[12115] <= 15'b111010101101110;
		Coeff[12116] <= 15'b111010101101111;
		Coeff[12117] <= 15'b111010101110000;
		Coeff[12118] <= 15'b111010101110001;
		Coeff[12119] <= 15'b111010101110011;
		Coeff[12120] <= 15'b111010101110100;
		Coeff[12121] <= 15'b111010101110101;
		Coeff[12122] <= 15'b111010101110110;
		Coeff[12123] <= 15'b111010101111000;
		Coeff[12124] <= 15'b111010101111001;
		Coeff[12125] <= 15'b111010101111010;
		Coeff[12126] <= 15'b111010101111011;
		Coeff[12127] <= 15'b111010101111101;
		Coeff[12128] <= 15'b111010101111110;
		Coeff[12129] <= 15'b111010101111111;
		Coeff[12130] <= 15'b111010110000000;
		Coeff[12131] <= 15'b111010110000010;
		Coeff[12132] <= 15'b111010110000011;
		Coeff[12133] <= 15'b111010110000100;
		Coeff[12134] <= 15'b111010110000101;
		Coeff[12135] <= 15'b111010110000110;
		Coeff[12136] <= 15'b111010110001000;
		Coeff[12137] <= 15'b111010110001001;
		Coeff[12138] <= 15'b111010110001010;
		Coeff[12139] <= 15'b111010110001011;
		Coeff[12140] <= 15'b111010110001101;
		Coeff[12141] <= 15'b111010110001110;
		Coeff[12142] <= 15'b111010110001111;
		Coeff[12143] <= 15'b111010110010000;
		Coeff[12144] <= 15'b111010110010010;
		Coeff[12145] <= 15'b111010110010011;
		Coeff[12146] <= 15'b111010110010100;
		Coeff[12147] <= 15'b111010110010101;
		Coeff[12148] <= 15'b111010110010111;
		Coeff[12149] <= 15'b111010110011000;
		Coeff[12150] <= 15'b111010110011001;
		Coeff[12151] <= 15'b111010110011010;
		Coeff[12152] <= 15'b111010110011100;
		Coeff[12153] <= 15'b111010110011101;
		Coeff[12154] <= 15'b111010110011110;
		Coeff[12155] <= 15'b111010110011111;
		Coeff[12156] <= 15'b111010110100001;
		Coeff[12157] <= 15'b111010110100010;
		Coeff[12158] <= 15'b111010110100011;
		Coeff[12159] <= 15'b111010110100100;
		Coeff[12160] <= 15'b111010110100110;
		Coeff[12161] <= 15'b111010110100111;
		Coeff[12162] <= 15'b111010110101000;
		Coeff[12163] <= 15'b111010110101001;
		Coeff[12164] <= 15'b111010110101010;
		Coeff[12165] <= 15'b111010110101100;
		Coeff[12166] <= 15'b111010110101101;
		Coeff[12167] <= 15'b111010110101110;
		Coeff[12168] <= 15'b111010110101111;
		Coeff[12169] <= 15'b111010110110001;
		Coeff[12170] <= 15'b111010110110010;
		Coeff[12171] <= 15'b111010110110011;
		Coeff[12172] <= 15'b111010110110100;
		Coeff[12173] <= 15'b111010110110110;
		Coeff[12174] <= 15'b111010110110111;
		Coeff[12175] <= 15'b111010110111000;
		Coeff[12176] <= 15'b111010110111001;
		Coeff[12177] <= 15'b111010110111011;
		Coeff[12178] <= 15'b111010110111100;
		Coeff[12179] <= 15'b111010110111101;
		Coeff[12180] <= 15'b111010110111110;
		Coeff[12181] <= 15'b111010110111111;
		Coeff[12182] <= 15'b111010111000001;
		Coeff[12183] <= 15'b111010111000010;
		Coeff[12184] <= 15'b111010111000011;
		Coeff[12185] <= 15'b111010111000100;
		Coeff[12186] <= 15'b111010111000110;
		Coeff[12187] <= 15'b111010111000111;
		Coeff[12188] <= 15'b111010111001000;
		Coeff[12189] <= 15'b111010111001001;
		Coeff[12190] <= 15'b111010111001011;
		Coeff[12191] <= 15'b111010111001100;
		Coeff[12192] <= 15'b111010111001101;
		Coeff[12193] <= 15'b111010111001110;
		Coeff[12194] <= 15'b111010111001111;
		Coeff[12195] <= 15'b111010111010001;
		Coeff[12196] <= 15'b111010111010010;
		Coeff[12197] <= 15'b111010111010011;
		Coeff[12198] <= 15'b111010111010100;
		Coeff[12199] <= 15'b111010111010110;
		Coeff[12200] <= 15'b111010111010111;
		Coeff[12201] <= 15'b111010111011000;
		Coeff[12202] <= 15'b111010111011001;
		Coeff[12203] <= 15'b111010111011010;
		Coeff[12204] <= 15'b111010111011100;
		Coeff[12205] <= 15'b111010111011101;
		Coeff[12206] <= 15'b111010111011110;
		Coeff[12207] <= 15'b111010111011111;
		Coeff[12208] <= 15'b111010111100001;
		Coeff[12209] <= 15'b111010111100010;
		Coeff[12210] <= 15'b111010111100011;
		Coeff[12211] <= 15'b111010111100100;
		Coeff[12212] <= 15'b111010111100110;
		Coeff[12213] <= 15'b111010111100111;
		Coeff[12214] <= 15'b111010111101000;
		Coeff[12215] <= 15'b111010111101001;
		Coeff[12216] <= 15'b111010111101010;
		Coeff[12217] <= 15'b111010111101100;
		Coeff[12218] <= 15'b111010111101101;
		Coeff[12219] <= 15'b111010111101110;
		Coeff[12220] <= 15'b111010111101111;
		Coeff[12221] <= 15'b111010111110001;
		Coeff[12222] <= 15'b111010111110010;
		Coeff[12223] <= 15'b111010111110011;
		Coeff[12224] <= 15'b111010111110100;
		Coeff[12225] <= 15'b111010111110101;
		Coeff[12226] <= 15'b111010111110111;
		Coeff[12227] <= 15'b111010111111000;
		Coeff[12228] <= 15'b111010111111001;
		Coeff[12229] <= 15'b111010111111010;
		Coeff[12230] <= 15'b111010111111011;
		Coeff[12231] <= 15'b111010111111101;
		Coeff[12232] <= 15'b111010111111110;
		Coeff[12233] <= 15'b111010111111111;
		Coeff[12234] <= 15'b111011000000000;
		Coeff[12235] <= 15'b111011000000010;
		Coeff[12236] <= 15'b111011000000011;
		Coeff[12237] <= 15'b111011000000100;
		Coeff[12238] <= 15'b111011000000101;
		Coeff[12239] <= 15'b111011000000110;
		Coeff[12240] <= 15'b111011000001000;
		Coeff[12241] <= 15'b111011000001001;
		Coeff[12242] <= 15'b111011000001010;
		Coeff[12243] <= 15'b111011000001011;
		Coeff[12244] <= 15'b111011000001101;
		Coeff[12245] <= 15'b111011000001110;
		Coeff[12246] <= 15'b111011000001111;
		Coeff[12247] <= 15'b111011000010000;
		Coeff[12248] <= 15'b111011000010001;
		Coeff[12249] <= 15'b111011000010011;
		Coeff[12250] <= 15'b111011000010100;
		Coeff[12251] <= 15'b111011000010101;
		Coeff[12252] <= 15'b111011000010110;
		Coeff[12253] <= 15'b111011000010111;
		Coeff[12254] <= 15'b111011000011001;
		Coeff[12255] <= 15'b111011000011010;
		Coeff[12256] <= 15'b111011000011011;
		Coeff[12257] <= 15'b111011000011100;
		Coeff[12258] <= 15'b111011000011101;
		Coeff[12259] <= 15'b111011000011111;
		Coeff[12260] <= 15'b111011000100000;
		Coeff[12261] <= 15'b111011000100001;
		Coeff[12262] <= 15'b111011000100010;
		Coeff[12263] <= 15'b111011000100100;
		Coeff[12264] <= 15'b111011000100101;
		Coeff[12265] <= 15'b111011000100110;
		Coeff[12266] <= 15'b111011000100111;
		Coeff[12267] <= 15'b111011000101000;
		Coeff[12268] <= 15'b111011000101010;
		Coeff[12269] <= 15'b111011000101011;
		Coeff[12270] <= 15'b111011000101100;
		Coeff[12271] <= 15'b111011000101101;
		Coeff[12272] <= 15'b111011000101110;
		Coeff[12273] <= 15'b111011000110000;
		Coeff[12274] <= 15'b111011000110001;
		Coeff[12275] <= 15'b111011000110010;
		Coeff[12276] <= 15'b111011000110011;
		Coeff[12277] <= 15'b111011000110100;
		Coeff[12278] <= 15'b111011000110110;
		Coeff[12279] <= 15'b111011000110111;
		Coeff[12280] <= 15'b111011000111000;
		Coeff[12281] <= 15'b111011000111001;
		Coeff[12282] <= 15'b111011000111010;
		Coeff[12283] <= 15'b111011000111100;
		Coeff[12284] <= 15'b111011000111101;
		Coeff[12285] <= 15'b111011000111110;
		Coeff[12286] <= 15'b111011000111111;
		Coeff[12287] <= 15'b111011001000000;
		Coeff[12288] <= 15'b111011001000010;
		Coeff[12289] <= 15'b111011001000011;
		Coeff[12290] <= 15'b111011001000100;
		Coeff[12291] <= 15'b111011001000101;
		Coeff[12292] <= 15'b111011001000110;
		Coeff[12293] <= 15'b111011001001000;
		Coeff[12294] <= 15'b111011001001001;
		Coeff[12295] <= 15'b111011001001010;
		Coeff[12296] <= 15'b111011001001011;
		Coeff[12297] <= 15'b111011001001100;
		Coeff[12298] <= 15'b111011001001110;
		Coeff[12299] <= 15'b111011001001111;
		Coeff[12300] <= 15'b111011001010000;
		Coeff[12301] <= 15'b111011001010001;
		Coeff[12302] <= 15'b111011001010010;
		Coeff[12303] <= 15'b111011001010100;
		Coeff[12304] <= 15'b111011001010101;
		Coeff[12305] <= 15'b111011001010110;
		Coeff[12306] <= 15'b111011001010111;
		Coeff[12307] <= 15'b111011001011000;
		Coeff[12308] <= 15'b111011001011010;
		Coeff[12309] <= 15'b111011001011011;
		Coeff[12310] <= 15'b111011001011100;
		Coeff[12311] <= 15'b111011001011101;
		Coeff[12312] <= 15'b111011001011110;
		Coeff[12313] <= 15'b111011001100000;
		Coeff[12314] <= 15'b111011001100001;
		Coeff[12315] <= 15'b111011001100010;
		Coeff[12316] <= 15'b111011001100011;
		Coeff[12317] <= 15'b111011001100100;
		Coeff[12318] <= 15'b111011001100110;
		Coeff[12319] <= 15'b111011001100111;
		Coeff[12320] <= 15'b111011001101000;
		Coeff[12321] <= 15'b111011001101001;
		Coeff[12322] <= 15'b111011001101010;
		Coeff[12323] <= 15'b111011001101100;
		Coeff[12324] <= 15'b111011001101101;
		Coeff[12325] <= 15'b111011001101110;
		Coeff[12326] <= 15'b111011001101111;
		Coeff[12327] <= 15'b111011001110000;
		Coeff[12328] <= 15'b111011001110010;
		Coeff[12329] <= 15'b111011001110011;
		Coeff[12330] <= 15'b111011001110100;
		Coeff[12331] <= 15'b111011001110101;
		Coeff[12332] <= 15'b111011001110110;
		Coeff[12333] <= 15'b111011001111000;
		Coeff[12334] <= 15'b111011001111001;
		Coeff[12335] <= 15'b111011001111010;
		Coeff[12336] <= 15'b111011001111011;
		Coeff[12337] <= 15'b111011001111100;
		Coeff[12338] <= 15'b111011001111101;
		Coeff[12339] <= 15'b111011001111111;
		Coeff[12340] <= 15'b111011010000000;
		Coeff[12341] <= 15'b111011010000001;
		Coeff[12342] <= 15'b111011010000010;
		Coeff[12343] <= 15'b111011010000011;
		Coeff[12344] <= 15'b111011010000101;
		Coeff[12345] <= 15'b111011010000110;
		Coeff[12346] <= 15'b111011010000111;
		Coeff[12347] <= 15'b111011010001000;
		Coeff[12348] <= 15'b111011010001001;
		Coeff[12349] <= 15'b111011010001011;
		Coeff[12350] <= 15'b111011010001100;
		Coeff[12351] <= 15'b111011010001101;
		Coeff[12352] <= 15'b111011010001110;
		Coeff[12353] <= 15'b111011010001111;
		Coeff[12354] <= 15'b111011010010000;
		Coeff[12355] <= 15'b111011010010010;
		Coeff[12356] <= 15'b111011010010011;
		Coeff[12357] <= 15'b111011010010100;
		Coeff[12358] <= 15'b111011010010101;
		Coeff[12359] <= 15'b111011010010110;
		Coeff[12360] <= 15'b111011010011000;
		Coeff[12361] <= 15'b111011010011001;
		Coeff[12362] <= 15'b111011010011010;
		Coeff[12363] <= 15'b111011010011011;
		Coeff[12364] <= 15'b111011010011100;
		Coeff[12365] <= 15'b111011010011101;
		Coeff[12366] <= 15'b111011010011111;
		Coeff[12367] <= 15'b111011010100000;
		Coeff[12368] <= 15'b111011010100001;
		Coeff[12369] <= 15'b111011010100010;
		Coeff[12370] <= 15'b111011010100011;
		Coeff[12371] <= 15'b111011010100101;
		Coeff[12372] <= 15'b111011010100110;
		Coeff[12373] <= 15'b111011010100111;
		Coeff[12374] <= 15'b111011010101000;
		Coeff[12375] <= 15'b111011010101001;
		Coeff[12376] <= 15'b111011010101010;
		Coeff[12377] <= 15'b111011010101100;
		Coeff[12378] <= 15'b111011010101101;
		Coeff[12379] <= 15'b111011010101110;
		Coeff[12380] <= 15'b111011010101111;
		Coeff[12381] <= 15'b111011010110000;
		Coeff[12382] <= 15'b111011010110001;
		Coeff[12383] <= 15'b111011010110011;
		Coeff[12384] <= 15'b111011010110100;
		Coeff[12385] <= 15'b111011010110101;
		Coeff[12386] <= 15'b111011010110110;
		Coeff[12387] <= 15'b111011010110111;
		Coeff[12388] <= 15'b111011010111001;
		Coeff[12389] <= 15'b111011010111010;
		Coeff[12390] <= 15'b111011010111011;
		Coeff[12391] <= 15'b111011010111100;
		Coeff[12392] <= 15'b111011010111101;
		Coeff[12393] <= 15'b111011010111110;
		Coeff[12394] <= 15'b111011011000000;
		Coeff[12395] <= 15'b111011011000001;
		Coeff[12396] <= 15'b111011011000010;
		Coeff[12397] <= 15'b111011011000011;
		Coeff[12398] <= 15'b111011011000100;
		Coeff[12399] <= 15'b111011011000101;
		Coeff[12400] <= 15'b111011011000111;
		Coeff[12401] <= 15'b111011011001000;
		Coeff[12402] <= 15'b111011011001001;
		Coeff[12403] <= 15'b111011011001010;
		Coeff[12404] <= 15'b111011011001011;
		Coeff[12405] <= 15'b111011011001100;
		Coeff[12406] <= 15'b111011011001110;
		Coeff[12407] <= 15'b111011011001111;
		Coeff[12408] <= 15'b111011011010000;
		Coeff[12409] <= 15'b111011011010001;
		Coeff[12410] <= 15'b111011011010010;
		Coeff[12411] <= 15'b111011011010011;
		Coeff[12412] <= 15'b111011011010101;
		Coeff[12413] <= 15'b111011011010110;
		Coeff[12414] <= 15'b111011011010111;
		Coeff[12415] <= 15'b111011011011000;
		Coeff[12416] <= 15'b111011011011001;
		Coeff[12417] <= 15'b111011011011010;
		Coeff[12418] <= 15'b111011011011100;
		Coeff[12419] <= 15'b111011011011101;
		Coeff[12420] <= 15'b111011011011110;
		Coeff[12421] <= 15'b111011011011111;
		Coeff[12422] <= 15'b111011011100000;
		Coeff[12423] <= 15'b111011011100001;
		Coeff[12424] <= 15'b111011011100011;
		Coeff[12425] <= 15'b111011011100100;
		Coeff[12426] <= 15'b111011011100101;
		Coeff[12427] <= 15'b111011011100110;
		Coeff[12428] <= 15'b111011011100111;
		Coeff[12429] <= 15'b111011011101000;
		Coeff[12430] <= 15'b111011011101010;
		Coeff[12431] <= 15'b111011011101011;
		Coeff[12432] <= 15'b111011011101100;
		Coeff[12433] <= 15'b111011011101101;
		Coeff[12434] <= 15'b111011011101110;
		Coeff[12435] <= 15'b111011011101111;
		Coeff[12436] <= 15'b111011011110001;
		Coeff[12437] <= 15'b111011011110010;
		Coeff[12438] <= 15'b111011011110011;
		Coeff[12439] <= 15'b111011011110100;
		Coeff[12440] <= 15'b111011011110101;
		Coeff[12441] <= 15'b111011011110110;
		Coeff[12442] <= 15'b111011011111000;
		Coeff[12443] <= 15'b111011011111001;
		Coeff[12444] <= 15'b111011011111010;
		Coeff[12445] <= 15'b111011011111011;
		Coeff[12446] <= 15'b111011011111100;
		Coeff[12447] <= 15'b111011011111101;
		Coeff[12448] <= 15'b111011011111110;
		Coeff[12449] <= 15'b111011100000000;
		Coeff[12450] <= 15'b111011100000001;
		Coeff[12451] <= 15'b111011100000010;
		Coeff[12452] <= 15'b111011100000011;
		Coeff[12453] <= 15'b111011100000100;
		Coeff[12454] <= 15'b111011100000101;
		Coeff[12455] <= 15'b111011100000111;
		Coeff[12456] <= 15'b111011100001000;
		Coeff[12457] <= 15'b111011100001001;
		Coeff[12458] <= 15'b111011100001010;
		Coeff[12459] <= 15'b111011100001011;
		Coeff[12460] <= 15'b111011100001100;
		Coeff[12461] <= 15'b111011100001101;
		Coeff[12462] <= 15'b111011100001111;
		Coeff[12463] <= 15'b111011100010000;
		Coeff[12464] <= 15'b111011100010001;
		Coeff[12465] <= 15'b111011100010010;
		Coeff[12466] <= 15'b111011100010011;
		Coeff[12467] <= 15'b111011100010100;
		Coeff[12468] <= 15'b111011100010110;
		Coeff[12469] <= 15'b111011100010111;
		Coeff[12470] <= 15'b111011100011000;
		Coeff[12471] <= 15'b111011100011001;
		Coeff[12472] <= 15'b111011100011010;
		Coeff[12473] <= 15'b111011100011011;
		Coeff[12474] <= 15'b111011100011100;
		Coeff[12475] <= 15'b111011100011110;
		Coeff[12476] <= 15'b111011100011111;
		Coeff[12477] <= 15'b111011100100000;
		Coeff[12478] <= 15'b111011100100001;
		Coeff[12479] <= 15'b111011100100010;
		Coeff[12480] <= 15'b111011100100011;
		Coeff[12481] <= 15'b111011100100101;
		Coeff[12482] <= 15'b111011100100110;
		Coeff[12483] <= 15'b111011100100111;
		Coeff[12484] <= 15'b111011100101000;
		Coeff[12485] <= 15'b111011100101001;
		Coeff[12486] <= 15'b111011100101010;
		Coeff[12487] <= 15'b111011100101011;
		Coeff[12488] <= 15'b111011100101101;
		Coeff[12489] <= 15'b111011100101110;
		Coeff[12490] <= 15'b111011100101111;
		Coeff[12491] <= 15'b111011100110000;
		Coeff[12492] <= 15'b111011100110001;
		Coeff[12493] <= 15'b111011100110010;
		Coeff[12494] <= 15'b111011100110011;
		Coeff[12495] <= 15'b111011100110101;
		Coeff[12496] <= 15'b111011100110110;
		Coeff[12497] <= 15'b111011100110111;
		Coeff[12498] <= 15'b111011100111000;
		Coeff[12499] <= 15'b111011100111001;
		Coeff[12500] <= 15'b111011100111010;
		Coeff[12501] <= 15'b111011100111011;
		Coeff[12502] <= 15'b111011100111101;
		Coeff[12503] <= 15'b111011100111110;
		Coeff[12504] <= 15'b111011100111111;
		Coeff[12505] <= 15'b111011101000000;
		Coeff[12506] <= 15'b111011101000001;
		Coeff[12507] <= 15'b111011101000010;
		Coeff[12508] <= 15'b111011101000011;
		Coeff[12509] <= 15'b111011101000101;
		Coeff[12510] <= 15'b111011101000110;
		Coeff[12511] <= 15'b111011101000111;
		Coeff[12512] <= 15'b111011101001000;
		Coeff[12513] <= 15'b111011101001001;
		Coeff[12514] <= 15'b111011101001010;
		Coeff[12515] <= 15'b111011101001011;
		Coeff[12516] <= 15'b111011101001101;
		Coeff[12517] <= 15'b111011101001110;
		Coeff[12518] <= 15'b111011101001111;
		Coeff[12519] <= 15'b111011101010000;
		Coeff[12520] <= 15'b111011101010001;
		Coeff[12521] <= 15'b111011101010010;
		Coeff[12522] <= 15'b111011101010011;
		Coeff[12523] <= 15'b111011101010101;
		Coeff[12524] <= 15'b111011101010110;
		Coeff[12525] <= 15'b111011101010111;
		Coeff[12526] <= 15'b111011101011000;
		Coeff[12527] <= 15'b111011101011001;
		Coeff[12528] <= 15'b111011101011010;
		Coeff[12529] <= 15'b111011101011011;
		Coeff[12530] <= 15'b111011101011100;
		Coeff[12531] <= 15'b111011101011110;
		Coeff[12532] <= 15'b111011101011111;
		Coeff[12533] <= 15'b111011101100000;
		Coeff[12534] <= 15'b111011101100001;
		Coeff[12535] <= 15'b111011101100010;
		Coeff[12536] <= 15'b111011101100011;
		Coeff[12537] <= 15'b111011101100100;
		Coeff[12538] <= 15'b111011101100110;
		Coeff[12539] <= 15'b111011101100111;
		Coeff[12540] <= 15'b111011101101000;
		Coeff[12541] <= 15'b111011101101001;
		Coeff[12542] <= 15'b111011101101010;
		Coeff[12543] <= 15'b111011101101011;
		Coeff[12544] <= 15'b111011101101100;
		Coeff[12545] <= 15'b111011101101101;
		Coeff[12546] <= 15'b111011101101111;
		Coeff[12547] <= 15'b111011101110000;
		Coeff[12548] <= 15'b111011101110001;
		Coeff[12549] <= 15'b111011101110010;
		Coeff[12550] <= 15'b111011101110011;
		Coeff[12551] <= 15'b111011101110100;
		Coeff[12552] <= 15'b111011101110101;
		Coeff[12553] <= 15'b111011101110110;
		Coeff[12554] <= 15'b111011101111000;
		Coeff[12555] <= 15'b111011101111001;
		Coeff[12556] <= 15'b111011101111010;
		Coeff[12557] <= 15'b111011101111011;
		Coeff[12558] <= 15'b111011101111100;
		Coeff[12559] <= 15'b111011101111101;
		Coeff[12560] <= 15'b111011101111110;
		Coeff[12561] <= 15'b111011101111111;
		Coeff[12562] <= 15'b111011110000001;
		Coeff[12563] <= 15'b111011110000010;
		Coeff[12564] <= 15'b111011110000011;
		Coeff[12565] <= 15'b111011110000100;
		Coeff[12566] <= 15'b111011110000101;
		Coeff[12567] <= 15'b111011110000110;
		Coeff[12568] <= 15'b111011110000111;
		Coeff[12569] <= 15'b111011110001000;
		Coeff[12570] <= 15'b111011110001010;
		Coeff[12571] <= 15'b111011110001011;
		Coeff[12572] <= 15'b111011110001100;
		Coeff[12573] <= 15'b111011110001101;
		Coeff[12574] <= 15'b111011110001110;
		Coeff[12575] <= 15'b111011110001111;
		Coeff[12576] <= 15'b111011110010000;
		Coeff[12577] <= 15'b111011110010001;
		Coeff[12578] <= 15'b111011110010011;
		Coeff[12579] <= 15'b111011110010100;
		Coeff[12580] <= 15'b111011110010101;
		Coeff[12581] <= 15'b111011110010110;
		Coeff[12582] <= 15'b111011110010111;
		Coeff[12583] <= 15'b111011110011000;
		Coeff[12584] <= 15'b111011110011001;
		Coeff[12585] <= 15'b111011110011010;
		Coeff[12586] <= 15'b111011110011100;
		Coeff[12587] <= 15'b111011110011101;
		Coeff[12588] <= 15'b111011110011110;
		Coeff[12589] <= 15'b111011110011111;
		Coeff[12590] <= 15'b111011110100000;
		Coeff[12591] <= 15'b111011110100001;
		Coeff[12592] <= 15'b111011110100010;
		Coeff[12593] <= 15'b111011110100011;
		Coeff[12594] <= 15'b111011110100100;
		Coeff[12595] <= 15'b111011110100110;
		Coeff[12596] <= 15'b111011110100111;
		Coeff[12597] <= 15'b111011110101000;
		Coeff[12598] <= 15'b111011110101001;
		Coeff[12599] <= 15'b111011110101010;
		Coeff[12600] <= 15'b111011110101011;
		Coeff[12601] <= 15'b111011110101100;
		Coeff[12602] <= 15'b111011110101101;
		Coeff[12603] <= 15'b111011110101111;
		Coeff[12604] <= 15'b111011110110000;
		Coeff[12605] <= 15'b111011110110001;
		Coeff[12606] <= 15'b111011110110010;
		Coeff[12607] <= 15'b111011110110011;
		Coeff[12608] <= 15'b111011110110100;
		Coeff[12609] <= 15'b111011110110101;
		Coeff[12610] <= 15'b111011110110110;
		Coeff[12611] <= 15'b111011110110111;
		Coeff[12612] <= 15'b111011110111001;
		Coeff[12613] <= 15'b111011110111010;
		Coeff[12614] <= 15'b111011110111011;
		Coeff[12615] <= 15'b111011110111100;
		Coeff[12616] <= 15'b111011110111101;
		Coeff[12617] <= 15'b111011110111110;
		Coeff[12618] <= 15'b111011110111111;
		Coeff[12619] <= 15'b111011111000000;
		Coeff[12620] <= 15'b111011111000001;
		Coeff[12621] <= 15'b111011111000011;
		Coeff[12622] <= 15'b111011111000100;
		Coeff[12623] <= 15'b111011111000101;
		Coeff[12624] <= 15'b111011111000110;
		Coeff[12625] <= 15'b111011111000111;
		Coeff[12626] <= 15'b111011111001000;
		Coeff[12627] <= 15'b111011111001001;
		Coeff[12628] <= 15'b111011111001010;
		Coeff[12629] <= 15'b111011111001011;
		Coeff[12630] <= 15'b111011111001101;
		Coeff[12631] <= 15'b111011111001110;
		Coeff[12632] <= 15'b111011111001111;
		Coeff[12633] <= 15'b111011111010000;
		Coeff[12634] <= 15'b111011111010001;
		Coeff[12635] <= 15'b111011111010010;
		Coeff[12636] <= 15'b111011111010011;
		Coeff[12637] <= 15'b111011111010100;
		Coeff[12638] <= 15'b111011111010101;
		Coeff[12639] <= 15'b111011111010110;
		Coeff[12640] <= 15'b111011111011000;
		Coeff[12641] <= 15'b111011111011001;
		Coeff[12642] <= 15'b111011111011010;
		Coeff[12643] <= 15'b111011111011011;
		Coeff[12644] <= 15'b111011111011100;
		Coeff[12645] <= 15'b111011111011101;
		Coeff[12646] <= 15'b111011111011110;
		Coeff[12647] <= 15'b111011111011111;
		Coeff[12648] <= 15'b111011111100000;
		Coeff[12649] <= 15'b111011111100001;
		Coeff[12650] <= 15'b111011111100011;
		Coeff[12651] <= 15'b111011111100100;
		Coeff[12652] <= 15'b111011111100101;
		Coeff[12653] <= 15'b111011111100110;
		Coeff[12654] <= 15'b111011111100111;
		Coeff[12655] <= 15'b111011111101000;
		Coeff[12656] <= 15'b111011111101001;
		Coeff[12657] <= 15'b111011111101010;
		Coeff[12658] <= 15'b111011111101011;
		Coeff[12659] <= 15'b111011111101100;
		Coeff[12660] <= 15'b111011111101110;
		Coeff[12661] <= 15'b111011111101111;
		Coeff[12662] <= 15'b111011111110000;
		Coeff[12663] <= 15'b111011111110001;
		Coeff[12664] <= 15'b111011111110010;
		Coeff[12665] <= 15'b111011111110011;
		Coeff[12666] <= 15'b111011111110100;
		Coeff[12667] <= 15'b111011111110101;
		Coeff[12668] <= 15'b111011111110110;
		Coeff[12669] <= 15'b111011111110111;
		Coeff[12670] <= 15'b111011111111001;
		Coeff[12671] <= 15'b111011111111010;
		Coeff[12672] <= 15'b111011111111011;
		Coeff[12673] <= 15'b111011111111100;
		Coeff[12674] <= 15'b111011111111101;
		Coeff[12675] <= 15'b111011111111110;
		Coeff[12676] <= 15'b111011111111111;
		Coeff[12677] <= 15'b111100000000000;
		Coeff[12678] <= 15'b111100000000001;
		Coeff[12679] <= 15'b111100000000010;
		Coeff[12680] <= 15'b111100000000011;
		Coeff[12681] <= 15'b111100000000101;
		Coeff[12682] <= 15'b111100000000110;
		Coeff[12683] <= 15'b111100000000111;
		Coeff[12684] <= 15'b111100000001000;
		Coeff[12685] <= 15'b111100000001001;
		Coeff[12686] <= 15'b111100000001010;
		Coeff[12687] <= 15'b111100000001011;
		Coeff[12688] <= 15'b111100000001100;
		Coeff[12689] <= 15'b111100000001101;
		Coeff[12690] <= 15'b111100000001110;
		Coeff[12691] <= 15'b111100000001111;
		Coeff[12692] <= 15'b111100000010001;
		Coeff[12693] <= 15'b111100000010010;
		Coeff[12694] <= 15'b111100000010011;
		Coeff[12695] <= 15'b111100000010100;
		Coeff[12696] <= 15'b111100000010101;
		Coeff[12697] <= 15'b111100000010110;
		Coeff[12698] <= 15'b111100000010111;
		Coeff[12699] <= 15'b111100000011000;
		Coeff[12700] <= 15'b111100000011001;
		Coeff[12701] <= 15'b111100000011010;
		Coeff[12702] <= 15'b111100000011011;
		Coeff[12703] <= 15'b111100000011101;
		Coeff[12704] <= 15'b111100000011110;
		Coeff[12705] <= 15'b111100000011111;
		Coeff[12706] <= 15'b111100000100000;
		Coeff[12707] <= 15'b111100000100001;
		Coeff[12708] <= 15'b111100000100010;
		Coeff[12709] <= 15'b111100000100011;
		Coeff[12710] <= 15'b111100000100100;
		Coeff[12711] <= 15'b111100000100101;
		Coeff[12712] <= 15'b111100000100110;
		Coeff[12713] <= 15'b111100000100111;
		Coeff[12714] <= 15'b111100000101000;
		Coeff[12715] <= 15'b111100000101010;
		Coeff[12716] <= 15'b111100000101011;
		Coeff[12717] <= 15'b111100000101100;
		Coeff[12718] <= 15'b111100000101101;
		Coeff[12719] <= 15'b111100000101110;
		Coeff[12720] <= 15'b111100000101111;
		Coeff[12721] <= 15'b111100000110000;
		Coeff[12722] <= 15'b111100000110001;
		Coeff[12723] <= 15'b111100000110010;
		Coeff[12724] <= 15'b111100000110011;
		Coeff[12725] <= 15'b111100000110100;
		Coeff[12726] <= 15'b111100000110101;
		Coeff[12727] <= 15'b111100000110110;
		Coeff[12728] <= 15'b111100000111000;
		Coeff[12729] <= 15'b111100000111001;
		Coeff[12730] <= 15'b111100000111010;
		Coeff[12731] <= 15'b111100000111011;
		Coeff[12732] <= 15'b111100000111100;
		Coeff[12733] <= 15'b111100000111101;
		Coeff[12734] <= 15'b111100000111110;
		Coeff[12735] <= 15'b111100000111111;
		Coeff[12736] <= 15'b111100001000000;
		Coeff[12737] <= 15'b111100001000001;
		Coeff[12738] <= 15'b111100001000010;
		Coeff[12739] <= 15'b111100001000011;
		Coeff[12740] <= 15'b111100001000101;
		Coeff[12741] <= 15'b111100001000110;
		Coeff[12742] <= 15'b111100001000111;
		Coeff[12743] <= 15'b111100001001000;
		Coeff[12744] <= 15'b111100001001001;
		Coeff[12745] <= 15'b111100001001010;
		Coeff[12746] <= 15'b111100001001011;
		Coeff[12747] <= 15'b111100001001100;
		Coeff[12748] <= 15'b111100001001101;
		Coeff[12749] <= 15'b111100001001110;
		Coeff[12750] <= 15'b111100001001111;
		Coeff[12751] <= 15'b111100001010000;
		Coeff[12752] <= 15'b111100001010001;
		Coeff[12753] <= 15'b111100001010010;
		Coeff[12754] <= 15'b111100001010100;
		Coeff[12755] <= 15'b111100001010101;
		Coeff[12756] <= 15'b111100001010110;
		Coeff[12757] <= 15'b111100001010111;
		Coeff[12758] <= 15'b111100001011000;
		Coeff[12759] <= 15'b111100001011001;
		Coeff[12760] <= 15'b111100001011010;
		Coeff[12761] <= 15'b111100001011011;
		Coeff[12762] <= 15'b111100001011100;
		Coeff[12763] <= 15'b111100001011101;
		Coeff[12764] <= 15'b111100001011110;
		Coeff[12765] <= 15'b111100001011111;
		Coeff[12766] <= 15'b111100001100000;
		Coeff[12767] <= 15'b111100001100001;
		Coeff[12768] <= 15'b111100001100011;
		Coeff[12769] <= 15'b111100001100100;
		Coeff[12770] <= 15'b111100001100101;
		Coeff[12771] <= 15'b111100001100110;
		Coeff[12772] <= 15'b111100001100111;
		Coeff[12773] <= 15'b111100001101000;
		Coeff[12774] <= 15'b111100001101001;
		Coeff[12775] <= 15'b111100001101010;
		Coeff[12776] <= 15'b111100001101011;
		Coeff[12777] <= 15'b111100001101100;
		Coeff[12778] <= 15'b111100001101101;
		Coeff[12779] <= 15'b111100001101110;
		Coeff[12780] <= 15'b111100001101111;
		Coeff[12781] <= 15'b111100001110000;
		Coeff[12782] <= 15'b111100001110001;
		Coeff[12783] <= 15'b111100001110010;
		Coeff[12784] <= 15'b111100001110100;
		Coeff[12785] <= 15'b111100001110101;
		Coeff[12786] <= 15'b111100001110110;
		Coeff[12787] <= 15'b111100001110111;
		Coeff[12788] <= 15'b111100001111000;
		Coeff[12789] <= 15'b111100001111001;
		Coeff[12790] <= 15'b111100001111010;
		Coeff[12791] <= 15'b111100001111011;
		Coeff[12792] <= 15'b111100001111100;
		Coeff[12793] <= 15'b111100001111101;
		Coeff[12794] <= 15'b111100001111110;
		Coeff[12795] <= 15'b111100001111111;
		Coeff[12796] <= 15'b111100010000000;
		Coeff[12797] <= 15'b111100010000001;
		Coeff[12798] <= 15'b111100010000010;
		Coeff[12799] <= 15'b111100010000011;
		Coeff[12800] <= 15'b111100010000101;
		Coeff[12801] <= 15'b111100010000110;
		Coeff[12802] <= 15'b111100010000111;
		Coeff[12803] <= 15'b111100010001000;
		Coeff[12804] <= 15'b111100010001001;
		Coeff[12805] <= 15'b111100010001010;
		Coeff[12806] <= 15'b111100010001011;
		Coeff[12807] <= 15'b111100010001100;
		Coeff[12808] <= 15'b111100010001101;
		Coeff[12809] <= 15'b111100010001110;
		Coeff[12810] <= 15'b111100010001111;
		Coeff[12811] <= 15'b111100010010000;
		Coeff[12812] <= 15'b111100010010001;
		Coeff[12813] <= 15'b111100010010010;
		Coeff[12814] <= 15'b111100010010011;
		Coeff[12815] <= 15'b111100010010100;
		Coeff[12816] <= 15'b111100010010101;
		Coeff[12817] <= 15'b111100010010110;
		Coeff[12818] <= 15'b111100010011000;
		Coeff[12819] <= 15'b111100010011001;
		Coeff[12820] <= 15'b111100010011010;
		Coeff[12821] <= 15'b111100010011011;
		Coeff[12822] <= 15'b111100010011100;
		Coeff[12823] <= 15'b111100010011101;
		Coeff[12824] <= 15'b111100010011110;
		Coeff[12825] <= 15'b111100010011111;
		Coeff[12826] <= 15'b111100010100000;
		Coeff[12827] <= 15'b111100010100001;
		Coeff[12828] <= 15'b111100010100010;
		Coeff[12829] <= 15'b111100010100011;
		Coeff[12830] <= 15'b111100010100100;
		Coeff[12831] <= 15'b111100010100101;
		Coeff[12832] <= 15'b111100010100110;
		Coeff[12833] <= 15'b111100010100111;
		Coeff[12834] <= 15'b111100010101000;
		Coeff[12835] <= 15'b111100010101001;
		Coeff[12836] <= 15'b111100010101010;
		Coeff[12837] <= 15'b111100010101011;
		Coeff[12838] <= 15'b111100010101101;
		Coeff[12839] <= 15'b111100010101110;
		Coeff[12840] <= 15'b111100010101111;
		Coeff[12841] <= 15'b111100010110000;
		Coeff[12842] <= 15'b111100010110001;
		Coeff[12843] <= 15'b111100010110010;
		Coeff[12844] <= 15'b111100010110011;
		Coeff[12845] <= 15'b111100010110100;
		Coeff[12846] <= 15'b111100010110101;
		Coeff[12847] <= 15'b111100010110110;
		Coeff[12848] <= 15'b111100010110111;
		Coeff[12849] <= 15'b111100010111000;
		Coeff[12850] <= 15'b111100010111001;
		Coeff[12851] <= 15'b111100010111010;
		Coeff[12852] <= 15'b111100010111011;
		Coeff[12853] <= 15'b111100010111100;
		Coeff[12854] <= 15'b111100010111101;
		Coeff[12855] <= 15'b111100010111110;
		Coeff[12856] <= 15'b111100010111111;
		Coeff[12857] <= 15'b111100011000000;
		Coeff[12858] <= 15'b111100011000001;
		Coeff[12859] <= 15'b111100011000010;
		Coeff[12860] <= 15'b111100011000100;
		Coeff[12861] <= 15'b111100011000101;
		Coeff[12862] <= 15'b111100011000110;
		Coeff[12863] <= 15'b111100011000111;
		Coeff[12864] <= 15'b111100011001000;
		Coeff[12865] <= 15'b111100011001001;
		Coeff[12866] <= 15'b111100011001010;
		Coeff[12867] <= 15'b111100011001011;
		Coeff[12868] <= 15'b111100011001100;
		Coeff[12869] <= 15'b111100011001101;
		Coeff[12870] <= 15'b111100011001110;
		Coeff[12871] <= 15'b111100011001111;
		Coeff[12872] <= 15'b111100011010000;
		Coeff[12873] <= 15'b111100011010001;
		Coeff[12874] <= 15'b111100011010010;
		Coeff[12875] <= 15'b111100011010011;
		Coeff[12876] <= 15'b111100011010100;
		Coeff[12877] <= 15'b111100011010101;
		Coeff[12878] <= 15'b111100011010110;
		Coeff[12879] <= 15'b111100011010111;
		Coeff[12880] <= 15'b111100011011000;
		Coeff[12881] <= 15'b111100011011001;
		Coeff[12882] <= 15'b111100011011010;
		Coeff[12883] <= 15'b111100011011011;
		Coeff[12884] <= 15'b111100011011100;
		Coeff[12885] <= 15'b111100011011101;
		Coeff[12886] <= 15'b111100011011110;
		Coeff[12887] <= 15'b111100011100000;
		Coeff[12888] <= 15'b111100011100001;
		Coeff[12889] <= 15'b111100011100010;
		Coeff[12890] <= 15'b111100011100011;
		Coeff[12891] <= 15'b111100011100100;
		Coeff[12892] <= 15'b111100011100101;
		Coeff[12893] <= 15'b111100011100110;
		Coeff[12894] <= 15'b111100011100111;
		Coeff[12895] <= 15'b111100011101000;
		Coeff[12896] <= 15'b111100011101001;
		Coeff[12897] <= 15'b111100011101010;
		Coeff[12898] <= 15'b111100011101011;
		Coeff[12899] <= 15'b111100011101100;
		Coeff[12900] <= 15'b111100011101101;
		Coeff[12901] <= 15'b111100011101110;
		Coeff[12902] <= 15'b111100011101111;
		Coeff[12903] <= 15'b111100011110000;
		Coeff[12904] <= 15'b111100011110001;
		Coeff[12905] <= 15'b111100011110010;
		Coeff[12906] <= 15'b111100011110011;
		Coeff[12907] <= 15'b111100011110100;
		Coeff[12908] <= 15'b111100011110101;
		Coeff[12909] <= 15'b111100011110110;
		Coeff[12910] <= 15'b111100011110111;
		Coeff[12911] <= 15'b111100011111000;
		Coeff[12912] <= 15'b111100011111001;
		Coeff[12913] <= 15'b111100011111010;
		Coeff[12914] <= 15'b111100011111011;
		Coeff[12915] <= 15'b111100011111100;
		Coeff[12916] <= 15'b111100011111101;
		Coeff[12917] <= 15'b111100011111110;
		Coeff[12918] <= 15'b111100011111111;
		Coeff[12919] <= 15'b111100100000000;
		Coeff[12920] <= 15'b111100100000001;
		Coeff[12921] <= 15'b111100100000010;
		Coeff[12922] <= 15'b111100100000100;
		Coeff[12923] <= 15'b111100100000101;
		Coeff[12924] <= 15'b111100100000110;
		Coeff[12925] <= 15'b111100100000111;
		Coeff[12926] <= 15'b111100100001000;
		Coeff[12927] <= 15'b111100100001001;
		Coeff[12928] <= 15'b111100100001010;
		Coeff[12929] <= 15'b111100100001011;
		Coeff[12930] <= 15'b111100100001100;
		Coeff[12931] <= 15'b111100100001101;
		Coeff[12932] <= 15'b111100100001110;
		Coeff[12933] <= 15'b111100100001111;
		Coeff[12934] <= 15'b111100100010000;
		Coeff[12935] <= 15'b111100100010001;
		Coeff[12936] <= 15'b111100100010010;
		Coeff[12937] <= 15'b111100100010011;
		Coeff[12938] <= 15'b111100100010100;
		Coeff[12939] <= 15'b111100100010101;
		Coeff[12940] <= 15'b111100100010110;
		Coeff[12941] <= 15'b111100100010111;
		Coeff[12942] <= 15'b111100100011000;
		Coeff[12943] <= 15'b111100100011001;
		Coeff[12944] <= 15'b111100100011010;
		Coeff[12945] <= 15'b111100100011011;
		Coeff[12946] <= 15'b111100100011100;
		Coeff[12947] <= 15'b111100100011101;
		Coeff[12948] <= 15'b111100100011110;
		Coeff[12949] <= 15'b111100100011111;
		Coeff[12950] <= 15'b111100100100000;
		Coeff[12951] <= 15'b111100100100001;
		Coeff[12952] <= 15'b111100100100010;
		Coeff[12953] <= 15'b111100100100011;
		Coeff[12954] <= 15'b111100100100100;
		Coeff[12955] <= 15'b111100100100101;
		Coeff[12956] <= 15'b111100100100110;
		Coeff[12957] <= 15'b111100100100111;
		Coeff[12958] <= 15'b111100100101000;
		Coeff[12959] <= 15'b111100100101001;
		Coeff[12960] <= 15'b111100100101010;
		Coeff[12961] <= 15'b111100100101011;
		Coeff[12962] <= 15'b111100100101100;
		Coeff[12963] <= 15'b111100100101101;
		Coeff[12964] <= 15'b111100100101110;
		Coeff[12965] <= 15'b111100100101111;
		Coeff[12966] <= 15'b111100100110000;
		Coeff[12967] <= 15'b111100100110001;
		Coeff[12968] <= 15'b111100100110010;
		Coeff[12969] <= 15'b111100100110011;
		Coeff[12970] <= 15'b111100100110100;
		Coeff[12971] <= 15'b111100100110101;
		Coeff[12972] <= 15'b111100100110110;
		Coeff[12973] <= 15'b111100100110111;
		Coeff[12974] <= 15'b111100100111000;
		Coeff[12975] <= 15'b111100100111001;
		Coeff[12976] <= 15'b111100100111010;
		Coeff[12977] <= 15'b111100100111011;
		Coeff[12978] <= 15'b111100100111100;
		Coeff[12979] <= 15'b111100100111101;
		Coeff[12980] <= 15'b111100100111110;
		Coeff[12981] <= 15'b111100100111111;
		Coeff[12982] <= 15'b111100101000000;
		Coeff[12983] <= 15'b111100101000001;
		Coeff[12984] <= 15'b111100101000010;
		Coeff[12985] <= 15'b111100101000011;
		Coeff[12986] <= 15'b111100101000100;
		Coeff[12987] <= 15'b111100101000101;
		Coeff[12988] <= 15'b111100101000110;
		Coeff[12989] <= 15'b111100101000111;
		Coeff[12990] <= 15'b111100101001000;
		Coeff[12991] <= 15'b111100101001001;
		Coeff[12992] <= 15'b111100101001010;
		Coeff[12993] <= 15'b111100101001011;
		Coeff[12994] <= 15'b111100101001100;
		Coeff[12995] <= 15'b111100101001101;
		Coeff[12996] <= 15'b111100101001110;
		Coeff[12997] <= 15'b111100101001111;
		Coeff[12998] <= 15'b111100101010001;
		Coeff[12999] <= 15'b111100101010010;
		Coeff[13000] <= 15'b111100101010011;
		Coeff[13001] <= 15'b111100101010100;
		Coeff[13002] <= 15'b111100101010101;
		Coeff[13003] <= 15'b111100101010110;
		Coeff[13004] <= 15'b111100101010111;
		Coeff[13005] <= 15'b111100101011000;
		Coeff[13006] <= 15'b111100101011001;
		Coeff[13007] <= 15'b111100101011010;
		Coeff[13008] <= 15'b111100101011011;
		Coeff[13009] <= 15'b111100101011100;
		Coeff[13010] <= 15'b111100101011101;
		Coeff[13011] <= 15'b111100101011110;
		Coeff[13012] <= 15'b111100101011111;
		Coeff[13013] <= 15'b111100101100000;
		Coeff[13014] <= 15'b111100101100000;
		Coeff[13015] <= 15'b111100101100001;
		Coeff[13016] <= 15'b111100101100010;
		Coeff[13017] <= 15'b111100101100011;
		Coeff[13018] <= 15'b111100101100100;
		Coeff[13019] <= 15'b111100101100101;
		Coeff[13020] <= 15'b111100101100110;
		Coeff[13021] <= 15'b111100101100111;
		Coeff[13022] <= 15'b111100101101000;
		Coeff[13023] <= 15'b111100101101001;
		Coeff[13024] <= 15'b111100101101010;
		Coeff[13025] <= 15'b111100101101011;
		Coeff[13026] <= 15'b111100101101100;
		Coeff[13027] <= 15'b111100101101101;
		Coeff[13028] <= 15'b111100101101110;
		Coeff[13029] <= 15'b111100101101111;
		Coeff[13030] <= 15'b111100101110000;
		Coeff[13031] <= 15'b111100101110001;
		Coeff[13032] <= 15'b111100101110010;
		Coeff[13033] <= 15'b111100101110011;
		Coeff[13034] <= 15'b111100101110100;
		Coeff[13035] <= 15'b111100101110101;
		Coeff[13036] <= 15'b111100101110110;
		Coeff[13037] <= 15'b111100101110111;
		Coeff[13038] <= 15'b111100101111000;
		Coeff[13039] <= 15'b111100101111001;
		Coeff[13040] <= 15'b111100101111010;
		Coeff[13041] <= 15'b111100101111011;
		Coeff[13042] <= 15'b111100101111100;
		Coeff[13043] <= 15'b111100101111101;
		Coeff[13044] <= 15'b111100101111110;
		Coeff[13045] <= 15'b111100101111111;
		Coeff[13046] <= 15'b111100110000000;
		Coeff[13047] <= 15'b111100110000001;
		Coeff[13048] <= 15'b111100110000010;
		Coeff[13049] <= 15'b111100110000011;
		Coeff[13050] <= 15'b111100110000100;
		Coeff[13051] <= 15'b111100110000101;
		Coeff[13052] <= 15'b111100110000110;
		Coeff[13053] <= 15'b111100110000111;
		Coeff[13054] <= 15'b111100110001000;
		Coeff[13055] <= 15'b111100110001001;
		Coeff[13056] <= 15'b111100110001010;
		Coeff[13057] <= 15'b111100110001011;
		Coeff[13058] <= 15'b111100110001100;
		Coeff[13059] <= 15'b111100110001101;
		Coeff[13060] <= 15'b111100110001110;
		Coeff[13061] <= 15'b111100110001111;
		Coeff[13062] <= 15'b111100110010000;
		Coeff[13063] <= 15'b111100110010001;
		Coeff[13064] <= 15'b111100110010010;
		Coeff[13065] <= 15'b111100110010011;
		Coeff[13066] <= 15'b111100110010100;
		Coeff[13067] <= 15'b111100110010101;
		Coeff[13068] <= 15'b111100110010110;
		Coeff[13069] <= 15'b111100110010111;
		Coeff[13070] <= 15'b111100110011000;
		Coeff[13071] <= 15'b111100110011001;
		Coeff[13072] <= 15'b111100110011010;
		Coeff[13073] <= 15'b111100110011011;
		Coeff[13074] <= 15'b111100110011100;
		Coeff[13075] <= 15'b111100110011101;
		Coeff[13076] <= 15'b111100110011110;
		Coeff[13077] <= 15'b111100110011111;
		Coeff[13078] <= 15'b111100110100000;
		Coeff[13079] <= 15'b111100110100001;
		Coeff[13080] <= 15'b111100110100010;
		Coeff[13081] <= 15'b111100110100011;
		Coeff[13082] <= 15'b111100110100100;
		Coeff[13083] <= 15'b111100110100101;
		Coeff[13084] <= 15'b111100110100110;
		Coeff[13085] <= 15'b111100110100111;
		Coeff[13086] <= 15'b111100110101000;
		Coeff[13087] <= 15'b111100110101001;
		Coeff[13088] <= 15'b111100110101010;
		Coeff[13089] <= 15'b111100110101011;
		Coeff[13090] <= 15'b111100110101011;
		Coeff[13091] <= 15'b111100110101100;
		Coeff[13092] <= 15'b111100110101101;
		Coeff[13093] <= 15'b111100110101110;
		Coeff[13094] <= 15'b111100110101111;
		Coeff[13095] <= 15'b111100110110000;
		Coeff[13096] <= 15'b111100110110001;
		Coeff[13097] <= 15'b111100110110010;
		Coeff[13098] <= 15'b111100110110011;
		Coeff[13099] <= 15'b111100110110100;
		Coeff[13100] <= 15'b111100110110101;
		Coeff[13101] <= 15'b111100110110110;
		Coeff[13102] <= 15'b111100110110111;
		Coeff[13103] <= 15'b111100110111000;
		Coeff[13104] <= 15'b111100110111001;
		Coeff[13105] <= 15'b111100110111010;
		Coeff[13106] <= 15'b111100110111011;
		Coeff[13107] <= 15'b111100110111100;
		Coeff[13108] <= 15'b111100110111101;
		Coeff[13109] <= 15'b111100110111110;
		Coeff[13110] <= 15'b111100110111111;
		Coeff[13111] <= 15'b111100111000000;
		Coeff[13112] <= 15'b111100111000001;
		Coeff[13113] <= 15'b111100111000010;
		Coeff[13114] <= 15'b111100111000011;
		Coeff[13115] <= 15'b111100111000100;
		Coeff[13116] <= 15'b111100111000101;
		Coeff[13117] <= 15'b111100111000110;
		Coeff[13118] <= 15'b111100111000111;
		Coeff[13119] <= 15'b111100111001000;
		Coeff[13120] <= 15'b111100111001001;
		Coeff[13121] <= 15'b111100111001010;
		Coeff[13122] <= 15'b111100111001011;
		Coeff[13123] <= 15'b111100111001100;
		Coeff[13124] <= 15'b111100111001100;
		Coeff[13125] <= 15'b111100111001101;
		Coeff[13126] <= 15'b111100111001110;
		Coeff[13127] <= 15'b111100111001111;
		Coeff[13128] <= 15'b111100111010000;
		Coeff[13129] <= 15'b111100111010001;
		Coeff[13130] <= 15'b111100111010010;
		Coeff[13131] <= 15'b111100111010011;
		Coeff[13132] <= 15'b111100111010100;
		Coeff[13133] <= 15'b111100111010101;
		Coeff[13134] <= 15'b111100111010110;
		Coeff[13135] <= 15'b111100111010111;
		Coeff[13136] <= 15'b111100111011000;
		Coeff[13137] <= 15'b111100111011001;
		Coeff[13138] <= 15'b111100111011010;
		Coeff[13139] <= 15'b111100111011011;
		Coeff[13140] <= 15'b111100111011100;
		Coeff[13141] <= 15'b111100111011101;
		Coeff[13142] <= 15'b111100111011110;
		Coeff[13143] <= 15'b111100111011111;
		Coeff[13144] <= 15'b111100111100000;
		Coeff[13145] <= 15'b111100111100001;
		Coeff[13146] <= 15'b111100111100010;
		Coeff[13147] <= 15'b111100111100011;
		Coeff[13148] <= 15'b111100111100100;
		Coeff[13149] <= 15'b111100111100101;
		Coeff[13150] <= 15'b111100111100110;
		Coeff[13151] <= 15'b111100111100110;
		Coeff[13152] <= 15'b111100111100111;
		Coeff[13153] <= 15'b111100111101000;
		Coeff[13154] <= 15'b111100111101001;
		Coeff[13155] <= 15'b111100111101010;
		Coeff[13156] <= 15'b111100111101011;
		Coeff[13157] <= 15'b111100111101100;
		Coeff[13158] <= 15'b111100111101101;
		Coeff[13159] <= 15'b111100111101110;
		Coeff[13160] <= 15'b111100111101111;
		Coeff[13161] <= 15'b111100111110000;
		Coeff[13162] <= 15'b111100111110001;
		Coeff[13163] <= 15'b111100111110010;
		Coeff[13164] <= 15'b111100111110011;
		Coeff[13165] <= 15'b111100111110100;
		Coeff[13166] <= 15'b111100111110101;
		Coeff[13167] <= 15'b111100111110110;
		Coeff[13168] <= 15'b111100111110111;
		Coeff[13169] <= 15'b111100111111000;
		Coeff[13170] <= 15'b111100111111001;
		Coeff[13171] <= 15'b111100111111010;
		Coeff[13172] <= 15'b111100111111011;
		Coeff[13173] <= 15'b111100111111011;
		Coeff[13174] <= 15'b111100111111100;
		Coeff[13175] <= 15'b111100111111101;
		Coeff[13176] <= 15'b111100111111110;
		Coeff[13177] <= 15'b111100111111111;
		Coeff[13178] <= 15'b111101000000000;
		Coeff[13179] <= 15'b111101000000001;
		Coeff[13180] <= 15'b111101000000010;
		Coeff[13181] <= 15'b111101000000011;
		Coeff[13182] <= 15'b111101000000100;
		Coeff[13183] <= 15'b111101000000101;
		Coeff[13184] <= 15'b111101000000110;
		Coeff[13185] <= 15'b111101000000111;
		Coeff[13186] <= 15'b111101000001000;
		Coeff[13187] <= 15'b111101000001001;
		Coeff[13188] <= 15'b111101000001010;
		Coeff[13189] <= 15'b111101000001011;
		Coeff[13190] <= 15'b111101000001100;
		Coeff[13191] <= 15'b111101000001101;
		Coeff[13192] <= 15'b111101000001110;
		Coeff[13193] <= 15'b111101000001110;
		Coeff[13194] <= 15'b111101000001111;
		Coeff[13195] <= 15'b111101000010000;
		Coeff[13196] <= 15'b111101000010001;
		Coeff[13197] <= 15'b111101000010010;
		Coeff[13198] <= 15'b111101000010011;
		Coeff[13199] <= 15'b111101000010100;
		Coeff[13200] <= 15'b111101000010101;
		Coeff[13201] <= 15'b111101000010110;
		Coeff[13202] <= 15'b111101000010111;
		Coeff[13203] <= 15'b111101000011000;
		Coeff[13204] <= 15'b111101000011001;
		Coeff[13205] <= 15'b111101000011010;
		Coeff[13206] <= 15'b111101000011011;
		Coeff[13207] <= 15'b111101000011100;
		Coeff[13208] <= 15'b111101000011101;
		Coeff[13209] <= 15'b111101000011110;
		Coeff[13210] <= 15'b111101000011111;
		Coeff[13211] <= 15'b111101000011111;
		Coeff[13212] <= 15'b111101000100000;
		Coeff[13213] <= 15'b111101000100001;
		Coeff[13214] <= 15'b111101000100010;
		Coeff[13215] <= 15'b111101000100011;
		Coeff[13216] <= 15'b111101000100100;
		Coeff[13217] <= 15'b111101000100101;
		Coeff[13218] <= 15'b111101000100110;
		Coeff[13219] <= 15'b111101000100111;
		Coeff[13220] <= 15'b111101000101000;
		Coeff[13221] <= 15'b111101000101001;
		Coeff[13222] <= 15'b111101000101010;
		Coeff[13223] <= 15'b111101000101011;
		Coeff[13224] <= 15'b111101000101100;
		Coeff[13225] <= 15'b111101000101101;
		Coeff[13226] <= 15'b111101000101110;
		Coeff[13227] <= 15'b111101000101110;
		Coeff[13228] <= 15'b111101000101111;
		Coeff[13229] <= 15'b111101000110000;
		Coeff[13230] <= 15'b111101000110001;
		Coeff[13231] <= 15'b111101000110010;
		Coeff[13232] <= 15'b111101000110011;
		Coeff[13233] <= 15'b111101000110100;
		Coeff[13234] <= 15'b111101000110101;
		Coeff[13235] <= 15'b111101000110110;
		Coeff[13236] <= 15'b111101000110111;
		Coeff[13237] <= 15'b111101000111000;
		Coeff[13238] <= 15'b111101000111001;
		Coeff[13239] <= 15'b111101000111010;
		Coeff[13240] <= 15'b111101000111011;
		Coeff[13241] <= 15'b111101000111100;
		Coeff[13242] <= 15'b111101000111100;
		Coeff[13243] <= 15'b111101000111101;
		Coeff[13244] <= 15'b111101000111110;
		Coeff[13245] <= 15'b111101000111111;
		Coeff[13246] <= 15'b111101001000000;
		Coeff[13247] <= 15'b111101001000001;
		Coeff[13248] <= 15'b111101001000010;
		Coeff[13249] <= 15'b111101001000011;
		Coeff[13250] <= 15'b111101001000100;
		Coeff[13251] <= 15'b111101001000101;
		Coeff[13252] <= 15'b111101001000110;
		Coeff[13253] <= 15'b111101001000111;
		Coeff[13254] <= 15'b111101001001000;
		Coeff[13255] <= 15'b111101001001001;
		Coeff[13256] <= 15'b111101001001001;
		Coeff[13257] <= 15'b111101001001010;
		Coeff[13258] <= 15'b111101001001011;
		Coeff[13259] <= 15'b111101001001100;
		Coeff[13260] <= 15'b111101001001101;
		Coeff[13261] <= 15'b111101001001110;
		Coeff[13262] <= 15'b111101001001111;
		Coeff[13263] <= 15'b111101001010000;
		Coeff[13264] <= 15'b111101001010001;
		Coeff[13265] <= 15'b111101001010010;
		Coeff[13266] <= 15'b111101001010011;
		Coeff[13267] <= 15'b111101001010100;
		Coeff[13268] <= 15'b111101001010101;
		Coeff[13269] <= 15'b111101001010110;
		Coeff[13270] <= 15'b111101001010110;
		Coeff[13271] <= 15'b111101001010111;
		Coeff[13272] <= 15'b111101001011000;
		Coeff[13273] <= 15'b111101001011001;
		Coeff[13274] <= 15'b111101001011010;
		Coeff[13275] <= 15'b111101001011011;
		Coeff[13276] <= 15'b111101001011100;
		Coeff[13277] <= 15'b111101001011101;
		Coeff[13278] <= 15'b111101001011110;
		Coeff[13279] <= 15'b111101001011111;
		Coeff[13280] <= 15'b111101001100000;
		Coeff[13281] <= 15'b111101001100001;
		Coeff[13282] <= 15'b111101001100010;
		Coeff[13283] <= 15'b111101001100010;
		Coeff[13284] <= 15'b111101001100011;
		Coeff[13285] <= 15'b111101001100100;
		Coeff[13286] <= 15'b111101001100101;
		Coeff[13287] <= 15'b111101001100110;
		Coeff[13288] <= 15'b111101001100111;
		Coeff[13289] <= 15'b111101001101000;
		Coeff[13290] <= 15'b111101001101001;
		Coeff[13291] <= 15'b111101001101010;
		Coeff[13292] <= 15'b111101001101011;
		Coeff[13293] <= 15'b111101001101100;
		Coeff[13294] <= 15'b111101001101101;
		Coeff[13295] <= 15'b111101001101101;
		Coeff[13296] <= 15'b111101001101110;
		Coeff[13297] <= 15'b111101001101111;
		Coeff[13298] <= 15'b111101001110000;
		Coeff[13299] <= 15'b111101001110001;
		Coeff[13300] <= 15'b111101001110010;
		Coeff[13301] <= 15'b111101001110011;
		Coeff[13302] <= 15'b111101001110100;
		Coeff[13303] <= 15'b111101001110101;
		Coeff[13304] <= 15'b111101001110110;
		Coeff[13305] <= 15'b111101001110111;
		Coeff[13306] <= 15'b111101001111000;
		Coeff[13307] <= 15'b111101001111000;
		Coeff[13308] <= 15'b111101001111001;
		Coeff[13309] <= 15'b111101001111010;
		Coeff[13310] <= 15'b111101001111011;
		Coeff[13311] <= 15'b111101001111100;
		Coeff[13312] <= 15'b111101001111101;
		Coeff[13313] <= 15'b111101001111110;
		Coeff[13314] <= 15'b111101001111111;
		Coeff[13315] <= 15'b111101010000000;
		Coeff[13316] <= 15'b111101010000001;
		Coeff[13317] <= 15'b111101010000010;
		Coeff[13318] <= 15'b111101010000010;
		Coeff[13319] <= 15'b111101010000011;
		Coeff[13320] <= 15'b111101010000100;
		Coeff[13321] <= 15'b111101010000101;
		Coeff[13322] <= 15'b111101010000110;
		Coeff[13323] <= 15'b111101010000111;
		Coeff[13324] <= 15'b111101010001000;
		Coeff[13325] <= 15'b111101010001001;
		Coeff[13326] <= 15'b111101010001010;
		Coeff[13327] <= 15'b111101010001011;
		Coeff[13328] <= 15'b111101010001100;
		Coeff[13329] <= 15'b111101010001100;
		Coeff[13330] <= 15'b111101010001101;
		Coeff[13331] <= 15'b111101010001110;
		Coeff[13332] <= 15'b111101010001111;
		Coeff[13333] <= 15'b111101010010000;
		Coeff[13334] <= 15'b111101010010001;
		Coeff[13335] <= 15'b111101010010010;
		Coeff[13336] <= 15'b111101010010011;
		Coeff[13337] <= 15'b111101010010100;
		Coeff[13338] <= 15'b111101010010101;
		Coeff[13339] <= 15'b111101010010110;
		Coeff[13340] <= 15'b111101010010110;
		Coeff[13341] <= 15'b111101010010111;
		Coeff[13342] <= 15'b111101010011000;
		Coeff[13343] <= 15'b111101010011001;
		Coeff[13344] <= 15'b111101010011010;
		Coeff[13345] <= 15'b111101010011011;
		Coeff[13346] <= 15'b111101010011100;
		Coeff[13347] <= 15'b111101010011101;
		Coeff[13348] <= 15'b111101010011110;
		Coeff[13349] <= 15'b111101010011111;
		Coeff[13350] <= 15'b111101010011111;
		Coeff[13351] <= 15'b111101010100000;
		Coeff[13352] <= 15'b111101010100001;
		Coeff[13353] <= 15'b111101010100010;
		Coeff[13354] <= 15'b111101010100011;
		Coeff[13355] <= 15'b111101010100100;
		Coeff[13356] <= 15'b111101010100101;
		Coeff[13357] <= 15'b111101010100110;
		Coeff[13358] <= 15'b111101010100111;
		Coeff[13359] <= 15'b111101010101000;
		Coeff[13360] <= 15'b111101010101000;
		Coeff[13361] <= 15'b111101010101001;
		Coeff[13362] <= 15'b111101010101010;
		Coeff[13363] <= 15'b111101010101011;
		Coeff[13364] <= 15'b111101010101100;
		Coeff[13365] <= 15'b111101010101101;
		Coeff[13366] <= 15'b111101010101110;
		Coeff[13367] <= 15'b111101010101111;
		Coeff[13368] <= 15'b111101010110000;
		Coeff[13369] <= 15'b111101010110001;
		Coeff[13370] <= 15'b111101010110001;
		Coeff[13371] <= 15'b111101010110010;
		Coeff[13372] <= 15'b111101010110011;
		Coeff[13373] <= 15'b111101010110100;
		Coeff[13374] <= 15'b111101010110101;
		Coeff[13375] <= 15'b111101010110110;
		Coeff[13376] <= 15'b111101010110111;
		Coeff[13377] <= 15'b111101010111000;
		Coeff[13378] <= 15'b111101010111001;
		Coeff[13379] <= 15'b111101010111001;
		Coeff[13380] <= 15'b111101010111010;
		Coeff[13381] <= 15'b111101010111011;
		Coeff[13382] <= 15'b111101010111100;
		Coeff[13383] <= 15'b111101010111101;
		Coeff[13384] <= 15'b111101010111110;
		Coeff[13385] <= 15'b111101010111111;
		Coeff[13386] <= 15'b111101011000000;
		Coeff[13387] <= 15'b111101011000001;
		Coeff[13388] <= 15'b111101011000001;
		Coeff[13389] <= 15'b111101011000010;
		Coeff[13390] <= 15'b111101011000011;
		Coeff[13391] <= 15'b111101011000100;
		Coeff[13392] <= 15'b111101011000101;
		Coeff[13393] <= 15'b111101011000110;
		Coeff[13394] <= 15'b111101011000111;
		Coeff[13395] <= 15'b111101011001000;
		Coeff[13396] <= 15'b111101011001001;
		Coeff[13397] <= 15'b111101011001001;
		Coeff[13398] <= 15'b111101011001010;
		Coeff[13399] <= 15'b111101011001011;
		Coeff[13400] <= 15'b111101011001100;
		Coeff[13401] <= 15'b111101011001101;
		Coeff[13402] <= 15'b111101011001110;
		Coeff[13403] <= 15'b111101011001111;
		Coeff[13404] <= 15'b111101011010000;
		Coeff[13405] <= 15'b111101011010001;
		Coeff[13406] <= 15'b111101011010001;
		Coeff[13407] <= 15'b111101011010010;
		Coeff[13408] <= 15'b111101011010011;
		Coeff[13409] <= 15'b111101011010100;
		Coeff[13410] <= 15'b111101011010101;
		Coeff[13411] <= 15'b111101011010110;
		Coeff[13412] <= 15'b111101011010111;
		Coeff[13413] <= 15'b111101011011000;
		Coeff[13414] <= 15'b111101011011001;
		Coeff[13415] <= 15'b111101011011001;
		Coeff[13416] <= 15'b111101011011010;
		Coeff[13417] <= 15'b111101011011011;
		Coeff[13418] <= 15'b111101011011100;
		Coeff[13419] <= 15'b111101011011101;
		Coeff[13420] <= 15'b111101011011110;
		Coeff[13421] <= 15'b111101011011111;
		Coeff[13422] <= 15'b111101011100000;
		Coeff[13423] <= 15'b111101011100000;
		Coeff[13424] <= 15'b111101011100001;
		Coeff[13425] <= 15'b111101011100010;
		Coeff[13426] <= 15'b111101011100011;
		Coeff[13427] <= 15'b111101011100100;
		Coeff[13428] <= 15'b111101011100101;
		Coeff[13429] <= 15'b111101011100110;
		Coeff[13430] <= 15'b111101011100111;
		Coeff[13431] <= 15'b111101011101000;
		Coeff[13432] <= 15'b111101011101000;
		Coeff[13433] <= 15'b111101011101001;
		Coeff[13434] <= 15'b111101011101010;
		Coeff[13435] <= 15'b111101011101011;
		Coeff[13436] <= 15'b111101011101100;
		Coeff[13437] <= 15'b111101011101101;
		Coeff[13438] <= 15'b111101011101110;
		Coeff[13439] <= 15'b111101011101111;
		Coeff[13440] <= 15'b111101011101111;
		Coeff[13441] <= 15'b111101011110000;
		Coeff[13442] <= 15'b111101011110001;
		Coeff[13443] <= 15'b111101011110010;
		Coeff[13444] <= 15'b111101011110011;
		Coeff[13445] <= 15'b111101011110100;
		Coeff[13446] <= 15'b111101011110101;
		Coeff[13447] <= 15'b111101011110110;
		Coeff[13448] <= 15'b111101011110110;
		Coeff[13449] <= 15'b111101011110111;
		Coeff[13450] <= 15'b111101011111000;
		Coeff[13451] <= 15'b111101011111001;
		Coeff[13452] <= 15'b111101011111010;
		Coeff[13453] <= 15'b111101011111011;
		Coeff[13454] <= 15'b111101011111100;
		Coeff[13455] <= 15'b111101011111100;
		Coeff[13456] <= 15'b111101011111101;
		Coeff[13457] <= 15'b111101011111110;
		Coeff[13458] <= 15'b111101011111111;
		Coeff[13459] <= 15'b111101100000000;
		Coeff[13460] <= 15'b111101100000001;
		Coeff[13461] <= 15'b111101100000010;
		Coeff[13462] <= 15'b111101100000011;
		Coeff[13463] <= 15'b111101100000011;
		Coeff[13464] <= 15'b111101100000100;
		Coeff[13465] <= 15'b111101100000101;
		Coeff[13466] <= 15'b111101100000110;
		Coeff[13467] <= 15'b111101100000111;
		Coeff[13468] <= 15'b111101100001000;
		Coeff[13469] <= 15'b111101100001001;
		Coeff[13470] <= 15'b111101100001010;
		Coeff[13471] <= 15'b111101100001010;
		Coeff[13472] <= 15'b111101100001011;
		Coeff[13473] <= 15'b111101100001100;
		Coeff[13474] <= 15'b111101100001101;
		Coeff[13475] <= 15'b111101100001110;
		Coeff[13476] <= 15'b111101100001111;
		Coeff[13477] <= 15'b111101100010000;
		Coeff[13478] <= 15'b111101100010000;
		Coeff[13479] <= 15'b111101100010001;
		Coeff[13480] <= 15'b111101100010010;
		Coeff[13481] <= 15'b111101100010011;
		Coeff[13482] <= 15'b111101100010100;
		Coeff[13483] <= 15'b111101100010101;
		Coeff[13484] <= 15'b111101100010110;
		Coeff[13485] <= 15'b111101100010110;
		Coeff[13486] <= 15'b111101100010111;
		Coeff[13487] <= 15'b111101100011000;
		Coeff[13488] <= 15'b111101100011001;
		Coeff[13489] <= 15'b111101100011010;
		Coeff[13490] <= 15'b111101100011011;
		Coeff[13491] <= 15'b111101100011100;
		Coeff[13492] <= 15'b111101100011100;
		Coeff[13493] <= 15'b111101100011101;
		Coeff[13494] <= 15'b111101100011110;
		Coeff[13495] <= 15'b111101100011111;
		Coeff[13496] <= 15'b111101100100000;
		Coeff[13497] <= 15'b111101100100001;
		Coeff[13498] <= 15'b111101100100010;
		Coeff[13499] <= 15'b111101100100011;
		Coeff[13500] <= 15'b111101100100011;
		Coeff[13501] <= 15'b111101100100100;
		Coeff[13502] <= 15'b111101100100101;
		Coeff[13503] <= 15'b111101100100110;
		Coeff[13504] <= 15'b111101100100111;
		Coeff[13505] <= 15'b111101100101000;
		Coeff[13506] <= 15'b111101100101001;
		Coeff[13507] <= 15'b111101100101001;
		Coeff[13508] <= 15'b111101100101010;
		Coeff[13509] <= 15'b111101100101011;
		Coeff[13510] <= 15'b111101100101100;
		Coeff[13511] <= 15'b111101100101101;
		Coeff[13512] <= 15'b111101100101110;
		Coeff[13513] <= 15'b111101100101110;
		Coeff[13514] <= 15'b111101100101111;
		Coeff[13515] <= 15'b111101100110000;
		Coeff[13516] <= 15'b111101100110001;
		Coeff[13517] <= 15'b111101100110010;
		Coeff[13518] <= 15'b111101100110011;
		Coeff[13519] <= 15'b111101100110100;
		Coeff[13520] <= 15'b111101100110100;
		Coeff[13521] <= 15'b111101100110101;
		Coeff[13522] <= 15'b111101100110110;
		Coeff[13523] <= 15'b111101100110111;
		Coeff[13524] <= 15'b111101100111000;
		Coeff[13525] <= 15'b111101100111001;
		Coeff[13526] <= 15'b111101100111010;
		Coeff[13527] <= 15'b111101100111010;
		Coeff[13528] <= 15'b111101100111011;
		Coeff[13529] <= 15'b111101100111100;
		Coeff[13530] <= 15'b111101100111101;
		Coeff[13531] <= 15'b111101100111110;
		Coeff[13532] <= 15'b111101100111111;
		Coeff[13533] <= 15'b111101101000000;
		Coeff[13534] <= 15'b111101101000000;
		Coeff[13535] <= 15'b111101101000001;
		Coeff[13536] <= 15'b111101101000010;
		Coeff[13537] <= 15'b111101101000011;
		Coeff[13538] <= 15'b111101101000100;
		Coeff[13539] <= 15'b111101101000101;
		Coeff[13540] <= 15'b111101101000101;
		Coeff[13541] <= 15'b111101101000110;
		Coeff[13542] <= 15'b111101101000111;
		Coeff[13543] <= 15'b111101101001000;
		Coeff[13544] <= 15'b111101101001001;
		Coeff[13545] <= 15'b111101101001010;
		Coeff[13546] <= 15'b111101101001011;
		Coeff[13547] <= 15'b111101101001011;
		Coeff[13548] <= 15'b111101101001100;
		Coeff[13549] <= 15'b111101101001101;
		Coeff[13550] <= 15'b111101101001110;
		Coeff[13551] <= 15'b111101101001111;
		Coeff[13552] <= 15'b111101101010000;
		Coeff[13553] <= 15'b111101101010000;
		Coeff[13554] <= 15'b111101101010001;
		Coeff[13555] <= 15'b111101101010010;
		Coeff[13556] <= 15'b111101101010011;
		Coeff[13557] <= 15'b111101101010100;
		Coeff[13558] <= 15'b111101101010101;
		Coeff[13559] <= 15'b111101101010101;
		Coeff[13560] <= 15'b111101101010110;
		Coeff[13561] <= 15'b111101101010111;
		Coeff[13562] <= 15'b111101101011000;
		Coeff[13563] <= 15'b111101101011001;
		Coeff[13564] <= 15'b111101101011010;
		Coeff[13565] <= 15'b111101101011010;
		Coeff[13566] <= 15'b111101101011011;
		Coeff[13567] <= 15'b111101101011100;
		Coeff[13568] <= 15'b111101101011101;
		Coeff[13569] <= 15'b111101101011110;
		Coeff[13570] <= 15'b111101101011111;
		Coeff[13571] <= 15'b111101101100000;
		Coeff[13572] <= 15'b111101101100000;
		Coeff[13573] <= 15'b111101101100001;
		Coeff[13574] <= 15'b111101101100010;
		Coeff[13575] <= 15'b111101101100011;
		Coeff[13576] <= 15'b111101101100100;
		Coeff[13577] <= 15'b111101101100101;
		Coeff[13578] <= 15'b111101101100101;
		Coeff[13579] <= 15'b111101101100110;
		Coeff[13580] <= 15'b111101101100111;
		Coeff[13581] <= 15'b111101101101000;
		Coeff[13582] <= 15'b111101101101001;
		Coeff[13583] <= 15'b111101101101010;
		Coeff[13584] <= 15'b111101101101010;
		Coeff[13585] <= 15'b111101101101011;
		Coeff[13586] <= 15'b111101101101100;
		Coeff[13587] <= 15'b111101101101101;
		Coeff[13588] <= 15'b111101101101110;
		Coeff[13589] <= 15'b111101101101111;
		Coeff[13590] <= 15'b111101101101111;
		Coeff[13591] <= 15'b111101101110000;
		Coeff[13592] <= 15'b111101101110001;
		Coeff[13593] <= 15'b111101101110010;
		Coeff[13594] <= 15'b111101101110011;
		Coeff[13595] <= 15'b111101101110100;
		Coeff[13596] <= 15'b111101101110100;
		Coeff[13597] <= 15'b111101101110101;
		Coeff[13598] <= 15'b111101101110110;
		Coeff[13599] <= 15'b111101101110111;
		Coeff[13600] <= 15'b111101101111000;
		Coeff[13601] <= 15'b111101101111001;
		Coeff[13602] <= 15'b111101101111001;
		Coeff[13603] <= 15'b111101101111010;
		Coeff[13604] <= 15'b111101101111011;
		Coeff[13605] <= 15'b111101101111100;
		Coeff[13606] <= 15'b111101101111101;
		Coeff[13607] <= 15'b111101101111101;
		Coeff[13608] <= 15'b111101101111110;
		Coeff[13609] <= 15'b111101101111111;
		Coeff[13610] <= 15'b111101110000000;
		Coeff[13611] <= 15'b111101110000001;
		Coeff[13612] <= 15'b111101110000010;
		Coeff[13613] <= 15'b111101110000010;
		Coeff[13614] <= 15'b111101110000011;
		Coeff[13615] <= 15'b111101110000100;
		Coeff[13616] <= 15'b111101110000101;
		Coeff[13617] <= 15'b111101110000110;
		Coeff[13618] <= 15'b111101110000111;
		Coeff[13619] <= 15'b111101110000111;
		Coeff[13620] <= 15'b111101110001000;
		Coeff[13621] <= 15'b111101110001001;
		Coeff[13622] <= 15'b111101110001010;
		Coeff[13623] <= 15'b111101110001011;
		Coeff[13624] <= 15'b111101110001011;
		Coeff[13625] <= 15'b111101110001100;
		Coeff[13626] <= 15'b111101110001101;
		Coeff[13627] <= 15'b111101110001110;
		Coeff[13628] <= 15'b111101110001111;
		Coeff[13629] <= 15'b111101110010000;
		Coeff[13630] <= 15'b111101110010000;
		Coeff[13631] <= 15'b111101110010001;
		Coeff[13632] <= 15'b111101110010010;
		Coeff[13633] <= 15'b111101110010011;
		Coeff[13634] <= 15'b111101110010100;
		Coeff[13635] <= 15'b111101110010101;
		Coeff[13636] <= 15'b111101110010101;
		Coeff[13637] <= 15'b111101110010110;
		Coeff[13638] <= 15'b111101110010111;
		Coeff[13639] <= 15'b111101110011000;
		Coeff[13640] <= 15'b111101110011001;
		Coeff[13641] <= 15'b111101110011001;
		Coeff[13642] <= 15'b111101110011010;
		Coeff[13643] <= 15'b111101110011011;
		Coeff[13644] <= 15'b111101110011100;
		Coeff[13645] <= 15'b111101110011101;
		Coeff[13646] <= 15'b111101110011101;
		Coeff[13647] <= 15'b111101110011110;
		Coeff[13648] <= 15'b111101110011111;
		Coeff[13649] <= 15'b111101110100000;
		Coeff[13650] <= 15'b111101110100001;
		Coeff[13651] <= 15'b111101110100010;
		Coeff[13652] <= 15'b111101110100010;
		Coeff[13653] <= 15'b111101110100011;
		Coeff[13654] <= 15'b111101110100100;
		Coeff[13655] <= 15'b111101110100101;
		Coeff[13656] <= 15'b111101110100110;
		Coeff[13657] <= 15'b111101110100110;
		Coeff[13658] <= 15'b111101110100111;
		Coeff[13659] <= 15'b111101110101000;
		Coeff[13660] <= 15'b111101110101001;
		Coeff[13661] <= 15'b111101110101010;
		Coeff[13662] <= 15'b111101110101010;
		Coeff[13663] <= 15'b111101110101011;
		Coeff[13664] <= 15'b111101110101100;
		Coeff[13665] <= 15'b111101110101101;
		Coeff[13666] <= 15'b111101110101110;
		Coeff[13667] <= 15'b111101110101111;
		Coeff[13668] <= 15'b111101110101111;
		Coeff[13669] <= 15'b111101110110000;
		Coeff[13670] <= 15'b111101110110001;
		Coeff[13671] <= 15'b111101110110010;
		Coeff[13672] <= 15'b111101110110011;
		Coeff[13673] <= 15'b111101110110011;
		Coeff[13674] <= 15'b111101110110100;
		Coeff[13675] <= 15'b111101110110101;
		Coeff[13676] <= 15'b111101110110110;
		Coeff[13677] <= 15'b111101110110111;
		Coeff[13678] <= 15'b111101110110111;
		Coeff[13679] <= 15'b111101110111000;
		Coeff[13680] <= 15'b111101110111001;
		Coeff[13681] <= 15'b111101110111010;
		Coeff[13682] <= 15'b111101110111011;
		Coeff[13683] <= 15'b111101110111011;
		Coeff[13684] <= 15'b111101110111100;
		Coeff[13685] <= 15'b111101110111101;
		Coeff[13686] <= 15'b111101110111110;
		Coeff[13687] <= 15'b111101110111111;
		Coeff[13688] <= 15'b111101110111111;
		Coeff[13689] <= 15'b111101111000000;
		Coeff[13690] <= 15'b111101111000001;
		Coeff[13691] <= 15'b111101111000010;
		Coeff[13692] <= 15'b111101111000011;
		Coeff[13693] <= 15'b111101111000011;
		Coeff[13694] <= 15'b111101111000100;
		Coeff[13695] <= 15'b111101111000101;
		Coeff[13696] <= 15'b111101111000110;
		Coeff[13697] <= 15'b111101111000111;
		Coeff[13698] <= 15'b111101111000111;
		Coeff[13699] <= 15'b111101111001000;
		Coeff[13700] <= 15'b111101111001001;
		Coeff[13701] <= 15'b111101111001010;
		Coeff[13702] <= 15'b111101111001011;
		Coeff[13703] <= 15'b111101111001011;
		Coeff[13704] <= 15'b111101111001100;
		Coeff[13705] <= 15'b111101111001101;
		Coeff[13706] <= 15'b111101111001110;
		Coeff[13707] <= 15'b111101111001111;
		Coeff[13708] <= 15'b111101111001111;
		Coeff[13709] <= 15'b111101111010000;
		Coeff[13710] <= 15'b111101111010001;
		Coeff[13711] <= 15'b111101111010010;
		Coeff[13712] <= 15'b111101111010011;
		Coeff[13713] <= 15'b111101111010011;
		Coeff[13714] <= 15'b111101111010100;
		Coeff[13715] <= 15'b111101111010101;
		Coeff[13716] <= 15'b111101111010110;
		Coeff[13717] <= 15'b111101111010111;
		Coeff[13718] <= 15'b111101111010111;
		Coeff[13719] <= 15'b111101111011000;
		Coeff[13720] <= 15'b111101111011001;
		Coeff[13721] <= 15'b111101111011010;
		Coeff[13722] <= 15'b111101111011011;
		Coeff[13723] <= 15'b111101111011011;
		Coeff[13724] <= 15'b111101111011100;
		Coeff[13725] <= 15'b111101111011101;
		Coeff[13726] <= 15'b111101111011110;
		Coeff[13727] <= 15'b111101111011111;
		Coeff[13728] <= 15'b111101111011111;
		Coeff[13729] <= 15'b111101111100000;
		Coeff[13730] <= 15'b111101111100001;
		Coeff[13731] <= 15'b111101111100010;
		Coeff[13732] <= 15'b111101111100011;
		Coeff[13733] <= 15'b111101111100011;
		Coeff[13734] <= 15'b111101111100100;
		Coeff[13735] <= 15'b111101111100101;
		Coeff[13736] <= 15'b111101111100110;
		Coeff[13737] <= 15'b111101111100110;
		Coeff[13738] <= 15'b111101111100111;
		Coeff[13739] <= 15'b111101111101000;
		Coeff[13740] <= 15'b111101111101001;
		Coeff[13741] <= 15'b111101111101010;
		Coeff[13742] <= 15'b111101111101010;
		Coeff[13743] <= 15'b111101111101011;
		Coeff[13744] <= 15'b111101111101100;
		Coeff[13745] <= 15'b111101111101101;
		Coeff[13746] <= 15'b111101111101110;
		Coeff[13747] <= 15'b111101111101110;
		Coeff[13748] <= 15'b111101111101111;
		Coeff[13749] <= 15'b111101111110000;
		Coeff[13750] <= 15'b111101111110001;
		Coeff[13751] <= 15'b111101111110001;
		Coeff[13752] <= 15'b111101111110010;
		Coeff[13753] <= 15'b111101111110011;
		Coeff[13754] <= 15'b111101111110100;
		Coeff[13755] <= 15'b111101111110101;
		Coeff[13756] <= 15'b111101111110101;
		Coeff[13757] <= 15'b111101111110110;
		Coeff[13758] <= 15'b111101111110111;
		Coeff[13759] <= 15'b111101111111000;
		Coeff[13760] <= 15'b111101111111001;
		Coeff[13761] <= 15'b111101111111001;
		Coeff[13762] <= 15'b111101111111010;
		Coeff[13763] <= 15'b111101111111011;
		Coeff[13764] <= 15'b111101111111100;
		Coeff[13765] <= 15'b111101111111100;
		Coeff[13766] <= 15'b111101111111101;
		Coeff[13767] <= 15'b111101111111110;
		Coeff[13768] <= 15'b111101111111111;
		Coeff[13769] <= 15'b111110000000000;
		Coeff[13770] <= 15'b111110000000000;
		Coeff[13771] <= 15'b111110000000001;
		Coeff[13772] <= 15'b111110000000010;
		Coeff[13773] <= 15'b111110000000011;
		Coeff[13774] <= 15'b111110000000011;
		Coeff[13775] <= 15'b111110000000100;
		Coeff[13776] <= 15'b111110000000101;
		Coeff[13777] <= 15'b111110000000110;
		Coeff[13778] <= 15'b111110000000111;
		Coeff[13779] <= 15'b111110000000111;
		Coeff[13780] <= 15'b111110000001000;
		Coeff[13781] <= 15'b111110000001001;
		Coeff[13782] <= 15'b111110000001010;
		Coeff[13783] <= 15'b111110000001010;
		Coeff[13784] <= 15'b111110000001011;
		Coeff[13785] <= 15'b111110000001100;
		Coeff[13786] <= 15'b111110000001101;
		Coeff[13787] <= 15'b111110000001110;
		Coeff[13788] <= 15'b111110000001110;
		Coeff[13789] <= 15'b111110000001111;
		Coeff[13790] <= 15'b111110000010000;
		Coeff[13791] <= 15'b111110000010001;
		Coeff[13792] <= 15'b111110000010001;
		Coeff[13793] <= 15'b111110000010010;
		Coeff[13794] <= 15'b111110000010011;
		Coeff[13795] <= 15'b111110000010100;
		Coeff[13796] <= 15'b111110000010100;
		Coeff[13797] <= 15'b111110000010101;
		Coeff[13798] <= 15'b111110000010110;
		Coeff[13799] <= 15'b111110000010111;
		Coeff[13800] <= 15'b111110000011000;
		Coeff[13801] <= 15'b111110000011000;
		Coeff[13802] <= 15'b111110000011001;
		Coeff[13803] <= 15'b111110000011010;
		Coeff[13804] <= 15'b111110000011011;
		Coeff[13805] <= 15'b111110000011011;
		Coeff[13806] <= 15'b111110000011100;
		Coeff[13807] <= 15'b111110000011101;
		Coeff[13808] <= 15'b111110000011110;
		Coeff[13809] <= 15'b111110000011111;
		Coeff[13810] <= 15'b111110000011111;
		Coeff[13811] <= 15'b111110000100000;
		Coeff[13812] <= 15'b111110000100001;
		Coeff[13813] <= 15'b111110000100010;
		Coeff[13814] <= 15'b111110000100010;
		Coeff[13815] <= 15'b111110000100011;
		Coeff[13816] <= 15'b111110000100100;
		Coeff[13817] <= 15'b111110000100101;
		Coeff[13818] <= 15'b111110000100101;
		Coeff[13819] <= 15'b111110000100110;
		Coeff[13820] <= 15'b111110000100111;
		Coeff[13821] <= 15'b111110000101000;
		Coeff[13822] <= 15'b111110000101000;
		Coeff[13823] <= 15'b111110000101001;
		Coeff[13824] <= 15'b111110000101010;
		Coeff[13825] <= 15'b111110000101011;
		Coeff[13826] <= 15'b111110000101100;
		Coeff[13827] <= 15'b111110000101100;
		Coeff[13828] <= 15'b111110000101101;
		Coeff[13829] <= 15'b111110000101110;
		Coeff[13830] <= 15'b111110000101111;
		Coeff[13831] <= 15'b111110000101111;
		Coeff[13832] <= 15'b111110000110000;
		Coeff[13833] <= 15'b111110000110001;
		Coeff[13834] <= 15'b111110000110010;
		Coeff[13835] <= 15'b111110000110010;
		Coeff[13836] <= 15'b111110000110011;
		Coeff[13837] <= 15'b111110000110100;
		Coeff[13838] <= 15'b111110000110101;
		Coeff[13839] <= 15'b111110000110101;
		Coeff[13840] <= 15'b111110000110110;
		Coeff[13841] <= 15'b111110000110111;
		Coeff[13842] <= 15'b111110000111000;
		Coeff[13843] <= 15'b111110000111000;
		Coeff[13844] <= 15'b111110000111001;
		Coeff[13845] <= 15'b111110000111010;
		Coeff[13846] <= 15'b111110000111011;
		Coeff[13847] <= 15'b111110000111011;
		Coeff[13848] <= 15'b111110000111100;
		Coeff[13849] <= 15'b111110000111101;
		Coeff[13850] <= 15'b111110000111110;
		Coeff[13851] <= 15'b111110000111110;
		Coeff[13852] <= 15'b111110000111111;
		Coeff[13853] <= 15'b111110001000000;
		Coeff[13854] <= 15'b111110001000001;
		Coeff[13855] <= 15'b111110001000010;
		Coeff[13856] <= 15'b111110001000010;
		Coeff[13857] <= 15'b111110001000011;
		Coeff[13858] <= 15'b111110001000100;
		Coeff[13859] <= 15'b111110001000101;
		Coeff[13860] <= 15'b111110001000101;
		Coeff[13861] <= 15'b111110001000110;
		Coeff[13862] <= 15'b111110001000111;
		Coeff[13863] <= 15'b111110001001000;
		Coeff[13864] <= 15'b111110001001000;
		Coeff[13865] <= 15'b111110001001001;
		Coeff[13866] <= 15'b111110001001010;
		Coeff[13867] <= 15'b111110001001011;
		Coeff[13868] <= 15'b111110001001011;
		Coeff[13869] <= 15'b111110001001100;
		Coeff[13870] <= 15'b111110001001101;
		Coeff[13871] <= 15'b111110001001110;
		Coeff[13872] <= 15'b111110001001110;
		Coeff[13873] <= 15'b111110001001111;
		Coeff[13874] <= 15'b111110001010000;
		Coeff[13875] <= 15'b111110001010001;
		Coeff[13876] <= 15'b111110001010001;
		Coeff[13877] <= 15'b111110001010010;
		Coeff[13878] <= 15'b111110001010011;
		Coeff[13879] <= 15'b111110001010100;
		Coeff[13880] <= 15'b111110001010100;
		Coeff[13881] <= 15'b111110001010101;
		Coeff[13882] <= 15'b111110001010110;
		Coeff[13883] <= 15'b111110001010111;
		Coeff[13884] <= 15'b111110001010111;
		Coeff[13885] <= 15'b111110001011000;
		Coeff[13886] <= 15'b111110001011001;
		Coeff[13887] <= 15'b111110001011001;
		Coeff[13888] <= 15'b111110001011010;
		Coeff[13889] <= 15'b111110001011011;
		Coeff[13890] <= 15'b111110001011100;
		Coeff[13891] <= 15'b111110001011100;
		Coeff[13892] <= 15'b111110001011101;
		Coeff[13893] <= 15'b111110001011110;
		Coeff[13894] <= 15'b111110001011111;
		Coeff[13895] <= 15'b111110001011111;
		Coeff[13896] <= 15'b111110001100000;
		Coeff[13897] <= 15'b111110001100001;
		Coeff[13898] <= 15'b111110001100010;
		Coeff[13899] <= 15'b111110001100010;
		Coeff[13900] <= 15'b111110001100011;
		Coeff[13901] <= 15'b111110001100100;
		Coeff[13902] <= 15'b111110001100101;
		Coeff[13903] <= 15'b111110001100101;
		Coeff[13904] <= 15'b111110001100110;
		Coeff[13905] <= 15'b111110001100111;
		Coeff[13906] <= 15'b111110001101000;
		Coeff[13907] <= 15'b111110001101000;
		Coeff[13908] <= 15'b111110001101001;
		Coeff[13909] <= 15'b111110001101010;
		Coeff[13910] <= 15'b111110001101011;
		Coeff[13911] <= 15'b111110001101011;
		Coeff[13912] <= 15'b111110001101100;
		Coeff[13913] <= 15'b111110001101101;
		Coeff[13914] <= 15'b111110001101110;
		Coeff[13915] <= 15'b111110001101110;
		Coeff[13916] <= 15'b111110001101111;
		Coeff[13917] <= 15'b111110001110000;
		Coeff[13918] <= 15'b111110001110000;
		Coeff[13919] <= 15'b111110001110001;
		Coeff[13920] <= 15'b111110001110010;
		Coeff[13921] <= 15'b111110001110011;
		Coeff[13922] <= 15'b111110001110011;
		Coeff[13923] <= 15'b111110001110100;
		Coeff[13924] <= 15'b111110001110101;
		Coeff[13925] <= 15'b111110001110110;
		Coeff[13926] <= 15'b111110001110110;
		Coeff[13927] <= 15'b111110001110111;
		Coeff[13928] <= 15'b111110001111000;
		Coeff[13929] <= 15'b111110001111001;
		Coeff[13930] <= 15'b111110001111001;
		Coeff[13931] <= 15'b111110001111010;
		Coeff[13932] <= 15'b111110001111011;
		Coeff[13933] <= 15'b111110001111011;
		Coeff[13934] <= 15'b111110001111100;
		Coeff[13935] <= 15'b111110001111101;
		Coeff[13936] <= 15'b111110001111110;
		Coeff[13937] <= 15'b111110001111110;
		Coeff[13938] <= 15'b111110001111111;
		Coeff[13939] <= 15'b111110010000000;
		Coeff[13940] <= 15'b111110010000001;
		Coeff[13941] <= 15'b111110010000001;
		Coeff[13942] <= 15'b111110010000010;
		Coeff[13943] <= 15'b111110010000011;
		Coeff[13944] <= 15'b111110010000011;
		Coeff[13945] <= 15'b111110010000100;
		Coeff[13946] <= 15'b111110010000101;
		Coeff[13947] <= 15'b111110010000110;
		Coeff[13948] <= 15'b111110010000110;
		Coeff[13949] <= 15'b111110010000111;
		Coeff[13950] <= 15'b111110010001000;
		Coeff[13951] <= 15'b111110010001001;
		Coeff[13952] <= 15'b111110010001001;
		Coeff[13953] <= 15'b111110010001010;
		Coeff[13954] <= 15'b111110010001011;
		Coeff[13955] <= 15'b111110010001011;
		Coeff[13956] <= 15'b111110010001100;
		Coeff[13957] <= 15'b111110010001101;
		Coeff[13958] <= 15'b111110010001110;
		Coeff[13959] <= 15'b111110010001110;
		Coeff[13960] <= 15'b111110010001111;
		Coeff[13961] <= 15'b111110010010000;
		Coeff[13962] <= 15'b111110010010001;
		Coeff[13963] <= 15'b111110010010001;
		Coeff[13964] <= 15'b111110010010010;
		Coeff[13965] <= 15'b111110010010011;
		Coeff[13966] <= 15'b111110010010011;
		Coeff[13967] <= 15'b111110010010100;
		Coeff[13968] <= 15'b111110010010101;
		Coeff[13969] <= 15'b111110010010110;
		Coeff[13970] <= 15'b111110010010110;
		Coeff[13971] <= 15'b111110010010111;
		Coeff[13972] <= 15'b111110010011000;
		Coeff[13973] <= 15'b111110010011000;
		Coeff[13974] <= 15'b111110010011001;
		Coeff[13975] <= 15'b111110010011010;
		Coeff[13976] <= 15'b111110010011011;
		Coeff[13977] <= 15'b111110010011011;
		Coeff[13978] <= 15'b111110010011100;
		Coeff[13979] <= 15'b111110010011101;
		Coeff[13980] <= 15'b111110010011110;
		Coeff[13981] <= 15'b111110010011110;
		Coeff[13982] <= 15'b111110010011111;
		Coeff[13983] <= 15'b111110010100000;
		Coeff[13984] <= 15'b111110010100000;
		Coeff[13985] <= 15'b111110010100001;
		Coeff[13986] <= 15'b111110010100010;
		Coeff[13987] <= 15'b111110010100011;
		Coeff[13988] <= 15'b111110010100011;
		Coeff[13989] <= 15'b111110010100100;
		Coeff[13990] <= 15'b111110010100101;
		Coeff[13991] <= 15'b111110010100101;
		Coeff[13992] <= 15'b111110010100110;
		Coeff[13993] <= 15'b111110010100111;
		Coeff[13994] <= 15'b111110010101000;
		Coeff[13995] <= 15'b111110010101000;
		Coeff[13996] <= 15'b111110010101001;
		Coeff[13997] <= 15'b111110010101010;
		Coeff[13998] <= 15'b111110010101010;
		Coeff[13999] <= 15'b111110010101011;
		Coeff[14000] <= 15'b111110010101100;
		Coeff[14001] <= 15'b111110010101101;
		Coeff[14002] <= 15'b111110010101101;
		Coeff[14003] <= 15'b111110010101110;
		Coeff[14004] <= 15'b111110010101111;
		Coeff[14005] <= 15'b111110010101111;
		Coeff[14006] <= 15'b111110010110000;
		Coeff[14007] <= 15'b111110010110001;
		Coeff[14008] <= 15'b111110010110001;
		Coeff[14009] <= 15'b111110010110010;
		Coeff[14010] <= 15'b111110010110011;
		Coeff[14011] <= 15'b111110010110100;
		Coeff[14012] <= 15'b111110010110100;
		Coeff[14013] <= 15'b111110010110101;
		Coeff[14014] <= 15'b111110010110110;
		Coeff[14015] <= 15'b111110010110110;
		Coeff[14016] <= 15'b111110010110111;
		Coeff[14017] <= 15'b111110010111000;
		Coeff[14018] <= 15'b111110010111001;
		Coeff[14019] <= 15'b111110010111001;
		Coeff[14020] <= 15'b111110010111010;
		Coeff[14021] <= 15'b111110010111011;
		Coeff[14022] <= 15'b111110010111011;
		Coeff[14023] <= 15'b111110010111100;
		Coeff[14024] <= 15'b111110010111101;
		Coeff[14025] <= 15'b111110010111110;
		Coeff[14026] <= 15'b111110010111110;
		Coeff[14027] <= 15'b111110010111111;
		Coeff[14028] <= 15'b111110011000000;
		Coeff[14029] <= 15'b111110011000000;
		Coeff[14030] <= 15'b111110011000001;
		Coeff[14031] <= 15'b111110011000010;
		Coeff[14032] <= 15'b111110011000010;
		Coeff[14033] <= 15'b111110011000011;
		Coeff[14034] <= 15'b111110011000100;
		Coeff[14035] <= 15'b111110011000101;
		Coeff[14036] <= 15'b111110011000101;
		Coeff[14037] <= 15'b111110011000110;
		Coeff[14038] <= 15'b111110011000111;
		Coeff[14039] <= 15'b111110011000111;
		Coeff[14040] <= 15'b111110011001000;
		Coeff[14041] <= 15'b111110011001001;
		Coeff[14042] <= 15'b111110011001001;
		Coeff[14043] <= 15'b111110011001010;
		Coeff[14044] <= 15'b111110011001011;
		Coeff[14045] <= 15'b111110011001100;
		Coeff[14046] <= 15'b111110011001100;
		Coeff[14047] <= 15'b111110011001101;
		Coeff[14048] <= 15'b111110011001110;
		Coeff[14049] <= 15'b111110011001110;
		Coeff[14050] <= 15'b111110011001111;
		Coeff[14051] <= 15'b111110011010000;
		Coeff[14052] <= 15'b111110011010000;
		Coeff[14053] <= 15'b111110011010001;
		Coeff[14054] <= 15'b111110011010010;
		Coeff[14055] <= 15'b111110011010011;
		Coeff[14056] <= 15'b111110011010011;
		Coeff[14057] <= 15'b111110011010100;
		Coeff[14058] <= 15'b111110011010101;
		Coeff[14059] <= 15'b111110011010101;
		Coeff[14060] <= 15'b111110011010110;
		Coeff[14061] <= 15'b111110011010111;
		Coeff[14062] <= 15'b111110011010111;
		Coeff[14063] <= 15'b111110011011000;
		Coeff[14064] <= 15'b111110011011001;
		Coeff[14065] <= 15'b111110011011001;
		Coeff[14066] <= 15'b111110011011010;
		Coeff[14067] <= 15'b111110011011011;
		Coeff[14068] <= 15'b111110011011100;
		Coeff[14069] <= 15'b111110011011100;
		Coeff[14070] <= 15'b111110011011101;
		Coeff[14071] <= 15'b111110011011110;
		Coeff[14072] <= 15'b111110011011110;
		Coeff[14073] <= 15'b111110011011111;
		Coeff[14074] <= 15'b111110011100000;
		Coeff[14075] <= 15'b111110011100000;
		Coeff[14076] <= 15'b111110011100001;
		Coeff[14077] <= 15'b111110011100010;
		Coeff[14078] <= 15'b111110011100010;
		Coeff[14079] <= 15'b111110011100011;
		Coeff[14080] <= 15'b111110011100100;
		Coeff[14081] <= 15'b111110011100100;
		Coeff[14082] <= 15'b111110011100101;
		Coeff[14083] <= 15'b111110011100110;
		Coeff[14084] <= 15'b111110011100111;
		Coeff[14085] <= 15'b111110011100111;
		Coeff[14086] <= 15'b111110011101000;
		Coeff[14087] <= 15'b111110011101001;
		Coeff[14088] <= 15'b111110011101001;
		Coeff[14089] <= 15'b111110011101010;
		Coeff[14090] <= 15'b111110011101011;
		Coeff[14091] <= 15'b111110011101011;
		Coeff[14092] <= 15'b111110011101100;
		Coeff[14093] <= 15'b111110011101101;
		Coeff[14094] <= 15'b111110011101101;
		Coeff[14095] <= 15'b111110011101110;
		Coeff[14096] <= 15'b111110011101111;
		Coeff[14097] <= 15'b111110011101111;
		Coeff[14098] <= 15'b111110011110000;
		Coeff[14099] <= 15'b111110011110001;
		Coeff[14100] <= 15'b111110011110010;
		Coeff[14101] <= 15'b111110011110010;
		Coeff[14102] <= 15'b111110011110011;
		Coeff[14103] <= 15'b111110011110100;
		Coeff[14104] <= 15'b111110011110100;
		Coeff[14105] <= 15'b111110011110101;
		Coeff[14106] <= 15'b111110011110110;
		Coeff[14107] <= 15'b111110011110110;
		Coeff[14108] <= 15'b111110011110111;
		Coeff[14109] <= 15'b111110011111000;
		Coeff[14110] <= 15'b111110011111000;
		Coeff[14111] <= 15'b111110011111001;
		Coeff[14112] <= 15'b111110011111010;
		Coeff[14113] <= 15'b111110011111010;
		Coeff[14114] <= 15'b111110011111011;
		Coeff[14115] <= 15'b111110011111100;
		Coeff[14116] <= 15'b111110011111100;
		Coeff[14117] <= 15'b111110011111101;
		Coeff[14118] <= 15'b111110011111110;
		Coeff[14119] <= 15'b111110011111110;
		Coeff[14120] <= 15'b111110011111111;
		Coeff[14121] <= 15'b111110100000000;
		Coeff[14122] <= 15'b111110100000000;
		Coeff[14123] <= 15'b111110100000001;
		Coeff[14124] <= 15'b111110100000010;
		Coeff[14125] <= 15'b111110100000010;
		Coeff[14126] <= 15'b111110100000011;
		Coeff[14127] <= 15'b111110100000100;
		Coeff[14128] <= 15'b111110100000101;
		Coeff[14129] <= 15'b111110100000101;
		Coeff[14130] <= 15'b111110100000110;
		Coeff[14131] <= 15'b111110100000111;
		Coeff[14132] <= 15'b111110100000111;
		Coeff[14133] <= 15'b111110100001000;
		Coeff[14134] <= 15'b111110100001001;
		Coeff[14135] <= 15'b111110100001001;
		Coeff[14136] <= 15'b111110100001010;
		Coeff[14137] <= 15'b111110100001011;
		Coeff[14138] <= 15'b111110100001011;
		Coeff[14139] <= 15'b111110100001100;
		Coeff[14140] <= 15'b111110100001101;
		Coeff[14141] <= 15'b111110100001101;
		Coeff[14142] <= 15'b111110100001110;
		Coeff[14143] <= 15'b111110100001111;
		Coeff[14144] <= 15'b111110100001111;
		Coeff[14145] <= 15'b111110100010000;
		Coeff[14146] <= 15'b111110100010001;
		Coeff[14147] <= 15'b111110100010001;
		Coeff[14148] <= 15'b111110100010010;
		Coeff[14149] <= 15'b111110100010011;
		Coeff[14150] <= 15'b111110100010011;
		Coeff[14151] <= 15'b111110100010100;
		Coeff[14152] <= 15'b111110100010101;
		Coeff[14153] <= 15'b111110100010101;
		Coeff[14154] <= 15'b111110100010110;
		Coeff[14155] <= 15'b111110100010111;
		Coeff[14156] <= 15'b111110100010111;
		Coeff[14157] <= 15'b111110100011000;
		Coeff[14158] <= 15'b111110100011001;
		Coeff[14159] <= 15'b111110100011001;
		Coeff[14160] <= 15'b111110100011010;
		Coeff[14161] <= 15'b111110100011011;
		Coeff[14162] <= 15'b111110100011011;
		Coeff[14163] <= 15'b111110100011100;
		Coeff[14164] <= 15'b111110100011101;
		Coeff[14165] <= 15'b111110100011101;
		Coeff[14166] <= 15'b111110100011110;
		Coeff[14167] <= 15'b111110100011111;
		Coeff[14168] <= 15'b111110100011111;
		Coeff[14169] <= 15'b111110100100000;
		Coeff[14170] <= 15'b111110100100001;
		Coeff[14171] <= 15'b111110100100001;
		Coeff[14172] <= 15'b111110100100010;
		Coeff[14173] <= 15'b111110100100011;
		Coeff[14174] <= 15'b111110100100011;
		Coeff[14175] <= 15'b111110100100100;
		Coeff[14176] <= 15'b111110100100101;
		Coeff[14177] <= 15'b111110100100101;
		Coeff[14178] <= 15'b111110100100110;
		Coeff[14179] <= 15'b111110100100111;
		Coeff[14180] <= 15'b111110100100111;
		Coeff[14181] <= 15'b111110100101000;
		Coeff[14182] <= 15'b111110100101000;
		Coeff[14183] <= 15'b111110100101001;
		Coeff[14184] <= 15'b111110100101010;
		Coeff[14185] <= 15'b111110100101010;
		Coeff[14186] <= 15'b111110100101011;
		Coeff[14187] <= 15'b111110100101100;
		Coeff[14188] <= 15'b111110100101100;
		Coeff[14189] <= 15'b111110100101101;
		Coeff[14190] <= 15'b111110100101110;
		Coeff[14191] <= 15'b111110100101110;
		Coeff[14192] <= 15'b111110100101111;
		Coeff[14193] <= 15'b111110100110000;
		Coeff[14194] <= 15'b111110100110000;
		Coeff[14195] <= 15'b111110100110001;
		Coeff[14196] <= 15'b111110100110010;
		Coeff[14197] <= 15'b111110100110010;
		Coeff[14198] <= 15'b111110100110011;
		Coeff[14199] <= 15'b111110100110100;
		Coeff[14200] <= 15'b111110100110100;
		Coeff[14201] <= 15'b111110100110101;
		Coeff[14202] <= 15'b111110100110110;
		Coeff[14203] <= 15'b111110100110110;
		Coeff[14204] <= 15'b111110100110111;
		Coeff[14205] <= 15'b111110100111000;
		Coeff[14206] <= 15'b111110100111000;
		Coeff[14207] <= 15'b111110100111001;
		Coeff[14208] <= 15'b111110100111010;
		Coeff[14209] <= 15'b111110100111010;
		Coeff[14210] <= 15'b111110100111011;
		Coeff[14211] <= 15'b111110100111011;
		Coeff[14212] <= 15'b111110100111100;
		Coeff[14213] <= 15'b111110100111101;
		Coeff[14214] <= 15'b111110100111101;
		Coeff[14215] <= 15'b111110100111110;
		Coeff[14216] <= 15'b111110100111111;
		Coeff[14217] <= 15'b111110100111111;
		Coeff[14218] <= 15'b111110101000000;
		Coeff[14219] <= 15'b111110101000001;
		Coeff[14220] <= 15'b111110101000001;
		Coeff[14221] <= 15'b111110101000010;
		Coeff[14222] <= 15'b111110101000011;
		Coeff[14223] <= 15'b111110101000011;
		Coeff[14224] <= 15'b111110101000100;
		Coeff[14225] <= 15'b111110101000101;
		Coeff[14226] <= 15'b111110101000101;
		Coeff[14227] <= 15'b111110101000110;
		Coeff[14228] <= 15'b111110101000110;
		Coeff[14229] <= 15'b111110101000111;
		Coeff[14230] <= 15'b111110101001000;
		Coeff[14231] <= 15'b111110101001000;
		Coeff[14232] <= 15'b111110101001001;
		Coeff[14233] <= 15'b111110101001010;
		Coeff[14234] <= 15'b111110101001010;
		Coeff[14235] <= 15'b111110101001011;
		Coeff[14236] <= 15'b111110101001100;
		Coeff[14237] <= 15'b111110101001100;
		Coeff[14238] <= 15'b111110101001101;
		Coeff[14239] <= 15'b111110101001110;
		Coeff[14240] <= 15'b111110101001110;
		Coeff[14241] <= 15'b111110101001111;
		Coeff[14242] <= 15'b111110101001111;
		Coeff[14243] <= 15'b111110101010000;
		Coeff[14244] <= 15'b111110101010001;
		Coeff[14245] <= 15'b111110101010001;
		Coeff[14246] <= 15'b111110101010010;
		Coeff[14247] <= 15'b111110101010011;
		Coeff[14248] <= 15'b111110101010011;
		Coeff[14249] <= 15'b111110101010100;
		Coeff[14250] <= 15'b111110101010101;
		Coeff[14251] <= 15'b111110101010101;
		Coeff[14252] <= 15'b111110101010110;
		Coeff[14253] <= 15'b111110101010110;
		Coeff[14254] <= 15'b111110101010111;
		Coeff[14255] <= 15'b111110101011000;
		Coeff[14256] <= 15'b111110101011000;
		Coeff[14257] <= 15'b111110101011001;
		Coeff[14258] <= 15'b111110101011010;
		Coeff[14259] <= 15'b111110101011010;
		Coeff[14260] <= 15'b111110101011011;
		Coeff[14261] <= 15'b111110101011100;
		Coeff[14262] <= 15'b111110101011100;
		Coeff[14263] <= 15'b111110101011101;
		Coeff[14264] <= 15'b111110101011101;
		Coeff[14265] <= 15'b111110101011110;
		Coeff[14266] <= 15'b111110101011111;
		Coeff[14267] <= 15'b111110101011111;
		Coeff[14268] <= 15'b111110101100000;
		Coeff[14269] <= 15'b111110101100001;
		Coeff[14270] <= 15'b111110101100001;
		Coeff[14271] <= 15'b111110101100010;
		Coeff[14272] <= 15'b111110101100011;
		Coeff[14273] <= 15'b111110101100011;
		Coeff[14274] <= 15'b111110101100100;
		Coeff[14275] <= 15'b111110101100100;
		Coeff[14276] <= 15'b111110101100101;
		Coeff[14277] <= 15'b111110101100110;
		Coeff[14278] <= 15'b111110101100110;
		Coeff[14279] <= 15'b111110101100111;
		Coeff[14280] <= 15'b111110101101000;
		Coeff[14281] <= 15'b111110101101000;
		Coeff[14282] <= 15'b111110101101001;
		Coeff[14283] <= 15'b111110101101001;
		Coeff[14284] <= 15'b111110101101010;
		Coeff[14285] <= 15'b111110101101011;
		Coeff[14286] <= 15'b111110101101011;
		Coeff[14287] <= 15'b111110101101100;
		Coeff[14288] <= 15'b111110101101101;
		Coeff[14289] <= 15'b111110101101101;
		Coeff[14290] <= 15'b111110101101110;
		Coeff[14291] <= 15'b111110101101110;
		Coeff[14292] <= 15'b111110101101111;
		Coeff[14293] <= 15'b111110101110000;
		Coeff[14294] <= 15'b111110101110000;
		Coeff[14295] <= 15'b111110101110001;
		Coeff[14296] <= 15'b111110101110010;
		Coeff[14297] <= 15'b111110101110010;
		Coeff[14298] <= 15'b111110101110011;
		Coeff[14299] <= 15'b111110101110011;
		Coeff[14300] <= 15'b111110101110100;
		Coeff[14301] <= 15'b111110101110101;
		Coeff[14302] <= 15'b111110101110101;
		Coeff[14303] <= 15'b111110101110110;
		Coeff[14304] <= 15'b111110101110111;
		Coeff[14305] <= 15'b111110101110111;
		Coeff[14306] <= 15'b111110101111000;
		Coeff[14307] <= 15'b111110101111000;
		Coeff[14308] <= 15'b111110101111001;
		Coeff[14309] <= 15'b111110101111010;
		Coeff[14310] <= 15'b111110101111010;
		Coeff[14311] <= 15'b111110101111011;
		Coeff[14312] <= 15'b111110101111100;
		Coeff[14313] <= 15'b111110101111100;
		Coeff[14314] <= 15'b111110101111101;
		Coeff[14315] <= 15'b111110101111101;
		Coeff[14316] <= 15'b111110101111110;
		Coeff[14317] <= 15'b111110101111111;
		Coeff[14318] <= 15'b111110101111111;
		Coeff[14319] <= 15'b111110110000000;
		Coeff[14320] <= 15'b111110110000001;
		Coeff[14321] <= 15'b111110110000001;
		Coeff[14322] <= 15'b111110110000010;
		Coeff[14323] <= 15'b111110110000010;
		Coeff[14324] <= 15'b111110110000011;
		Coeff[14325] <= 15'b111110110000100;
		Coeff[14326] <= 15'b111110110000100;
		Coeff[14327] <= 15'b111110110000101;
		Coeff[14328] <= 15'b111110110000101;
		Coeff[14329] <= 15'b111110110000110;
		Coeff[14330] <= 15'b111110110000111;
		Coeff[14331] <= 15'b111110110000111;
		Coeff[14332] <= 15'b111110110001000;
		Coeff[14333] <= 15'b111110110001001;
		Coeff[14334] <= 15'b111110110001001;
		Coeff[14335] <= 15'b111110110001010;
		Coeff[14336] <= 15'b111110110001010;
		Coeff[14337] <= 15'b111110110001011;
		Coeff[14338] <= 15'b111110110001100;
		Coeff[14339] <= 15'b111110110001100;
		Coeff[14340] <= 15'b111110110001101;
		Coeff[14341] <= 15'b111110110001101;
		Coeff[14342] <= 15'b111110110001110;
		Coeff[14343] <= 15'b111110110001111;
		Coeff[14344] <= 15'b111110110001111;
		Coeff[14345] <= 15'b111110110010000;
		Coeff[14346] <= 15'b111110110010000;
		Coeff[14347] <= 15'b111110110010001;
		Coeff[14348] <= 15'b111110110010010;
		Coeff[14349] <= 15'b111110110010010;
		Coeff[14350] <= 15'b111110110010011;
		Coeff[14351] <= 15'b111110110010100;
		Coeff[14352] <= 15'b111110110010100;
		Coeff[14353] <= 15'b111110110010101;
		Coeff[14354] <= 15'b111110110010101;
		Coeff[14355] <= 15'b111110110010110;
		Coeff[14356] <= 15'b111110110010111;
		Coeff[14357] <= 15'b111110110010111;
		Coeff[14358] <= 15'b111110110011000;
		Coeff[14359] <= 15'b111110110011000;
		Coeff[14360] <= 15'b111110110011001;
		Coeff[14361] <= 15'b111110110011010;
		Coeff[14362] <= 15'b111110110011010;
		Coeff[14363] <= 15'b111110110011011;
		Coeff[14364] <= 15'b111110110011011;
		Coeff[14365] <= 15'b111110110011100;
		Coeff[14366] <= 15'b111110110011101;
		Coeff[14367] <= 15'b111110110011101;
		Coeff[14368] <= 15'b111110110011110;
		Coeff[14369] <= 15'b111110110011110;
		Coeff[14370] <= 15'b111110110011111;
		Coeff[14371] <= 15'b111110110100000;
		Coeff[14372] <= 15'b111110110100000;
		Coeff[14373] <= 15'b111110110100001;
		Coeff[14374] <= 15'b111110110100001;
		Coeff[14375] <= 15'b111110110100010;
		Coeff[14376] <= 15'b111110110100011;
		Coeff[14377] <= 15'b111110110100011;
		Coeff[14378] <= 15'b111110110100100;
		Coeff[14379] <= 15'b111110110100100;
		Coeff[14380] <= 15'b111110110100101;
		Coeff[14381] <= 15'b111110110100110;
		Coeff[14382] <= 15'b111110110100110;
		Coeff[14383] <= 15'b111110110100111;
		Coeff[14384] <= 15'b111110110100111;
		Coeff[14385] <= 15'b111110110101000;
		Coeff[14386] <= 15'b111110110101001;
		Coeff[14387] <= 15'b111110110101001;
		Coeff[14388] <= 15'b111110110101010;
		Coeff[14389] <= 15'b111110110101010;
		Coeff[14390] <= 15'b111110110101011;
		Coeff[14391] <= 15'b111110110101100;
		Coeff[14392] <= 15'b111110110101100;
		Coeff[14393] <= 15'b111110110101101;
		Coeff[14394] <= 15'b111110110101101;
		Coeff[14395] <= 15'b111110110101110;
		Coeff[14396] <= 15'b111110110101111;
		Coeff[14397] <= 15'b111110110101111;
		Coeff[14398] <= 15'b111110110110000;
		Coeff[14399] <= 15'b111110110110000;
		Coeff[14400] <= 15'b111110110110001;
		Coeff[14401] <= 15'b111110110110010;
		Coeff[14402] <= 15'b111110110110010;
		Coeff[14403] <= 15'b111110110110011;
		Coeff[14404] <= 15'b111110110110011;
		Coeff[14405] <= 15'b111110110110100;
		Coeff[14406] <= 15'b111110110110101;
		Coeff[14407] <= 15'b111110110110101;
		Coeff[14408] <= 15'b111110110110110;
		Coeff[14409] <= 15'b111110110110110;
		Coeff[14410] <= 15'b111110110110111;
		Coeff[14411] <= 15'b111110110111000;
		Coeff[14412] <= 15'b111110110111000;
		Coeff[14413] <= 15'b111110110111001;
		Coeff[14414] <= 15'b111110110111001;
		Coeff[14415] <= 15'b111110110111010;
		Coeff[14416] <= 15'b111110110111010;
		Coeff[14417] <= 15'b111110110111011;
		Coeff[14418] <= 15'b111110110111100;
		Coeff[14419] <= 15'b111110110111100;
		Coeff[14420] <= 15'b111110110111101;
		Coeff[14421] <= 15'b111110110111101;
		Coeff[14422] <= 15'b111110110111110;
		Coeff[14423] <= 15'b111110110111111;
		Coeff[14424] <= 15'b111110110111111;
		Coeff[14425] <= 15'b111110111000000;
		Coeff[14426] <= 15'b111110111000000;
		Coeff[14427] <= 15'b111110111000001;
		Coeff[14428] <= 15'b111110111000010;
		Coeff[14429] <= 15'b111110111000010;
		Coeff[14430] <= 15'b111110111000011;
		Coeff[14431] <= 15'b111110111000011;
		Coeff[14432] <= 15'b111110111000100;
		Coeff[14433] <= 15'b111110111000100;
		Coeff[14434] <= 15'b111110111000101;
		Coeff[14435] <= 15'b111110111000110;
		Coeff[14436] <= 15'b111110111000110;
		Coeff[14437] <= 15'b111110111000111;
		Coeff[14438] <= 15'b111110111000111;
		Coeff[14439] <= 15'b111110111001000;
		Coeff[14440] <= 15'b111110111001001;
		Coeff[14441] <= 15'b111110111001001;
		Coeff[14442] <= 15'b111110111001010;
		Coeff[14443] <= 15'b111110111001010;
		Coeff[14444] <= 15'b111110111001011;
		Coeff[14445] <= 15'b111110111001011;
		Coeff[14446] <= 15'b111110111001100;
		Coeff[14447] <= 15'b111110111001101;
		Coeff[14448] <= 15'b111110111001101;
		Coeff[14449] <= 15'b111110111001110;
		Coeff[14450] <= 15'b111110111001110;
		Coeff[14451] <= 15'b111110111001111;
		Coeff[14452] <= 15'b111110111001111;
		Coeff[14453] <= 15'b111110111010000;
		Coeff[14454] <= 15'b111110111010001;
		Coeff[14455] <= 15'b111110111010001;
		Coeff[14456] <= 15'b111110111010010;
		Coeff[14457] <= 15'b111110111010010;
		Coeff[14458] <= 15'b111110111010011;
		Coeff[14459] <= 15'b111110111010100;
		Coeff[14460] <= 15'b111110111010100;
		Coeff[14461] <= 15'b111110111010101;
		Coeff[14462] <= 15'b111110111010101;
		Coeff[14463] <= 15'b111110111010110;
		Coeff[14464] <= 15'b111110111010110;
		Coeff[14465] <= 15'b111110111010111;
		Coeff[14466] <= 15'b111110111011000;
		Coeff[14467] <= 15'b111110111011000;
		Coeff[14468] <= 15'b111110111011001;
		Coeff[14469] <= 15'b111110111011001;
		Coeff[14470] <= 15'b111110111011010;
		Coeff[14471] <= 15'b111110111011010;
		Coeff[14472] <= 15'b111110111011011;
		Coeff[14473] <= 15'b111110111011100;
		Coeff[14474] <= 15'b111110111011100;
		Coeff[14475] <= 15'b111110111011101;
		Coeff[14476] <= 15'b111110111011101;
		Coeff[14477] <= 15'b111110111011110;
		Coeff[14478] <= 15'b111110111011110;
		Coeff[14479] <= 15'b111110111011111;
		Coeff[14480] <= 15'b111110111100000;
		Coeff[14481] <= 15'b111110111100000;
		Coeff[14482] <= 15'b111110111100001;
		Coeff[14483] <= 15'b111110111100001;
		Coeff[14484] <= 15'b111110111100010;
		Coeff[14485] <= 15'b111110111100010;
		Coeff[14486] <= 15'b111110111100011;
		Coeff[14487] <= 15'b111110111100100;
		Coeff[14488] <= 15'b111110111100100;
		Coeff[14489] <= 15'b111110111100101;
		Coeff[14490] <= 15'b111110111100101;
		Coeff[14491] <= 15'b111110111100110;
		Coeff[14492] <= 15'b111110111100110;
		Coeff[14493] <= 15'b111110111100111;
		Coeff[14494] <= 15'b111110111101000;
		Coeff[14495] <= 15'b111110111101000;
		Coeff[14496] <= 15'b111110111101001;
		Coeff[14497] <= 15'b111110111101001;
		Coeff[14498] <= 15'b111110111101010;
		Coeff[14499] <= 15'b111110111101010;
		Coeff[14500] <= 15'b111110111101011;
		Coeff[14501] <= 15'b111110111101011;
		Coeff[14502] <= 15'b111110111101100;
		Coeff[14503] <= 15'b111110111101101;
		Coeff[14504] <= 15'b111110111101101;
		Coeff[14505] <= 15'b111110111101110;
		Coeff[14506] <= 15'b111110111101110;
		Coeff[14507] <= 15'b111110111101111;
		Coeff[14508] <= 15'b111110111101111;
		Coeff[14509] <= 15'b111110111110000;
		Coeff[14510] <= 15'b111110111110001;
		Coeff[14511] <= 15'b111110111110001;
		Coeff[14512] <= 15'b111110111110010;
		Coeff[14513] <= 15'b111110111110010;
		Coeff[14514] <= 15'b111110111110011;
		Coeff[14515] <= 15'b111110111110011;
		Coeff[14516] <= 15'b111110111110100;
		Coeff[14517] <= 15'b111110111110100;
		Coeff[14518] <= 15'b111110111110101;
		Coeff[14519] <= 15'b111110111110110;
		Coeff[14520] <= 15'b111110111110110;
		Coeff[14521] <= 15'b111110111110111;
		Coeff[14522] <= 15'b111110111110111;
		Coeff[14523] <= 15'b111110111111000;
		Coeff[14524] <= 15'b111110111111000;
		Coeff[14525] <= 15'b111110111111001;
		Coeff[14526] <= 15'b111110111111001;
		Coeff[14527] <= 15'b111110111111010;
		Coeff[14528] <= 15'b111110111111011;
		Coeff[14529] <= 15'b111110111111011;
		Coeff[14530] <= 15'b111110111111100;
		Coeff[14531] <= 15'b111110111111100;
		Coeff[14532] <= 15'b111110111111101;
		Coeff[14533] <= 15'b111110111111101;
		Coeff[14534] <= 15'b111110111111110;
		Coeff[14535] <= 15'b111110111111110;
		Coeff[14536] <= 15'b111110111111111;
		Coeff[14537] <= 15'b111111000000000;
		Coeff[14538] <= 15'b111111000000000;
		Coeff[14539] <= 15'b111111000000001;
		Coeff[14540] <= 15'b111111000000001;
		Coeff[14541] <= 15'b111111000000010;
		Coeff[14542] <= 15'b111111000000010;
		Coeff[14543] <= 15'b111111000000011;
		Coeff[14544] <= 15'b111111000000011;
		Coeff[14545] <= 15'b111111000000100;
		Coeff[14546] <= 15'b111111000000101;
		Coeff[14547] <= 15'b111111000000101;
		Coeff[14548] <= 15'b111111000000110;
		Coeff[14549] <= 15'b111111000000110;
		Coeff[14550] <= 15'b111111000000111;
		Coeff[14551] <= 15'b111111000000111;
		Coeff[14552] <= 15'b111111000001000;
		Coeff[14553] <= 15'b111111000001000;
		Coeff[14554] <= 15'b111111000001001;
		Coeff[14555] <= 15'b111111000001010;
		Coeff[14556] <= 15'b111111000001010;
		Coeff[14557] <= 15'b111111000001011;
		Coeff[14558] <= 15'b111111000001011;
		Coeff[14559] <= 15'b111111000001100;
		Coeff[14560] <= 15'b111111000001100;
		Coeff[14561] <= 15'b111111000001101;
		Coeff[14562] <= 15'b111111000001101;
		Coeff[14563] <= 15'b111111000001110;
		Coeff[14564] <= 15'b111111000001110;
		Coeff[14565] <= 15'b111111000001111;
		Coeff[14566] <= 15'b111111000010000;
		Coeff[14567] <= 15'b111111000010000;
		Coeff[14568] <= 15'b111111000010001;
		Coeff[14569] <= 15'b111111000010001;
		Coeff[14570] <= 15'b111111000010010;
		Coeff[14571] <= 15'b111111000010010;
		Coeff[14572] <= 15'b111111000010011;
		Coeff[14573] <= 15'b111111000010011;
		Coeff[14574] <= 15'b111111000010100;
		Coeff[14575] <= 15'b111111000010100;
		Coeff[14576] <= 15'b111111000010101;
		Coeff[14577] <= 15'b111111000010101;
		Coeff[14578] <= 15'b111111000010110;
		Coeff[14579] <= 15'b111111000010111;
		Coeff[14580] <= 15'b111111000010111;
		Coeff[14581] <= 15'b111111000011000;
		Coeff[14582] <= 15'b111111000011000;
		Coeff[14583] <= 15'b111111000011001;
		Coeff[14584] <= 15'b111111000011001;
		Coeff[14585] <= 15'b111111000011010;
		Coeff[14586] <= 15'b111111000011010;
		Coeff[14587] <= 15'b111111000011011;
		Coeff[14588] <= 15'b111111000011011;
		Coeff[14589] <= 15'b111111000011100;
		Coeff[14590] <= 15'b111111000011101;
		Coeff[14591] <= 15'b111111000011101;
		Coeff[14592] <= 15'b111111000011110;
		Coeff[14593] <= 15'b111111000011110;
		Coeff[14594] <= 15'b111111000011111;
		Coeff[14595] <= 15'b111111000011111;
		Coeff[14596] <= 15'b111111000100000;
		Coeff[14597] <= 15'b111111000100000;
		Coeff[14598] <= 15'b111111000100001;
		Coeff[14599] <= 15'b111111000100001;
		Coeff[14600] <= 15'b111111000100010;
		Coeff[14601] <= 15'b111111000100010;
		Coeff[14602] <= 15'b111111000100011;
		Coeff[14603] <= 15'b111111000100011;
		Coeff[14604] <= 15'b111111000100100;
		Coeff[14605] <= 15'b111111000100101;
		Coeff[14606] <= 15'b111111000100101;
		Coeff[14607] <= 15'b111111000100110;
		Coeff[14608] <= 15'b111111000100110;
		Coeff[14609] <= 15'b111111000100111;
		Coeff[14610] <= 15'b111111000100111;
		Coeff[14611] <= 15'b111111000101000;
		Coeff[14612] <= 15'b111111000101000;
		Coeff[14613] <= 15'b111111000101001;
		Coeff[14614] <= 15'b111111000101001;
		Coeff[14615] <= 15'b111111000101010;
		Coeff[14616] <= 15'b111111000101010;
		Coeff[14617] <= 15'b111111000101011;
		Coeff[14618] <= 15'b111111000101011;
		Coeff[14619] <= 15'b111111000101100;
		Coeff[14620] <= 15'b111111000101101;
		Coeff[14621] <= 15'b111111000101101;
		Coeff[14622] <= 15'b111111000101110;
		Coeff[14623] <= 15'b111111000101110;
		Coeff[14624] <= 15'b111111000101111;
		Coeff[14625] <= 15'b111111000101111;
		Coeff[14626] <= 15'b111111000110000;
		Coeff[14627] <= 15'b111111000110000;
		Coeff[14628] <= 15'b111111000110001;
		Coeff[14629] <= 15'b111111000110001;
		Coeff[14630] <= 15'b111111000110010;
		Coeff[14631] <= 15'b111111000110010;
		Coeff[14632] <= 15'b111111000110011;
		Coeff[14633] <= 15'b111111000110011;
		Coeff[14634] <= 15'b111111000110100;
		Coeff[14635] <= 15'b111111000110100;
		Coeff[14636] <= 15'b111111000110101;
		Coeff[14637] <= 15'b111111000110101;
		Coeff[14638] <= 15'b111111000110110;
		Coeff[14639] <= 15'b111111000110110;
		Coeff[14640] <= 15'b111111000110111;
		Coeff[14641] <= 15'b111111000111000;
		Coeff[14642] <= 15'b111111000111000;
		Coeff[14643] <= 15'b111111000111001;
		Coeff[14644] <= 15'b111111000111001;
		Coeff[14645] <= 15'b111111000111010;
		Coeff[14646] <= 15'b111111000111010;
		Coeff[14647] <= 15'b111111000111011;
		Coeff[14648] <= 15'b111111000111011;
		Coeff[14649] <= 15'b111111000111100;
		Coeff[14650] <= 15'b111111000111100;
		Coeff[14651] <= 15'b111111000111101;
		Coeff[14652] <= 15'b111111000111101;
		Coeff[14653] <= 15'b111111000111110;
		Coeff[14654] <= 15'b111111000111110;
		Coeff[14655] <= 15'b111111000111111;
		Coeff[14656] <= 15'b111111000111111;
		Coeff[14657] <= 15'b111111001000000;
		Coeff[14658] <= 15'b111111001000000;
		Coeff[14659] <= 15'b111111001000001;
		Coeff[14660] <= 15'b111111001000001;
		Coeff[14661] <= 15'b111111001000010;
		Coeff[14662] <= 15'b111111001000010;
		Coeff[14663] <= 15'b111111001000011;
		Coeff[14664] <= 15'b111111001000011;
		Coeff[14665] <= 15'b111111001000100;
		Coeff[14666] <= 15'b111111001000101;
		Coeff[14667] <= 15'b111111001000101;
		Coeff[14668] <= 15'b111111001000110;
		Coeff[14669] <= 15'b111111001000110;
		Coeff[14670] <= 15'b111111001000111;
		Coeff[14671] <= 15'b111111001000111;
		Coeff[14672] <= 15'b111111001001000;
		Coeff[14673] <= 15'b111111001001000;
		Coeff[14674] <= 15'b111111001001001;
		Coeff[14675] <= 15'b111111001001001;
		Coeff[14676] <= 15'b111111001001010;
		Coeff[14677] <= 15'b111111001001010;
		Coeff[14678] <= 15'b111111001001011;
		Coeff[14679] <= 15'b111111001001011;
		Coeff[14680] <= 15'b111111001001100;
		Coeff[14681] <= 15'b111111001001100;
		Coeff[14682] <= 15'b111111001001101;
		Coeff[14683] <= 15'b111111001001101;
		Coeff[14684] <= 15'b111111001001110;
		Coeff[14685] <= 15'b111111001001110;
		Coeff[14686] <= 15'b111111001001111;
		Coeff[14687] <= 15'b111111001001111;
		Coeff[14688] <= 15'b111111001010000;
		Coeff[14689] <= 15'b111111001010000;
		Coeff[14690] <= 15'b111111001010001;
		Coeff[14691] <= 15'b111111001010001;
		Coeff[14692] <= 15'b111111001010010;
		Coeff[14693] <= 15'b111111001010010;
		Coeff[14694] <= 15'b111111001010011;
		Coeff[14695] <= 15'b111111001010011;
		Coeff[14696] <= 15'b111111001010100;
		Coeff[14697] <= 15'b111111001010100;
		Coeff[14698] <= 15'b111111001010101;
		Coeff[14699] <= 15'b111111001010101;
		Coeff[14700] <= 15'b111111001010110;
		Coeff[14701] <= 15'b111111001010110;
		Coeff[14702] <= 15'b111111001010111;
		Coeff[14703] <= 15'b111111001010111;
		Coeff[14704] <= 15'b111111001011000;
		Coeff[14705] <= 15'b111111001011000;
		Coeff[14706] <= 15'b111111001011001;
		Coeff[14707] <= 15'b111111001011001;
		Coeff[14708] <= 15'b111111001011010;
		Coeff[14709] <= 15'b111111001011010;
		Coeff[14710] <= 15'b111111001011011;
		Coeff[14711] <= 15'b111111001011011;
		Coeff[14712] <= 15'b111111001011100;
		Coeff[14713] <= 15'b111111001011100;
		Coeff[14714] <= 15'b111111001011101;
		Coeff[14715] <= 15'b111111001011101;
		Coeff[14716] <= 15'b111111001011110;
		Coeff[14717] <= 15'b111111001011110;
		Coeff[14718] <= 15'b111111001011111;
		Coeff[14719] <= 15'b111111001011111;
		Coeff[14720] <= 15'b111111001100000;
		Coeff[14721] <= 15'b111111001100000;
		Coeff[14722] <= 15'b111111001100001;
		Coeff[14723] <= 15'b111111001100001;
		Coeff[14724] <= 15'b111111001100010;
		Coeff[14725] <= 15'b111111001100010;
		Coeff[14726] <= 15'b111111001100011;
		Coeff[14727] <= 15'b111111001100011;
		Coeff[14728] <= 15'b111111001100100;
		Coeff[14729] <= 15'b111111001100100;
		Coeff[14730] <= 15'b111111001100101;
		Coeff[14731] <= 15'b111111001100101;
		Coeff[14732] <= 15'b111111001100110;
		Coeff[14733] <= 15'b111111001100110;
		Coeff[14734] <= 15'b111111001100111;
		Coeff[14735] <= 15'b111111001100111;
		Coeff[14736] <= 15'b111111001101000;
		Coeff[14737] <= 15'b111111001101000;
		Coeff[14738] <= 15'b111111001101001;
		Coeff[14739] <= 15'b111111001101001;
		Coeff[14740] <= 15'b111111001101010;
		Coeff[14741] <= 15'b111111001101010;
		Coeff[14742] <= 15'b111111001101011;
		Coeff[14743] <= 15'b111111001101011;
		Coeff[14744] <= 15'b111111001101100;
		Coeff[14745] <= 15'b111111001101100;
		Coeff[14746] <= 15'b111111001101101;
		Coeff[14747] <= 15'b111111001101101;
		Coeff[14748] <= 15'b111111001101110;
		Coeff[14749] <= 15'b111111001101110;
		Coeff[14750] <= 15'b111111001101111;
		Coeff[14751] <= 15'b111111001101111;
		Coeff[14752] <= 15'b111111001110000;
		Coeff[14753] <= 15'b111111001110000;
		Coeff[14754] <= 15'b111111001110001;
		Coeff[14755] <= 15'b111111001110001;
		Coeff[14756] <= 15'b111111001110010;
		Coeff[14757] <= 15'b111111001110010;
		Coeff[14758] <= 15'b111111001110011;
		Coeff[14759] <= 15'b111111001110011;
		Coeff[14760] <= 15'b111111001110100;
		Coeff[14761] <= 15'b111111001110100;
		Coeff[14762] <= 15'b111111001110101;
		Coeff[14763] <= 15'b111111001110101;
		Coeff[14764] <= 15'b111111001110110;
		Coeff[14765] <= 15'b111111001110110;
		Coeff[14766] <= 15'b111111001110111;
		Coeff[14767] <= 15'b111111001110111;
		Coeff[14768] <= 15'b111111001111000;
		Coeff[14769] <= 15'b111111001111000;
		Coeff[14770] <= 15'b111111001111000;
		Coeff[14771] <= 15'b111111001111001;
		Coeff[14772] <= 15'b111111001111001;
		Coeff[14773] <= 15'b111111001111010;
		Coeff[14774] <= 15'b111111001111010;
		Coeff[14775] <= 15'b111111001111011;
		Coeff[14776] <= 15'b111111001111011;
		Coeff[14777] <= 15'b111111001111100;
		Coeff[14778] <= 15'b111111001111100;
		Coeff[14779] <= 15'b111111001111101;
		Coeff[14780] <= 15'b111111001111101;
		Coeff[14781] <= 15'b111111001111110;
		Coeff[14782] <= 15'b111111001111110;
		Coeff[14783] <= 15'b111111001111111;
		Coeff[14784] <= 15'b111111001111111;
		Coeff[14785] <= 15'b111111010000000;
		Coeff[14786] <= 15'b111111010000000;
		Coeff[14787] <= 15'b111111010000001;
		Coeff[14788] <= 15'b111111010000001;
		Coeff[14789] <= 15'b111111010000010;
		Coeff[14790] <= 15'b111111010000010;
		Coeff[14791] <= 15'b111111010000011;
		Coeff[14792] <= 15'b111111010000011;
		Coeff[14793] <= 15'b111111010000100;
		Coeff[14794] <= 15'b111111010000100;
		Coeff[14795] <= 15'b111111010000100;
		Coeff[14796] <= 15'b111111010000101;
		Coeff[14797] <= 15'b111111010000101;
		Coeff[14798] <= 15'b111111010000110;
		Coeff[14799] <= 15'b111111010000110;
		Coeff[14800] <= 15'b111111010000111;
		Coeff[14801] <= 15'b111111010000111;
		Coeff[14802] <= 15'b111111010001000;
		Coeff[14803] <= 15'b111111010001000;
		Coeff[14804] <= 15'b111111010001001;
		Coeff[14805] <= 15'b111111010001001;
		Coeff[14806] <= 15'b111111010001010;
		Coeff[14807] <= 15'b111111010001010;
		Coeff[14808] <= 15'b111111010001011;
		Coeff[14809] <= 15'b111111010001011;
		Coeff[14810] <= 15'b111111010001100;
		Coeff[14811] <= 15'b111111010001100;
		Coeff[14812] <= 15'b111111010001101;
		Coeff[14813] <= 15'b111111010001101;
		Coeff[14814] <= 15'b111111010001101;
		Coeff[14815] <= 15'b111111010001110;
		Coeff[14816] <= 15'b111111010001110;
		Coeff[14817] <= 15'b111111010001111;
		Coeff[14818] <= 15'b111111010001111;
		Coeff[14819] <= 15'b111111010010000;
		Coeff[14820] <= 15'b111111010010000;
		Coeff[14821] <= 15'b111111010010001;
		Coeff[14822] <= 15'b111111010010001;
		Coeff[14823] <= 15'b111111010010010;
		Coeff[14824] <= 15'b111111010010010;
		Coeff[14825] <= 15'b111111010010011;
		Coeff[14826] <= 15'b111111010010011;
		Coeff[14827] <= 15'b111111010010100;
		Coeff[14828] <= 15'b111111010010100;
		Coeff[14829] <= 15'b111111010010101;
		Coeff[14830] <= 15'b111111010010101;
		Coeff[14831] <= 15'b111111010010101;
		Coeff[14832] <= 15'b111111010010110;
		Coeff[14833] <= 15'b111111010010110;
		Coeff[14834] <= 15'b111111010010111;
		Coeff[14835] <= 15'b111111010010111;
		Coeff[14836] <= 15'b111111010011000;
		Coeff[14837] <= 15'b111111010011000;
		Coeff[14838] <= 15'b111111010011001;
		Coeff[14839] <= 15'b111111010011001;
		Coeff[14840] <= 15'b111111010011010;
		Coeff[14841] <= 15'b111111010011010;
		Coeff[14842] <= 15'b111111010011011;
		Coeff[14843] <= 15'b111111010011011;
		Coeff[14844] <= 15'b111111010011011;
		Coeff[14845] <= 15'b111111010011100;
		Coeff[14846] <= 15'b111111010011100;
		Coeff[14847] <= 15'b111111010011101;
		Coeff[14848] <= 15'b111111010011101;
		Coeff[14849] <= 15'b111111010011110;
		Coeff[14850] <= 15'b111111010011110;
		Coeff[14851] <= 15'b111111010011111;
		Coeff[14852] <= 15'b111111010011111;
		Coeff[14853] <= 15'b111111010100000;
		Coeff[14854] <= 15'b111111010100000;
		Coeff[14855] <= 15'b111111010100001;
		Coeff[14856] <= 15'b111111010100001;
		Coeff[14857] <= 15'b111111010100001;
		Coeff[14858] <= 15'b111111010100010;
		Coeff[14859] <= 15'b111111010100010;
		Coeff[14860] <= 15'b111111010100011;
		Coeff[14861] <= 15'b111111010100011;
		Coeff[14862] <= 15'b111111010100100;
		Coeff[14863] <= 15'b111111010100100;
		Coeff[14864] <= 15'b111111010100101;
		Coeff[14865] <= 15'b111111010100101;
		Coeff[14866] <= 15'b111111010100110;
		Coeff[14867] <= 15'b111111010100110;
		Coeff[14868] <= 15'b111111010100110;
		Coeff[14869] <= 15'b111111010100111;
		Coeff[14870] <= 15'b111111010100111;
		Coeff[14871] <= 15'b111111010101000;
		Coeff[14872] <= 15'b111111010101000;
		Coeff[14873] <= 15'b111111010101001;
		Coeff[14874] <= 15'b111111010101001;
		Coeff[14875] <= 15'b111111010101010;
		Coeff[14876] <= 15'b111111010101010;
		Coeff[14877] <= 15'b111111010101011;
		Coeff[14878] <= 15'b111111010101011;
		Coeff[14879] <= 15'b111111010101011;
		Coeff[14880] <= 15'b111111010101100;
		Coeff[14881] <= 15'b111111010101100;
		Coeff[14882] <= 15'b111111010101101;
		Coeff[14883] <= 15'b111111010101101;
		Coeff[14884] <= 15'b111111010101110;
		Coeff[14885] <= 15'b111111010101110;
		Coeff[14886] <= 15'b111111010101111;
		Coeff[14887] <= 15'b111111010101111;
		Coeff[14888] <= 15'b111111010110000;
		Coeff[14889] <= 15'b111111010110000;
		Coeff[14890] <= 15'b111111010110000;
		Coeff[14891] <= 15'b111111010110001;
		Coeff[14892] <= 15'b111111010110001;
		Coeff[14893] <= 15'b111111010110010;
		Coeff[14894] <= 15'b111111010110010;
		Coeff[14895] <= 15'b111111010110011;
		Coeff[14896] <= 15'b111111010110011;
		Coeff[14897] <= 15'b111111010110100;
		Coeff[14898] <= 15'b111111010110100;
		Coeff[14899] <= 15'b111111010110100;
		Coeff[14900] <= 15'b111111010110101;
		Coeff[14901] <= 15'b111111010110101;
		Coeff[14902] <= 15'b111111010110110;
		Coeff[14903] <= 15'b111111010110110;
		Coeff[14904] <= 15'b111111010110111;
		Coeff[14905] <= 15'b111111010110111;
		Coeff[14906] <= 15'b111111010111000;
		Coeff[14907] <= 15'b111111010111000;
		Coeff[14908] <= 15'b111111010111000;
		Coeff[14909] <= 15'b111111010111001;
		Coeff[14910] <= 15'b111111010111001;
		Coeff[14911] <= 15'b111111010111010;
		Coeff[14912] <= 15'b111111010111010;
		Coeff[14913] <= 15'b111111010111011;
		Coeff[14914] <= 15'b111111010111011;
		Coeff[14915] <= 15'b111111010111100;
		Coeff[14916] <= 15'b111111010111100;
		Coeff[14917] <= 15'b111111010111100;
		Coeff[14918] <= 15'b111111010111101;
		Coeff[14919] <= 15'b111111010111101;
		Coeff[14920] <= 15'b111111010111110;
		Coeff[14921] <= 15'b111111010111110;
		Coeff[14922] <= 15'b111111010111111;
		Coeff[14923] <= 15'b111111010111111;
		Coeff[14924] <= 15'b111111011000000;
		Coeff[14925] <= 15'b111111011000000;
		Coeff[14926] <= 15'b111111011000000;
		Coeff[14927] <= 15'b111111011000001;
		Coeff[14928] <= 15'b111111011000001;
		Coeff[14929] <= 15'b111111011000010;
		Coeff[14930] <= 15'b111111011000010;
		Coeff[14931] <= 15'b111111011000011;
		Coeff[14932] <= 15'b111111011000011;
		Coeff[14933] <= 15'b111111011000011;
		Coeff[14934] <= 15'b111111011000100;
		Coeff[14935] <= 15'b111111011000100;
		Coeff[14936] <= 15'b111111011000101;
		Coeff[14937] <= 15'b111111011000101;
		Coeff[14938] <= 15'b111111011000110;
		Coeff[14939] <= 15'b111111011000110;
		Coeff[14940] <= 15'b111111011000110;
		Coeff[14941] <= 15'b111111011000111;
		Coeff[14942] <= 15'b111111011000111;
		Coeff[14943] <= 15'b111111011001000;
		Coeff[14944] <= 15'b111111011001000;
		Coeff[14945] <= 15'b111111011001001;
		Coeff[14946] <= 15'b111111011001001;
		Coeff[14947] <= 15'b111111011001010;
		Coeff[14948] <= 15'b111111011001010;
		Coeff[14949] <= 15'b111111011001010;
		Coeff[14950] <= 15'b111111011001011;
		Coeff[14951] <= 15'b111111011001011;
		Coeff[14952] <= 15'b111111011001100;
		Coeff[14953] <= 15'b111111011001100;
		Coeff[14954] <= 15'b111111011001101;
		Coeff[14955] <= 15'b111111011001101;
		Coeff[14956] <= 15'b111111011001101;
		Coeff[14957] <= 15'b111111011001110;
		Coeff[14958] <= 15'b111111011001110;
		Coeff[14959] <= 15'b111111011001111;
		Coeff[14960] <= 15'b111111011001111;
		Coeff[14961] <= 15'b111111011010000;
		Coeff[14962] <= 15'b111111011010000;
		Coeff[14963] <= 15'b111111011010000;
		Coeff[14964] <= 15'b111111011010001;
		Coeff[14965] <= 15'b111111011010001;
		Coeff[14966] <= 15'b111111011010010;
		Coeff[14967] <= 15'b111111011010010;
		Coeff[14968] <= 15'b111111011010011;
		Coeff[14969] <= 15'b111111011010011;
		Coeff[14970] <= 15'b111111011010011;
		Coeff[14971] <= 15'b111111011010100;
		Coeff[14972] <= 15'b111111011010100;
		Coeff[14973] <= 15'b111111011010101;
		Coeff[14974] <= 15'b111111011010101;
		Coeff[14975] <= 15'b111111011010101;
		Coeff[14976] <= 15'b111111011010110;
		Coeff[14977] <= 15'b111111011010110;
		Coeff[14978] <= 15'b111111011010111;
		Coeff[14979] <= 15'b111111011010111;
		Coeff[14980] <= 15'b111111011011000;
		Coeff[14981] <= 15'b111111011011000;
		Coeff[14982] <= 15'b111111011011000;
		Coeff[14983] <= 15'b111111011011001;
		Coeff[14984] <= 15'b111111011011001;
		Coeff[14985] <= 15'b111111011011010;
		Coeff[14986] <= 15'b111111011011010;
		Coeff[14987] <= 15'b111111011011011;
		Coeff[14988] <= 15'b111111011011011;
		Coeff[14989] <= 15'b111111011011011;
		Coeff[14990] <= 15'b111111011011100;
		Coeff[14991] <= 15'b111111011011100;
		Coeff[14992] <= 15'b111111011011101;
		Coeff[14993] <= 15'b111111011011101;
		Coeff[14994] <= 15'b111111011011101;
		Coeff[14995] <= 15'b111111011011110;
		Coeff[14996] <= 15'b111111011011110;
		Coeff[14997] <= 15'b111111011011111;
		Coeff[14998] <= 15'b111111011011111;
		Coeff[14999] <= 15'b111111011100000;
		Coeff[15000] <= 15'b111111011100000;
		Coeff[15001] <= 15'b111111011100000;
		Coeff[15002] <= 15'b111111011100001;
		Coeff[15003] <= 15'b111111011100001;
		Coeff[15004] <= 15'b111111011100010;
		Coeff[15005] <= 15'b111111011100010;
		Coeff[15006] <= 15'b111111011100010;
		Coeff[15007] <= 15'b111111011100011;
		Coeff[15008] <= 15'b111111011100011;
		Coeff[15009] <= 15'b111111011100100;
		Coeff[15010] <= 15'b111111011100100;
		Coeff[15011] <= 15'b111111011100101;
		Coeff[15012] <= 15'b111111011100101;
		Coeff[15013] <= 15'b111111011100101;
		Coeff[15014] <= 15'b111111011100110;
		Coeff[15015] <= 15'b111111011100110;
		Coeff[15016] <= 15'b111111011100111;
		Coeff[15017] <= 15'b111111011100111;
		Coeff[15018] <= 15'b111111011100111;
		Coeff[15019] <= 15'b111111011101000;
		Coeff[15020] <= 15'b111111011101000;
		Coeff[15021] <= 15'b111111011101001;
		Coeff[15022] <= 15'b111111011101001;
		Coeff[15023] <= 15'b111111011101001;
		Coeff[15024] <= 15'b111111011101010;
		Coeff[15025] <= 15'b111111011101010;
		Coeff[15026] <= 15'b111111011101011;
		Coeff[15027] <= 15'b111111011101011;
		Coeff[15028] <= 15'b111111011101011;
		Coeff[15029] <= 15'b111111011101100;
		Coeff[15030] <= 15'b111111011101100;
		Coeff[15031] <= 15'b111111011101101;
		Coeff[15032] <= 15'b111111011101101;
		Coeff[15033] <= 15'b111111011101110;
		Coeff[15034] <= 15'b111111011101110;
		Coeff[15035] <= 15'b111111011101110;
		Coeff[15036] <= 15'b111111011101111;
		Coeff[15037] <= 15'b111111011101111;
		Coeff[15038] <= 15'b111111011110000;
		Coeff[15039] <= 15'b111111011110000;
		Coeff[15040] <= 15'b111111011110000;
		Coeff[15041] <= 15'b111111011110001;
		Coeff[15042] <= 15'b111111011110001;
		Coeff[15043] <= 15'b111111011110010;
		Coeff[15044] <= 15'b111111011110010;
		Coeff[15045] <= 15'b111111011110010;
		Coeff[15046] <= 15'b111111011110011;
		Coeff[15047] <= 15'b111111011110011;
		Coeff[15048] <= 15'b111111011110100;
		Coeff[15049] <= 15'b111111011110100;
		Coeff[15050] <= 15'b111111011110100;
		Coeff[15051] <= 15'b111111011110101;
		Coeff[15052] <= 15'b111111011110101;
		Coeff[15053] <= 15'b111111011110110;
		Coeff[15054] <= 15'b111111011110110;
		Coeff[15055] <= 15'b111111011110110;
		Coeff[15056] <= 15'b111111011110111;
		Coeff[15057] <= 15'b111111011110111;
		Coeff[15058] <= 15'b111111011111000;
		Coeff[15059] <= 15'b111111011111000;
		Coeff[15060] <= 15'b111111011111000;
		Coeff[15061] <= 15'b111111011111001;
		Coeff[15062] <= 15'b111111011111001;
		Coeff[15063] <= 15'b111111011111010;
		Coeff[15064] <= 15'b111111011111010;
		Coeff[15065] <= 15'b111111011111010;
		Coeff[15066] <= 15'b111111011111011;
		Coeff[15067] <= 15'b111111011111011;
		Coeff[15068] <= 15'b111111011111100;
		Coeff[15069] <= 15'b111111011111100;
		Coeff[15070] <= 15'b111111011111100;
		Coeff[15071] <= 15'b111111011111101;
		Coeff[15072] <= 15'b111111011111101;
		Coeff[15073] <= 15'b111111011111110;
		Coeff[15074] <= 15'b111111011111110;
		Coeff[15075] <= 15'b111111011111110;
		Coeff[15076] <= 15'b111111011111111;
		Coeff[15077] <= 15'b111111011111111;
		Coeff[15078] <= 15'b111111011111111;
		Coeff[15079] <= 15'b111111100000000;
		Coeff[15080] <= 15'b111111100000000;
		Coeff[15081] <= 15'b111111100000001;
		Coeff[15082] <= 15'b111111100000001;
		Coeff[15083] <= 15'b111111100000001;
		Coeff[15084] <= 15'b111111100000010;
		Coeff[15085] <= 15'b111111100000010;
		Coeff[15086] <= 15'b111111100000011;
		Coeff[15087] <= 15'b111111100000011;
		Coeff[15088] <= 15'b111111100000011;
		Coeff[15089] <= 15'b111111100000100;
		Coeff[15090] <= 15'b111111100000100;
		Coeff[15091] <= 15'b111111100000101;
		Coeff[15092] <= 15'b111111100000101;
		Coeff[15093] <= 15'b111111100000101;
		Coeff[15094] <= 15'b111111100000110;
		Coeff[15095] <= 15'b111111100000110;
		Coeff[15096] <= 15'b111111100000110;
		Coeff[15097] <= 15'b111111100000111;
		Coeff[15098] <= 15'b111111100000111;
		Coeff[15099] <= 15'b111111100001000;
		Coeff[15100] <= 15'b111111100001000;
		Coeff[15101] <= 15'b111111100001000;
		Coeff[15102] <= 15'b111111100001001;
		Coeff[15103] <= 15'b111111100001001;
		Coeff[15104] <= 15'b111111100001010;
		Coeff[15105] <= 15'b111111100001010;
		Coeff[15106] <= 15'b111111100001010;
		Coeff[15107] <= 15'b111111100001011;
		Coeff[15108] <= 15'b111111100001011;
		Coeff[15109] <= 15'b111111100001011;
		Coeff[15110] <= 15'b111111100001100;
		Coeff[15111] <= 15'b111111100001100;
		Coeff[15112] <= 15'b111111100001101;
		Coeff[15113] <= 15'b111111100001101;
		Coeff[15114] <= 15'b111111100001101;
		Coeff[15115] <= 15'b111111100001110;
		Coeff[15116] <= 15'b111111100001110;
		Coeff[15117] <= 15'b111111100001111;
		Coeff[15118] <= 15'b111111100001111;
		Coeff[15119] <= 15'b111111100001111;
		Coeff[15120] <= 15'b111111100010000;
		Coeff[15121] <= 15'b111111100010000;
		Coeff[15122] <= 15'b111111100010000;
		Coeff[15123] <= 15'b111111100010001;
		Coeff[15124] <= 15'b111111100010001;
		Coeff[15125] <= 15'b111111100010010;
		Coeff[15126] <= 15'b111111100010010;
		Coeff[15127] <= 15'b111111100010010;
		Coeff[15128] <= 15'b111111100010011;
		Coeff[15129] <= 15'b111111100010011;
		Coeff[15130] <= 15'b111111100010011;
		Coeff[15131] <= 15'b111111100010100;
		Coeff[15132] <= 15'b111111100010100;
		Coeff[15133] <= 15'b111111100010101;
		Coeff[15134] <= 15'b111111100010101;
		Coeff[15135] <= 15'b111111100010101;
		Coeff[15136] <= 15'b111111100010110;
		Coeff[15137] <= 15'b111111100010110;
		Coeff[15138] <= 15'b111111100010110;
		Coeff[15139] <= 15'b111111100010111;
		Coeff[15140] <= 15'b111111100010111;
		Coeff[15141] <= 15'b111111100011000;
		Coeff[15142] <= 15'b111111100011000;
		Coeff[15143] <= 15'b111111100011000;
		Coeff[15144] <= 15'b111111100011001;
		Coeff[15145] <= 15'b111111100011001;
		Coeff[15146] <= 15'b111111100011001;
		Coeff[15147] <= 15'b111111100011010;
		Coeff[15148] <= 15'b111111100011010;
		Coeff[15149] <= 15'b111111100011011;
		Coeff[15150] <= 15'b111111100011011;
		Coeff[15151] <= 15'b111111100011011;
		Coeff[15152] <= 15'b111111100011100;
		Coeff[15153] <= 15'b111111100011100;
		Coeff[15154] <= 15'b111111100011100;
		Coeff[15155] <= 15'b111111100011101;
		Coeff[15156] <= 15'b111111100011101;
		Coeff[15157] <= 15'b111111100011110;
		Coeff[15158] <= 15'b111111100011110;
		Coeff[15159] <= 15'b111111100011110;
		Coeff[15160] <= 15'b111111100011111;
		Coeff[15161] <= 15'b111111100011111;
		Coeff[15162] <= 15'b111111100011111;
		Coeff[15163] <= 15'b111111100100000;
		Coeff[15164] <= 15'b111111100100000;
		Coeff[15165] <= 15'b111111100100000;
		Coeff[15166] <= 15'b111111100100001;
		Coeff[15167] <= 15'b111111100100001;
		Coeff[15168] <= 15'b111111100100010;
		Coeff[15169] <= 15'b111111100100010;
		Coeff[15170] <= 15'b111111100100010;
		Coeff[15171] <= 15'b111111100100011;
		Coeff[15172] <= 15'b111111100100011;
		Coeff[15173] <= 15'b111111100100011;
		Coeff[15174] <= 15'b111111100100100;
		Coeff[15175] <= 15'b111111100100100;
		Coeff[15176] <= 15'b111111100100100;
		Coeff[15177] <= 15'b111111100100101;
		Coeff[15178] <= 15'b111111100100101;
		Coeff[15179] <= 15'b111111100100110;
		Coeff[15180] <= 15'b111111100100110;
		Coeff[15181] <= 15'b111111100100110;
		Coeff[15182] <= 15'b111111100100111;
		Coeff[15183] <= 15'b111111100100111;
		Coeff[15184] <= 15'b111111100100111;
		Coeff[15185] <= 15'b111111100101000;
		Coeff[15186] <= 15'b111111100101000;
		Coeff[15187] <= 15'b111111100101000;
		Coeff[15188] <= 15'b111111100101001;
		Coeff[15189] <= 15'b111111100101001;
		Coeff[15190] <= 15'b111111100101010;
		Coeff[15191] <= 15'b111111100101010;
		Coeff[15192] <= 15'b111111100101010;
		Coeff[15193] <= 15'b111111100101011;
		Coeff[15194] <= 15'b111111100101011;
		Coeff[15195] <= 15'b111111100101011;
		Coeff[15196] <= 15'b111111100101100;
		Coeff[15197] <= 15'b111111100101100;
		Coeff[15198] <= 15'b111111100101100;
		Coeff[15199] <= 15'b111111100101101;
		Coeff[15200] <= 15'b111111100101101;
		Coeff[15201] <= 15'b111111100101101;
		Coeff[15202] <= 15'b111111100101110;
		Coeff[15203] <= 15'b111111100101110;
		Coeff[15204] <= 15'b111111100101111;
		Coeff[15205] <= 15'b111111100101111;
		Coeff[15206] <= 15'b111111100101111;
		Coeff[15207] <= 15'b111111100110000;
		Coeff[15208] <= 15'b111111100110000;
		Coeff[15209] <= 15'b111111100110000;
		Coeff[15210] <= 15'b111111100110001;
		Coeff[15211] <= 15'b111111100110001;
		Coeff[15212] <= 15'b111111100110001;
		Coeff[15213] <= 15'b111111100110010;
		Coeff[15214] <= 15'b111111100110010;
		Coeff[15215] <= 15'b111111100110010;
		Coeff[15216] <= 15'b111111100110011;
		Coeff[15217] <= 15'b111111100110011;
		Coeff[15218] <= 15'b111111100110011;
		Coeff[15219] <= 15'b111111100110100;
		Coeff[15220] <= 15'b111111100110100;
		Coeff[15221] <= 15'b111111100110101;
		Coeff[15222] <= 15'b111111100110101;
		Coeff[15223] <= 15'b111111100110101;
		Coeff[15224] <= 15'b111111100110110;
		Coeff[15225] <= 15'b111111100110110;
		Coeff[15226] <= 15'b111111100110110;
		Coeff[15227] <= 15'b111111100110111;
		Coeff[15228] <= 15'b111111100110111;
		Coeff[15229] <= 15'b111111100110111;
		Coeff[15230] <= 15'b111111100111000;
		Coeff[15231] <= 15'b111111100111000;
		Coeff[15232] <= 15'b111111100111000;
		Coeff[15233] <= 15'b111111100111001;
		Coeff[15234] <= 15'b111111100111001;
		Coeff[15235] <= 15'b111111100111001;
		Coeff[15236] <= 15'b111111100111010;
		Coeff[15237] <= 15'b111111100111010;
		Coeff[15238] <= 15'b111111100111010;
		Coeff[15239] <= 15'b111111100111011;
		Coeff[15240] <= 15'b111111100111011;
		Coeff[15241] <= 15'b111111100111011;
		Coeff[15242] <= 15'b111111100111100;
		Coeff[15243] <= 15'b111111100111100;
		Coeff[15244] <= 15'b111111100111100;
		Coeff[15245] <= 15'b111111100111101;
		Coeff[15246] <= 15'b111111100111101;
		Coeff[15247] <= 15'b111111100111110;
		Coeff[15248] <= 15'b111111100111110;
		Coeff[15249] <= 15'b111111100111110;
		Coeff[15250] <= 15'b111111100111111;
		Coeff[15251] <= 15'b111111100111111;
		Coeff[15252] <= 15'b111111100111111;
		Coeff[15253] <= 15'b111111101000000;
		Coeff[15254] <= 15'b111111101000000;
		Coeff[15255] <= 15'b111111101000000;
		Coeff[15256] <= 15'b111111101000001;
		Coeff[15257] <= 15'b111111101000001;
		Coeff[15258] <= 15'b111111101000001;
		Coeff[15259] <= 15'b111111101000010;
		Coeff[15260] <= 15'b111111101000010;
		Coeff[15261] <= 15'b111111101000010;
		Coeff[15262] <= 15'b111111101000011;
		Coeff[15263] <= 15'b111111101000011;
		Coeff[15264] <= 15'b111111101000011;
		Coeff[15265] <= 15'b111111101000100;
		Coeff[15266] <= 15'b111111101000100;
		Coeff[15267] <= 15'b111111101000100;
		Coeff[15268] <= 15'b111111101000101;
		Coeff[15269] <= 15'b111111101000101;
		Coeff[15270] <= 15'b111111101000101;
		Coeff[15271] <= 15'b111111101000110;
		Coeff[15272] <= 15'b111111101000110;
		Coeff[15273] <= 15'b111111101000110;
		Coeff[15274] <= 15'b111111101000111;
		Coeff[15275] <= 15'b111111101000111;
		Coeff[15276] <= 15'b111111101000111;
		Coeff[15277] <= 15'b111111101001000;
		Coeff[15278] <= 15'b111111101001000;
		Coeff[15279] <= 15'b111111101001000;
		Coeff[15280] <= 15'b111111101001001;
		Coeff[15281] <= 15'b111111101001001;
		Coeff[15282] <= 15'b111111101001001;
		Coeff[15283] <= 15'b111111101001010;
		Coeff[15284] <= 15'b111111101001010;
		Coeff[15285] <= 15'b111111101001010;
		Coeff[15286] <= 15'b111111101001011;
		Coeff[15287] <= 15'b111111101001011;
		Coeff[15288] <= 15'b111111101001011;
		Coeff[15289] <= 15'b111111101001100;
		Coeff[15290] <= 15'b111111101001100;
		Coeff[15291] <= 15'b111111101001100;
		Coeff[15292] <= 15'b111111101001101;
		Coeff[15293] <= 15'b111111101001101;
		Coeff[15294] <= 15'b111111101001101;
		Coeff[15295] <= 15'b111111101001110;
		Coeff[15296] <= 15'b111111101001110;
		Coeff[15297] <= 15'b111111101001110;
		Coeff[15298] <= 15'b111111101001111;
		Coeff[15299] <= 15'b111111101001111;
		Coeff[15300] <= 15'b111111101001111;
		Coeff[15301] <= 15'b111111101010000;
		Coeff[15302] <= 15'b111111101010000;
		Coeff[15303] <= 15'b111111101010000;
		Coeff[15304] <= 15'b111111101010000;
		Coeff[15305] <= 15'b111111101010001;
		Coeff[15306] <= 15'b111111101010001;
		Coeff[15307] <= 15'b111111101010001;
		Coeff[15308] <= 15'b111111101010010;
		Coeff[15309] <= 15'b111111101010010;
		Coeff[15310] <= 15'b111111101010010;
		Coeff[15311] <= 15'b111111101010011;
		Coeff[15312] <= 15'b111111101010011;
		Coeff[15313] <= 15'b111111101010011;
		Coeff[15314] <= 15'b111111101010100;
		Coeff[15315] <= 15'b111111101010100;
		Coeff[15316] <= 15'b111111101010100;
		Coeff[15317] <= 15'b111111101010101;
		Coeff[15318] <= 15'b111111101010101;
		Coeff[15319] <= 15'b111111101010101;
		Coeff[15320] <= 15'b111111101010110;
		Coeff[15321] <= 15'b111111101010110;
		Coeff[15322] <= 15'b111111101010110;
		Coeff[15323] <= 15'b111111101010111;
		Coeff[15324] <= 15'b111111101010111;
		Coeff[15325] <= 15'b111111101010111;
		Coeff[15326] <= 15'b111111101011000;
		Coeff[15327] <= 15'b111111101011000;
		Coeff[15328] <= 15'b111111101011000;
		Coeff[15329] <= 15'b111111101011001;
		Coeff[15330] <= 15'b111111101011001;
		Coeff[15331] <= 15'b111111101011001;
		Coeff[15332] <= 15'b111111101011001;
		Coeff[15333] <= 15'b111111101011010;
		Coeff[15334] <= 15'b111111101011010;
		Coeff[15335] <= 15'b111111101011010;
		Coeff[15336] <= 15'b111111101011011;
		Coeff[15337] <= 15'b111111101011011;
		Coeff[15338] <= 15'b111111101011011;
		Coeff[15339] <= 15'b111111101011100;
		Coeff[15340] <= 15'b111111101011100;
		Coeff[15341] <= 15'b111111101011100;
		Coeff[15342] <= 15'b111111101011101;
		Coeff[15343] <= 15'b111111101011101;
		Coeff[15344] <= 15'b111111101011101;
		Coeff[15345] <= 15'b111111101011110;
		Coeff[15346] <= 15'b111111101011110;
		Coeff[15347] <= 15'b111111101011110;
		Coeff[15348] <= 15'b111111101011110;
		Coeff[15349] <= 15'b111111101011111;
		Coeff[15350] <= 15'b111111101011111;
		Coeff[15351] <= 15'b111111101011111;
		Coeff[15352] <= 15'b111111101100000;
		Coeff[15353] <= 15'b111111101100000;
		Coeff[15354] <= 15'b111111101100000;
		Coeff[15355] <= 15'b111111101100001;
		Coeff[15356] <= 15'b111111101100001;
		Coeff[15357] <= 15'b111111101100001;
		Coeff[15358] <= 15'b111111101100010;
		Coeff[15359] <= 15'b111111101100010;
		Coeff[15360] <= 15'b111111101100010;
		Coeff[15361] <= 15'b111111101100011;
		Coeff[15362] <= 15'b111111101100011;
		Coeff[15363] <= 15'b111111101100011;
		Coeff[15364] <= 15'b111111101100011;
		Coeff[15365] <= 15'b111111101100100;
		Coeff[15366] <= 15'b111111101100100;
		Coeff[15367] <= 15'b111111101100100;
		Coeff[15368] <= 15'b111111101100101;
		Coeff[15369] <= 15'b111111101100101;
		Coeff[15370] <= 15'b111111101100101;
		Coeff[15371] <= 15'b111111101100110;
		Coeff[15372] <= 15'b111111101100110;
		Coeff[15373] <= 15'b111111101100110;
		Coeff[15374] <= 15'b111111101100110;
		Coeff[15375] <= 15'b111111101100111;
		Coeff[15376] <= 15'b111111101100111;
		Coeff[15377] <= 15'b111111101100111;
		Coeff[15378] <= 15'b111111101101000;
		Coeff[15379] <= 15'b111111101101000;
		Coeff[15380] <= 15'b111111101101000;
		Coeff[15381] <= 15'b111111101101001;
		Coeff[15382] <= 15'b111111101101001;
		Coeff[15383] <= 15'b111111101101001;
		Coeff[15384] <= 15'b111111101101010;
		Coeff[15385] <= 15'b111111101101010;
		Coeff[15386] <= 15'b111111101101010;
		Coeff[15387] <= 15'b111111101101010;
		Coeff[15388] <= 15'b111111101101011;
		Coeff[15389] <= 15'b111111101101011;
		Coeff[15390] <= 15'b111111101101011;
		Coeff[15391] <= 15'b111111101101100;
		Coeff[15392] <= 15'b111111101101100;
		Coeff[15393] <= 15'b111111101101100;
		Coeff[15394] <= 15'b111111101101101;
		Coeff[15395] <= 15'b111111101101101;
		Coeff[15396] <= 15'b111111101101101;
		Coeff[15397] <= 15'b111111101101101;
		Coeff[15398] <= 15'b111111101101110;
		Coeff[15399] <= 15'b111111101101110;
		Coeff[15400] <= 15'b111111101101110;
		Coeff[15401] <= 15'b111111101101111;
		Coeff[15402] <= 15'b111111101101111;
		Coeff[15403] <= 15'b111111101101111;
		Coeff[15404] <= 15'b111111101101111;
		Coeff[15405] <= 15'b111111101110000;
		Coeff[15406] <= 15'b111111101110000;
		Coeff[15407] <= 15'b111111101110000;
		Coeff[15408] <= 15'b111111101110001;
		Coeff[15409] <= 15'b111111101110001;
		Coeff[15410] <= 15'b111111101110001;
		Coeff[15411] <= 15'b111111101110010;
		Coeff[15412] <= 15'b111111101110010;
		Coeff[15413] <= 15'b111111101110010;
		Coeff[15414] <= 15'b111111101110010;
		Coeff[15415] <= 15'b111111101110011;
		Coeff[15416] <= 15'b111111101110011;
		Coeff[15417] <= 15'b111111101110011;
		Coeff[15418] <= 15'b111111101110100;
		Coeff[15419] <= 15'b111111101110100;
		Coeff[15420] <= 15'b111111101110100;
		Coeff[15421] <= 15'b111111101110100;
		Coeff[15422] <= 15'b111111101110101;
		Coeff[15423] <= 15'b111111101110101;
		Coeff[15424] <= 15'b111111101110101;
		Coeff[15425] <= 15'b111111101110110;
		Coeff[15426] <= 15'b111111101110110;
		Coeff[15427] <= 15'b111111101110110;
		Coeff[15428] <= 15'b111111101110110;
		Coeff[15429] <= 15'b111111101110111;
		Coeff[15430] <= 15'b111111101110111;
		Coeff[15431] <= 15'b111111101110111;
		Coeff[15432] <= 15'b111111101111000;
		Coeff[15433] <= 15'b111111101111000;
		Coeff[15434] <= 15'b111111101111000;
		Coeff[15435] <= 15'b111111101111000;
		Coeff[15436] <= 15'b111111101111001;
		Coeff[15437] <= 15'b111111101111001;
		Coeff[15438] <= 15'b111111101111001;
		Coeff[15439] <= 15'b111111101111010;
		Coeff[15440] <= 15'b111111101111010;
		Coeff[15441] <= 15'b111111101111010;
		Coeff[15442] <= 15'b111111101111010;
		Coeff[15443] <= 15'b111111101111011;
		Coeff[15444] <= 15'b111111101111011;
		Coeff[15445] <= 15'b111111101111011;
		Coeff[15446] <= 15'b111111101111100;
		Coeff[15447] <= 15'b111111101111100;
		Coeff[15448] <= 15'b111111101111100;
		Coeff[15449] <= 15'b111111101111100;
		Coeff[15450] <= 15'b111111101111101;
		Coeff[15451] <= 15'b111111101111101;
		Coeff[15452] <= 15'b111111101111101;
		Coeff[15453] <= 15'b111111101111110;
		Coeff[15454] <= 15'b111111101111110;
		Coeff[15455] <= 15'b111111101111110;
		Coeff[15456] <= 15'b111111101111110;
		Coeff[15457] <= 15'b111111101111111;
		Coeff[15458] <= 15'b111111101111111;
		Coeff[15459] <= 15'b111111101111111;
		Coeff[15460] <= 15'b111111110000000;
		Coeff[15461] <= 15'b111111110000000;
		Coeff[15462] <= 15'b111111110000000;
		Coeff[15463] <= 15'b111111110000000;
		Coeff[15464] <= 15'b111111110000001;
		Coeff[15465] <= 15'b111111110000001;
		Coeff[15466] <= 15'b111111110000001;
		Coeff[15467] <= 15'b111111110000001;
		Coeff[15468] <= 15'b111111110000010;
		Coeff[15469] <= 15'b111111110000010;
		Coeff[15470] <= 15'b111111110000010;
		Coeff[15471] <= 15'b111111110000011;
		Coeff[15472] <= 15'b111111110000011;
		Coeff[15473] <= 15'b111111110000011;
		Coeff[15474] <= 15'b111111110000011;
		Coeff[15475] <= 15'b111111110000100;
		Coeff[15476] <= 15'b111111110000100;
		Coeff[15477] <= 15'b111111110000100;
		Coeff[15478] <= 15'b111111110000100;
		Coeff[15479] <= 15'b111111110000101;
		Coeff[15480] <= 15'b111111110000101;
		Coeff[15481] <= 15'b111111110000101;
		Coeff[15482] <= 15'b111111110000110;
		Coeff[15483] <= 15'b111111110000110;
		Coeff[15484] <= 15'b111111110000110;
		Coeff[15485] <= 15'b111111110000110;
		Coeff[15486] <= 15'b111111110000111;
		Coeff[15487] <= 15'b111111110000111;
		Coeff[15488] <= 15'b111111110000111;
		Coeff[15489] <= 15'b111111110000111;
		Coeff[15490] <= 15'b111111110001000;
		Coeff[15491] <= 15'b111111110001000;
		Coeff[15492] <= 15'b111111110001000;
		Coeff[15493] <= 15'b111111110001001;
		Coeff[15494] <= 15'b111111110001001;
		Coeff[15495] <= 15'b111111110001001;
		Coeff[15496] <= 15'b111111110001001;
		Coeff[15497] <= 15'b111111110001010;
		Coeff[15498] <= 15'b111111110001010;
		Coeff[15499] <= 15'b111111110001010;
		Coeff[15500] <= 15'b111111110001010;
		Coeff[15501] <= 15'b111111110001011;
		Coeff[15502] <= 15'b111111110001011;
		Coeff[15503] <= 15'b111111110001011;
		Coeff[15504] <= 15'b111111110001011;
		Coeff[15505] <= 15'b111111110001100;
		Coeff[15506] <= 15'b111111110001100;
		Coeff[15507] <= 15'b111111110001100;
		Coeff[15508] <= 15'b111111110001101;
		Coeff[15509] <= 15'b111111110001101;
		Coeff[15510] <= 15'b111111110001101;
		Coeff[15511] <= 15'b111111110001101;
		Coeff[15512] <= 15'b111111110001110;
		Coeff[15513] <= 15'b111111110001110;
		Coeff[15514] <= 15'b111111110001110;
		Coeff[15515] <= 15'b111111110001110;
		Coeff[15516] <= 15'b111111110001111;
		Coeff[15517] <= 15'b111111110001111;
		Coeff[15518] <= 15'b111111110001111;
		Coeff[15519] <= 15'b111111110001111;
		Coeff[15520] <= 15'b111111110010000;
		Coeff[15521] <= 15'b111111110010000;
		Coeff[15522] <= 15'b111111110010000;
		Coeff[15523] <= 15'b111111110010000;
		Coeff[15524] <= 15'b111111110010001;
		Coeff[15525] <= 15'b111111110010001;
		Coeff[15526] <= 15'b111111110010001;
		Coeff[15527] <= 15'b111111110010001;
		Coeff[15528] <= 15'b111111110010010;
		Coeff[15529] <= 15'b111111110010010;
		Coeff[15530] <= 15'b111111110010010;
		Coeff[15531] <= 15'b111111110010010;
		Coeff[15532] <= 15'b111111110010011;
		Coeff[15533] <= 15'b111111110010011;
		Coeff[15534] <= 15'b111111110010011;
		Coeff[15535] <= 15'b111111110010100;
		Coeff[15536] <= 15'b111111110010100;
		Coeff[15537] <= 15'b111111110010100;
		Coeff[15538] <= 15'b111111110010100;
		Coeff[15539] <= 15'b111111110010101;
		Coeff[15540] <= 15'b111111110010101;
		Coeff[15541] <= 15'b111111110010101;
		Coeff[15542] <= 15'b111111110010101;
		Coeff[15543] <= 15'b111111110010110;
		Coeff[15544] <= 15'b111111110010110;
		Coeff[15545] <= 15'b111111110010110;
		Coeff[15546] <= 15'b111111110010110;
		Coeff[15547] <= 15'b111111110010111;
		Coeff[15548] <= 15'b111111110010111;
		Coeff[15549] <= 15'b111111110010111;
		Coeff[15550] <= 15'b111111110010111;
		Coeff[15551] <= 15'b111111110011000;
		Coeff[15552] <= 15'b111111110011000;
		Coeff[15553] <= 15'b111111110011000;
		Coeff[15554] <= 15'b111111110011000;
		Coeff[15555] <= 15'b111111110011001;
		Coeff[15556] <= 15'b111111110011001;
		Coeff[15557] <= 15'b111111110011001;
		Coeff[15558] <= 15'b111111110011001;
		Coeff[15559] <= 15'b111111110011010;
		Coeff[15560] <= 15'b111111110011010;
		Coeff[15561] <= 15'b111111110011010;
		Coeff[15562] <= 15'b111111110011010;
		Coeff[15563] <= 15'b111111110011011;
		Coeff[15564] <= 15'b111111110011011;
		Coeff[15565] <= 15'b111111110011011;
		Coeff[15566] <= 15'b111111110011011;
		Coeff[15567] <= 15'b111111110011100;
		Coeff[15568] <= 15'b111111110011100;
		Coeff[15569] <= 15'b111111110011100;
		Coeff[15570] <= 15'b111111110011100;
		Coeff[15571] <= 15'b111111110011101;
		Coeff[15572] <= 15'b111111110011101;
		Coeff[15573] <= 15'b111111110011101;
		Coeff[15574] <= 15'b111111110011101;
		Coeff[15575] <= 15'b111111110011101;
		Coeff[15576] <= 15'b111111110011110;
		Coeff[15577] <= 15'b111111110011110;
		Coeff[15578] <= 15'b111111110011110;
		Coeff[15579] <= 15'b111111110011110;
		Coeff[15580] <= 15'b111111110011111;
		Coeff[15581] <= 15'b111111110011111;
		Coeff[15582] <= 15'b111111110011111;
		Coeff[15583] <= 15'b111111110011111;
		Coeff[15584] <= 15'b111111110100000;
		Coeff[15585] <= 15'b111111110100000;
		Coeff[15586] <= 15'b111111110100000;
		Coeff[15587] <= 15'b111111110100000;
		Coeff[15588] <= 15'b111111110100001;
		Coeff[15589] <= 15'b111111110100001;
		Coeff[15590] <= 15'b111111110100001;
		Coeff[15591] <= 15'b111111110100001;
		Coeff[15592] <= 15'b111111110100010;
		Coeff[15593] <= 15'b111111110100010;
		Coeff[15594] <= 15'b111111110100010;
		Coeff[15595] <= 15'b111111110100010;
		Coeff[15596] <= 15'b111111110100011;
		Coeff[15597] <= 15'b111111110100011;
		Coeff[15598] <= 15'b111111110100011;
		Coeff[15599] <= 15'b111111110100011;
		Coeff[15600] <= 15'b111111110100011;
		Coeff[15601] <= 15'b111111110100100;
		Coeff[15602] <= 15'b111111110100100;
		Coeff[15603] <= 15'b111111110100100;
		Coeff[15604] <= 15'b111111110100100;
		Coeff[15605] <= 15'b111111110100101;
		Coeff[15606] <= 15'b111111110100101;
		Coeff[15607] <= 15'b111111110100101;
		Coeff[15608] <= 15'b111111110100101;
		Coeff[15609] <= 15'b111111110100110;
		Coeff[15610] <= 15'b111111110100110;
		Coeff[15611] <= 15'b111111110100110;
		Coeff[15612] <= 15'b111111110100110;
		Coeff[15613] <= 15'b111111110100111;
		Coeff[15614] <= 15'b111111110100111;
		Coeff[15615] <= 15'b111111110100111;
		Coeff[15616] <= 15'b111111110100111;
		Coeff[15617] <= 15'b111111110100111;
		Coeff[15618] <= 15'b111111110101000;
		Coeff[15619] <= 15'b111111110101000;
		Coeff[15620] <= 15'b111111110101000;
		Coeff[15621] <= 15'b111111110101000;
		Coeff[15622] <= 15'b111111110101001;
		Coeff[15623] <= 15'b111111110101001;
		Coeff[15624] <= 15'b111111110101001;
		Coeff[15625] <= 15'b111111110101001;
		Coeff[15626] <= 15'b111111110101010;
		Coeff[15627] <= 15'b111111110101010;
		Coeff[15628] <= 15'b111111110101010;
		Coeff[15629] <= 15'b111111110101010;
		Coeff[15630] <= 15'b111111110101010;
		Coeff[15631] <= 15'b111111110101011;
		Coeff[15632] <= 15'b111111110101011;
		Coeff[15633] <= 15'b111111110101011;
		Coeff[15634] <= 15'b111111110101011;
		Coeff[15635] <= 15'b111111110101100;
		Coeff[15636] <= 15'b111111110101100;
		Coeff[15637] <= 15'b111111110101100;
		Coeff[15638] <= 15'b111111110101100;
		Coeff[15639] <= 15'b111111110101100;
		Coeff[15640] <= 15'b111111110101101;
		Coeff[15641] <= 15'b111111110101101;
		Coeff[15642] <= 15'b111111110101101;
		Coeff[15643] <= 15'b111111110101101;
		Coeff[15644] <= 15'b111111110101110;
		Coeff[15645] <= 15'b111111110101110;
		Coeff[15646] <= 15'b111111110101110;
		Coeff[15647] <= 15'b111111110101110;
		Coeff[15648] <= 15'b111111110101110;
		Coeff[15649] <= 15'b111111110101111;
		Coeff[15650] <= 15'b111111110101111;
		Coeff[15651] <= 15'b111111110101111;
		Coeff[15652] <= 15'b111111110101111;
		Coeff[15653] <= 15'b111111110110000;
		Coeff[15654] <= 15'b111111110110000;
		Coeff[15655] <= 15'b111111110110000;
		Coeff[15656] <= 15'b111111110110000;
		Coeff[15657] <= 15'b111111110110000;
		Coeff[15658] <= 15'b111111110110001;
		Coeff[15659] <= 15'b111111110110001;
		Coeff[15660] <= 15'b111111110110001;
		Coeff[15661] <= 15'b111111110110001;
		Coeff[15662] <= 15'b111111110110010;
		Coeff[15663] <= 15'b111111110110010;
		Coeff[15664] <= 15'b111111110110010;
		Coeff[15665] <= 15'b111111110110010;
		Coeff[15666] <= 15'b111111110110010;
		Coeff[15667] <= 15'b111111110110011;
		Coeff[15668] <= 15'b111111110110011;
		Coeff[15669] <= 15'b111111110110011;
		Coeff[15670] <= 15'b111111110110011;
		Coeff[15671] <= 15'b111111110110011;
		Coeff[15672] <= 15'b111111110110100;
		Coeff[15673] <= 15'b111111110110100;
		Coeff[15674] <= 15'b111111110110100;
		Coeff[15675] <= 15'b111111110110100;
		Coeff[15676] <= 15'b111111110110101;
		Coeff[15677] <= 15'b111111110110101;
		Coeff[15678] <= 15'b111111110110101;
		Coeff[15679] <= 15'b111111110110101;
		Coeff[15680] <= 15'b111111110110101;
		Coeff[15681] <= 15'b111111110110110;
		Coeff[15682] <= 15'b111111110110110;
		Coeff[15683] <= 15'b111111110110110;
		Coeff[15684] <= 15'b111111110110110;
		Coeff[15685] <= 15'b111111110110110;
		Coeff[15686] <= 15'b111111110110111;
		Coeff[15687] <= 15'b111111110110111;
		Coeff[15688] <= 15'b111111110110111;
		Coeff[15689] <= 15'b111111110110111;
		Coeff[15690] <= 15'b111111110110111;
		Coeff[15691] <= 15'b111111110111000;
		Coeff[15692] <= 15'b111111110111000;
		Coeff[15693] <= 15'b111111110111000;
		Coeff[15694] <= 15'b111111110111000;
		Coeff[15695] <= 15'b111111110111001;
		Coeff[15696] <= 15'b111111110111001;
		Coeff[15697] <= 15'b111111110111001;
		Coeff[15698] <= 15'b111111110111001;
		Coeff[15699] <= 15'b111111110111001;
		Coeff[15700] <= 15'b111111110111010;
		Coeff[15701] <= 15'b111111110111010;
		Coeff[15702] <= 15'b111111110111010;
		Coeff[15703] <= 15'b111111110111010;
		Coeff[15704] <= 15'b111111110111010;
		Coeff[15705] <= 15'b111111110111011;
		Coeff[15706] <= 15'b111111110111011;
		Coeff[15707] <= 15'b111111110111011;
		Coeff[15708] <= 15'b111111110111011;
		Coeff[15709] <= 15'b111111110111011;
		Coeff[15710] <= 15'b111111110111100;
		Coeff[15711] <= 15'b111111110111100;
		Coeff[15712] <= 15'b111111110111100;
		Coeff[15713] <= 15'b111111110111100;
		Coeff[15714] <= 15'b111111110111100;
		Coeff[15715] <= 15'b111111110111101;
		Coeff[15716] <= 15'b111111110111101;
		Coeff[15717] <= 15'b111111110111101;
		Coeff[15718] <= 15'b111111110111101;
		Coeff[15719] <= 15'b111111110111101;
		Coeff[15720] <= 15'b111111110111110;
		Coeff[15721] <= 15'b111111110111110;
		Coeff[15722] <= 15'b111111110111110;
		Coeff[15723] <= 15'b111111110111110;
		Coeff[15724] <= 15'b111111110111110;
		Coeff[15725] <= 15'b111111110111111;
		Coeff[15726] <= 15'b111111110111111;
		Coeff[15727] <= 15'b111111110111111;
		Coeff[15728] <= 15'b111111110111111;
		Coeff[15729] <= 15'b111111110111111;
		Coeff[15730] <= 15'b111111111000000;
		Coeff[15731] <= 15'b111111111000000;
		Coeff[15732] <= 15'b111111111000000;
		Coeff[15733] <= 15'b111111111000000;
		Coeff[15734] <= 15'b111111111000000;
		Coeff[15735] <= 15'b111111111000001;
		Coeff[15736] <= 15'b111111111000001;
		Coeff[15737] <= 15'b111111111000001;
		Coeff[15738] <= 15'b111111111000001;
		Coeff[15739] <= 15'b111111111000001;
		Coeff[15740] <= 15'b111111111000010;
		Coeff[15741] <= 15'b111111111000010;
		Coeff[15742] <= 15'b111111111000010;
		Coeff[15743] <= 15'b111111111000010;
		Coeff[15744] <= 15'b111111111000010;
		Coeff[15745] <= 15'b111111111000011;
		Coeff[15746] <= 15'b111111111000011;
		Coeff[15747] <= 15'b111111111000011;
		Coeff[15748] <= 15'b111111111000011;
		Coeff[15749] <= 15'b111111111000011;
		Coeff[15750] <= 15'b111111111000011;
		Coeff[15751] <= 15'b111111111000100;
		Coeff[15752] <= 15'b111111111000100;
		Coeff[15753] <= 15'b111111111000100;
		Coeff[15754] <= 15'b111111111000100;
		Coeff[15755] <= 15'b111111111000100;
		Coeff[15756] <= 15'b111111111000101;
		Coeff[15757] <= 15'b111111111000101;
		Coeff[15758] <= 15'b111111111000101;
		Coeff[15759] <= 15'b111111111000101;
		Coeff[15760] <= 15'b111111111000101;
		Coeff[15761] <= 15'b111111111000110;
		Coeff[15762] <= 15'b111111111000110;
		Coeff[15763] <= 15'b111111111000110;
		Coeff[15764] <= 15'b111111111000110;
		Coeff[15765] <= 15'b111111111000110;
		Coeff[15766] <= 15'b111111111000110;
		Coeff[15767] <= 15'b111111111000111;
		Coeff[15768] <= 15'b111111111000111;
		Coeff[15769] <= 15'b111111111000111;
		Coeff[15770] <= 15'b111111111000111;
		Coeff[15771] <= 15'b111111111000111;
		Coeff[15772] <= 15'b111111111001000;
		Coeff[15773] <= 15'b111111111001000;
		Coeff[15774] <= 15'b111111111001000;
		Coeff[15775] <= 15'b111111111001000;
		Coeff[15776] <= 15'b111111111001000;
		Coeff[15777] <= 15'b111111111001001;
		Coeff[15778] <= 15'b111111111001001;
		Coeff[15779] <= 15'b111111111001001;
		Coeff[15780] <= 15'b111111111001001;
		Coeff[15781] <= 15'b111111111001001;
		Coeff[15782] <= 15'b111111111001001;
		Coeff[15783] <= 15'b111111111001010;
		Coeff[15784] <= 15'b111111111001010;
		Coeff[15785] <= 15'b111111111001010;
		Coeff[15786] <= 15'b111111111001010;
		Coeff[15787] <= 15'b111111111001010;
		Coeff[15788] <= 15'b111111111001011;
		Coeff[15789] <= 15'b111111111001011;
		Coeff[15790] <= 15'b111111111001011;
		Coeff[15791] <= 15'b111111111001011;
		Coeff[15792] <= 15'b111111111001011;
		Coeff[15793] <= 15'b111111111001011;
		Coeff[15794] <= 15'b111111111001100;
		Coeff[15795] <= 15'b111111111001100;
		Coeff[15796] <= 15'b111111111001100;
		Coeff[15797] <= 15'b111111111001100;
		Coeff[15798] <= 15'b111111111001100;
		Coeff[15799] <= 15'b111111111001100;
		Coeff[15800] <= 15'b111111111001101;
		Coeff[15801] <= 15'b111111111001101;
		Coeff[15802] <= 15'b111111111001101;
		Coeff[15803] <= 15'b111111111001101;
		Coeff[15804] <= 15'b111111111001101;
		Coeff[15805] <= 15'b111111111001110;
		Coeff[15806] <= 15'b111111111001110;
		Coeff[15807] <= 15'b111111111001110;
		Coeff[15808] <= 15'b111111111001110;
		Coeff[15809] <= 15'b111111111001110;
		Coeff[15810] <= 15'b111111111001110;
		Coeff[15811] <= 15'b111111111001111;
		Coeff[15812] <= 15'b111111111001111;
		Coeff[15813] <= 15'b111111111001111;
		Coeff[15814] <= 15'b111111111001111;
		Coeff[15815] <= 15'b111111111001111;
		Coeff[15816] <= 15'b111111111001111;
		Coeff[15817] <= 15'b111111111010000;
		Coeff[15818] <= 15'b111111111010000;
		Coeff[15819] <= 15'b111111111010000;
		Coeff[15820] <= 15'b111111111010000;
		Coeff[15821] <= 15'b111111111010000;
		Coeff[15822] <= 15'b111111111010000;
		Coeff[15823] <= 15'b111111111010001;
		Coeff[15824] <= 15'b111111111010001;
		Coeff[15825] <= 15'b111111111010001;
		Coeff[15826] <= 15'b111111111010001;
		Coeff[15827] <= 15'b111111111010001;
		Coeff[15828] <= 15'b111111111010001;
		Coeff[15829] <= 15'b111111111010010;
		Coeff[15830] <= 15'b111111111010010;
		Coeff[15831] <= 15'b111111111010010;
		Coeff[15832] <= 15'b111111111010010;
		Coeff[15833] <= 15'b111111111010010;
		Coeff[15834] <= 15'b111111111010010;
		Coeff[15835] <= 15'b111111111010011;
		Coeff[15836] <= 15'b111111111010011;
		Coeff[15837] <= 15'b111111111010011;
		Coeff[15838] <= 15'b111111111010011;
		Coeff[15839] <= 15'b111111111010011;
		Coeff[15840] <= 15'b111111111010011;
		Coeff[15841] <= 15'b111111111010100;
		Coeff[15842] <= 15'b111111111010100;
		Coeff[15843] <= 15'b111111111010100;
		Coeff[15844] <= 15'b111111111010100;
		Coeff[15845] <= 15'b111111111010100;
		Coeff[15846] <= 15'b111111111010100;
		Coeff[15847] <= 15'b111111111010101;
		Coeff[15848] <= 15'b111111111010101;
		Coeff[15849] <= 15'b111111111010101;
		Coeff[15850] <= 15'b111111111010101;
		Coeff[15851] <= 15'b111111111010101;
		Coeff[15852] <= 15'b111111111010101;
		Coeff[15853] <= 15'b111111111010110;
		Coeff[15854] <= 15'b111111111010110;
		Coeff[15855] <= 15'b111111111010110;
		Coeff[15856] <= 15'b111111111010110;
		Coeff[15857] <= 15'b111111111010110;
		Coeff[15858] <= 15'b111111111010110;
		Coeff[15859] <= 15'b111111111010111;
		Coeff[15860] <= 15'b111111111010111;
		Coeff[15861] <= 15'b111111111010111;
		Coeff[15862] <= 15'b111111111010111;
		Coeff[15863] <= 15'b111111111010111;
		Coeff[15864] <= 15'b111111111010111;
		Coeff[15865] <= 15'b111111111010111;
		Coeff[15866] <= 15'b111111111011000;
		Coeff[15867] <= 15'b111111111011000;
		Coeff[15868] <= 15'b111111111011000;
		Coeff[15869] <= 15'b111111111011000;
		Coeff[15870] <= 15'b111111111011000;
		Coeff[15871] <= 15'b111111111011000;
		Coeff[15872] <= 15'b111111111011001;
		Coeff[15873] <= 15'b111111111011001;
		Coeff[15874] <= 15'b111111111011001;
		Coeff[15875] <= 15'b111111111011001;
		Coeff[15876] <= 15'b111111111011001;
		Coeff[15877] <= 15'b111111111011001;
		Coeff[15878] <= 15'b111111111011001;
		Coeff[15879] <= 15'b111111111011010;
		Coeff[15880] <= 15'b111111111011010;
		Coeff[15881] <= 15'b111111111011010;
		Coeff[15882] <= 15'b111111111011010;
		Coeff[15883] <= 15'b111111111011010;
		Coeff[15884] <= 15'b111111111011010;
		Coeff[15885] <= 15'b111111111011011;
		Coeff[15886] <= 15'b111111111011011;
		Coeff[15887] <= 15'b111111111011011;
		Coeff[15888] <= 15'b111111111011011;
		Coeff[15889] <= 15'b111111111011011;
		Coeff[15890] <= 15'b111111111011011;
		Coeff[15891] <= 15'b111111111011011;
		Coeff[15892] <= 15'b111111111011100;
		Coeff[15893] <= 15'b111111111011100;
		Coeff[15894] <= 15'b111111111011100;
		Coeff[15895] <= 15'b111111111011100;
		Coeff[15896] <= 15'b111111111011100;
		Coeff[15897] <= 15'b111111111011100;
		Coeff[15898] <= 15'b111111111011100;
		Coeff[15899] <= 15'b111111111011101;
		Coeff[15900] <= 15'b111111111011101;
		Coeff[15901] <= 15'b111111111011101;
		Coeff[15902] <= 15'b111111111011101;
		Coeff[15903] <= 15'b111111111011101;
		Coeff[15904] <= 15'b111111111011101;
		Coeff[15905] <= 15'b111111111011101;
		Coeff[15906] <= 15'b111111111011110;
		Coeff[15907] <= 15'b111111111011110;
		Coeff[15908] <= 15'b111111111011110;
		Coeff[15909] <= 15'b111111111011110;
		Coeff[15910] <= 15'b111111111011110;
		Coeff[15911] <= 15'b111111111011110;
		Coeff[15912] <= 15'b111111111011110;
		Coeff[15913] <= 15'b111111111011111;
		Coeff[15914] <= 15'b111111111011111;
		Coeff[15915] <= 15'b111111111011111;
		Coeff[15916] <= 15'b111111111011111;
		Coeff[15917] <= 15'b111111111011111;
		Coeff[15918] <= 15'b111111111011111;
		Coeff[15919] <= 15'b111111111011111;
		Coeff[15920] <= 15'b111111111100000;
		Coeff[15921] <= 15'b111111111100000;
		Coeff[15922] <= 15'b111111111100000;
		Coeff[15923] <= 15'b111111111100000;
		Coeff[15924] <= 15'b111111111100000;
		Coeff[15925] <= 15'b111111111100000;
		Coeff[15926] <= 15'b111111111100000;
		Coeff[15927] <= 15'b111111111100001;
		Coeff[15928] <= 15'b111111111100001;
		Coeff[15929] <= 15'b111111111100001;
		Coeff[15930] <= 15'b111111111100001;
		Coeff[15931] <= 15'b111111111100001;
		Coeff[15932] <= 15'b111111111100001;
		Coeff[15933] <= 15'b111111111100001;
		Coeff[15934] <= 15'b111111111100010;
		Coeff[15935] <= 15'b111111111100010;
		Coeff[15936] <= 15'b111111111100010;
		Coeff[15937] <= 15'b111111111100010;
		Coeff[15938] <= 15'b111111111100010;
		Coeff[15939] <= 15'b111111111100010;
		Coeff[15940] <= 15'b111111111100010;
		Coeff[15941] <= 15'b111111111100010;
		Coeff[15942] <= 15'b111111111100011;
		Coeff[15943] <= 15'b111111111100011;
		Coeff[15944] <= 15'b111111111100011;
		Coeff[15945] <= 15'b111111111100011;
		Coeff[15946] <= 15'b111111111100011;
		Coeff[15947] <= 15'b111111111100011;
		Coeff[15948] <= 15'b111111111100011;
		Coeff[15949] <= 15'b111111111100100;
		Coeff[15950] <= 15'b111111111100100;
		Coeff[15951] <= 15'b111111111100100;
		Coeff[15952] <= 15'b111111111100100;
		Coeff[15953] <= 15'b111111111100100;
		Coeff[15954] <= 15'b111111111100100;
		Coeff[15955] <= 15'b111111111100100;
		Coeff[15956] <= 15'b111111111100100;
		Coeff[15957] <= 15'b111111111100101;
		Coeff[15958] <= 15'b111111111100101;
		Coeff[15959] <= 15'b111111111100101;
		Coeff[15960] <= 15'b111111111100101;
		Coeff[15961] <= 15'b111111111100101;
		Coeff[15962] <= 15'b111111111100101;
		Coeff[15963] <= 15'b111111111100101;
		Coeff[15964] <= 15'b111111111100101;
		Coeff[15965] <= 15'b111111111100110;
		Coeff[15966] <= 15'b111111111100110;
		Coeff[15967] <= 15'b111111111100110;
		Coeff[15968] <= 15'b111111111100110;
		Coeff[15969] <= 15'b111111111100110;
		Coeff[15970] <= 15'b111111111100110;
		Coeff[15971] <= 15'b111111111100110;
		Coeff[15972] <= 15'b111111111100110;
		Coeff[15973] <= 15'b111111111100111;
		Coeff[15974] <= 15'b111111111100111;
		Coeff[15975] <= 15'b111111111100111;
		Coeff[15976] <= 15'b111111111100111;
		Coeff[15977] <= 15'b111111111100111;
		Coeff[15978] <= 15'b111111111100111;
		Coeff[15979] <= 15'b111111111100111;
		Coeff[15980] <= 15'b111111111100111;
		Coeff[15981] <= 15'b111111111101000;
		Coeff[15982] <= 15'b111111111101000;
		Coeff[15983] <= 15'b111111111101000;
		Coeff[15984] <= 15'b111111111101000;
		Coeff[15985] <= 15'b111111111101000;
		Coeff[15986] <= 15'b111111111101000;
		Coeff[15987] <= 15'b111111111101000;
		Coeff[15988] <= 15'b111111111101000;
		Coeff[15989] <= 15'b111111111101001;
		Coeff[15990] <= 15'b111111111101001;
		Coeff[15991] <= 15'b111111111101001;
		Coeff[15992] <= 15'b111111111101001;
		Coeff[15993] <= 15'b111111111101001;
		Coeff[15994] <= 15'b111111111101001;
		Coeff[15995] <= 15'b111111111101001;
		Coeff[15996] <= 15'b111111111101001;
		Coeff[15997] <= 15'b111111111101001;
		Coeff[15998] <= 15'b111111111101010;
		Coeff[15999] <= 15'b111111111101010;
		Coeff[16000] <= 15'b111111111101010;
		Coeff[16001] <= 15'b111111111101010;
		Coeff[16002] <= 15'b111111111101010;
		Coeff[16003] <= 15'b111111111101010;
		Coeff[16004] <= 15'b111111111101010;
		Coeff[16005] <= 15'b111111111101010;
		Coeff[16006] <= 15'b111111111101010;
		Coeff[16007] <= 15'b111111111101011;
		Coeff[16008] <= 15'b111111111101011;
		Coeff[16009] <= 15'b111111111101011;
		Coeff[16010] <= 15'b111111111101011;
		Coeff[16011] <= 15'b111111111101011;
		Coeff[16012] <= 15'b111111111101011;
		Coeff[16013] <= 15'b111111111101011;
		Coeff[16014] <= 15'b111111111101011;
		Coeff[16015] <= 15'b111111111101011;
		Coeff[16016] <= 15'b111111111101100;
		Coeff[16017] <= 15'b111111111101100;
		Coeff[16018] <= 15'b111111111101100;
		Coeff[16019] <= 15'b111111111101100;
		Coeff[16020] <= 15'b111111111101100;
		Coeff[16021] <= 15'b111111111101100;
		Coeff[16022] <= 15'b111111111101100;
		Coeff[16023] <= 15'b111111111101100;
		Coeff[16024] <= 15'b111111111101100;
		Coeff[16025] <= 15'b111111111101101;
		Coeff[16026] <= 15'b111111111101101;
		Coeff[16027] <= 15'b111111111101101;
		Coeff[16028] <= 15'b111111111101101;
		Coeff[16029] <= 15'b111111111101101;
		Coeff[16030] <= 15'b111111111101101;
		Coeff[16031] <= 15'b111111111101101;
		Coeff[16032] <= 15'b111111111101101;
		Coeff[16033] <= 15'b111111111101101;
		Coeff[16034] <= 15'b111111111101110;
		Coeff[16035] <= 15'b111111111101110;
		Coeff[16036] <= 15'b111111111101110;
		Coeff[16037] <= 15'b111111111101110;
		Coeff[16038] <= 15'b111111111101110;
		Coeff[16039] <= 15'b111111111101110;
		Coeff[16040] <= 15'b111111111101110;
		Coeff[16041] <= 15'b111111111101110;
		Coeff[16042] <= 15'b111111111101110;
		Coeff[16043] <= 15'b111111111101110;
		Coeff[16044] <= 15'b111111111101111;
		Coeff[16045] <= 15'b111111111101111;
		Coeff[16046] <= 15'b111111111101111;
		Coeff[16047] <= 15'b111111111101111;
		Coeff[16048] <= 15'b111111111101111;
		Coeff[16049] <= 15'b111111111101111;
		Coeff[16050] <= 15'b111111111101111;
		Coeff[16051] <= 15'b111111111101111;
		Coeff[16052] <= 15'b111111111101111;
		Coeff[16053] <= 15'b111111111110000;
		Coeff[16054] <= 15'b111111111110000;
		Coeff[16055] <= 15'b111111111110000;
		Coeff[16056] <= 15'b111111111110000;
		Coeff[16057] <= 15'b111111111110000;
		Coeff[16058] <= 15'b111111111110000;
		Coeff[16059] <= 15'b111111111110000;
		Coeff[16060] <= 15'b111111111110000;
		Coeff[16061] <= 15'b111111111110000;
		Coeff[16062] <= 15'b111111111110000;
		Coeff[16063] <= 15'b111111111110000;
		Coeff[16064] <= 15'b111111111110001;
		Coeff[16065] <= 15'b111111111110001;
		Coeff[16066] <= 15'b111111111110001;
		Coeff[16067] <= 15'b111111111110001;
		Coeff[16068] <= 15'b111111111110001;
		Coeff[16069] <= 15'b111111111110001;
		Coeff[16070] <= 15'b111111111110001;
		Coeff[16071] <= 15'b111111111110001;
		Coeff[16072] <= 15'b111111111110001;
		Coeff[16073] <= 15'b111111111110001;
		Coeff[16074] <= 15'b111111111110010;
		Coeff[16075] <= 15'b111111111110010;
		Coeff[16076] <= 15'b111111111110010;
		Coeff[16077] <= 15'b111111111110010;
		Coeff[16078] <= 15'b111111111110010;
		Coeff[16079] <= 15'b111111111110010;
		Coeff[16080] <= 15'b111111111110010;
		Coeff[16081] <= 15'b111111111110010;
		Coeff[16082] <= 15'b111111111110010;
		Coeff[16083] <= 15'b111111111110010;
		Coeff[16084] <= 15'b111111111110010;
		Coeff[16085] <= 15'b111111111110011;
		Coeff[16086] <= 15'b111111111110011;
		Coeff[16087] <= 15'b111111111110011;
		Coeff[16088] <= 15'b111111111110011;
		Coeff[16089] <= 15'b111111111110011;
		Coeff[16090] <= 15'b111111111110011;
		Coeff[16091] <= 15'b111111111110011;
		Coeff[16092] <= 15'b111111111110011;
		Coeff[16093] <= 15'b111111111110011;
		Coeff[16094] <= 15'b111111111110011;
		Coeff[16095] <= 15'b111111111110011;
		Coeff[16096] <= 15'b111111111110100;
		Coeff[16097] <= 15'b111111111110100;
		Coeff[16098] <= 15'b111111111110100;
		Coeff[16099] <= 15'b111111111110100;
		Coeff[16100] <= 15'b111111111110100;
		Coeff[16101] <= 15'b111111111110100;
		Coeff[16102] <= 15'b111111111110100;
		Coeff[16103] <= 15'b111111111110100;
		Coeff[16104] <= 15'b111111111110100;
		Coeff[16105] <= 15'b111111111110100;
		Coeff[16106] <= 15'b111111111110100;
		Coeff[16107] <= 15'b111111111110100;
		Coeff[16108] <= 15'b111111111110101;
		Coeff[16109] <= 15'b111111111110101;
		Coeff[16110] <= 15'b111111111110101;
		Coeff[16111] <= 15'b111111111110101;
		Coeff[16112] <= 15'b111111111110101;
		Coeff[16113] <= 15'b111111111110101;
		Coeff[16114] <= 15'b111111111110101;
		Coeff[16115] <= 15'b111111111110101;
		Coeff[16116] <= 15'b111111111110101;
		Coeff[16117] <= 15'b111111111110101;
		Coeff[16118] <= 15'b111111111110101;
		Coeff[16119] <= 15'b111111111110101;
		Coeff[16120] <= 15'b111111111110110;
		Coeff[16121] <= 15'b111111111110110;
		Coeff[16122] <= 15'b111111111110110;
		Coeff[16123] <= 15'b111111111110110;
		Coeff[16124] <= 15'b111111111110110;
		Coeff[16125] <= 15'b111111111110110;
		Coeff[16126] <= 15'b111111111110110;
		Coeff[16127] <= 15'b111111111110110;
		Coeff[16128] <= 15'b111111111110110;
		Coeff[16129] <= 15'b111111111110110;
		Coeff[16130] <= 15'b111111111110110;
		Coeff[16131] <= 15'b111111111110110;
		Coeff[16132] <= 15'b111111111110110;
		Coeff[16133] <= 15'b111111111110111;
		Coeff[16134] <= 15'b111111111110111;
		Coeff[16135] <= 15'b111111111110111;
		Coeff[16136] <= 15'b111111111110111;
		Coeff[16137] <= 15'b111111111110111;
		Coeff[16138] <= 15'b111111111110111;
		Coeff[16139] <= 15'b111111111110111;
		Coeff[16140] <= 15'b111111111110111;
		Coeff[16141] <= 15'b111111111110111;
		Coeff[16142] <= 15'b111111111110111;
		Coeff[16143] <= 15'b111111111110111;
		Coeff[16144] <= 15'b111111111110111;
		Coeff[16145] <= 15'b111111111110111;
		Coeff[16146] <= 15'b111111111110111;
		Coeff[16147] <= 15'b111111111111000;
		Coeff[16148] <= 15'b111111111111000;
		Coeff[16149] <= 15'b111111111111000;
		Coeff[16150] <= 15'b111111111111000;
		Coeff[16151] <= 15'b111111111111000;
		Coeff[16152] <= 15'b111111111111000;
		Coeff[16153] <= 15'b111111111111000;
		Coeff[16154] <= 15'b111111111111000;
		Coeff[16155] <= 15'b111111111111000;
		Coeff[16156] <= 15'b111111111111000;
		Coeff[16157] <= 15'b111111111111000;
		Coeff[16158] <= 15'b111111111111000;
		Coeff[16159] <= 15'b111111111111000;
		Coeff[16160] <= 15'b111111111111000;
		Coeff[16161] <= 15'b111111111111001;
		Coeff[16162] <= 15'b111111111111001;
		Coeff[16163] <= 15'b111111111111001;
		Coeff[16164] <= 15'b111111111111001;
		Coeff[16165] <= 15'b111111111111001;
		Coeff[16166] <= 15'b111111111111001;
		Coeff[16167] <= 15'b111111111111001;
		Coeff[16168] <= 15'b111111111111001;
		Coeff[16169] <= 15'b111111111111001;
		Coeff[16170] <= 15'b111111111111001;
		Coeff[16171] <= 15'b111111111111001;
		Coeff[16172] <= 15'b111111111111001;
		Coeff[16173] <= 15'b111111111111001;
		Coeff[16174] <= 15'b111111111111001;
		Coeff[16175] <= 15'b111111111111001;
		Coeff[16176] <= 15'b111111111111001;
		Coeff[16177] <= 15'b111111111111010;
		Coeff[16178] <= 15'b111111111111010;
		Coeff[16179] <= 15'b111111111111010;
		Coeff[16180] <= 15'b111111111111010;
		Coeff[16181] <= 15'b111111111111010;
		Coeff[16182] <= 15'b111111111111010;
		Coeff[16183] <= 15'b111111111111010;
		Coeff[16184] <= 15'b111111111111010;
		Coeff[16185] <= 15'b111111111111010;
		Coeff[16186] <= 15'b111111111111010;
		Coeff[16187] <= 15'b111111111111010;
		Coeff[16188] <= 15'b111111111111010;
		Coeff[16189] <= 15'b111111111111010;
		Coeff[16190] <= 15'b111111111111010;
		Coeff[16191] <= 15'b111111111111010;
		Coeff[16192] <= 15'b111111111111010;
		Coeff[16193] <= 15'b111111111111011;
		Coeff[16194] <= 15'b111111111111011;
		Coeff[16195] <= 15'b111111111111011;
		Coeff[16196] <= 15'b111111111111011;
		Coeff[16197] <= 15'b111111111111011;
		Coeff[16198] <= 15'b111111111111011;
		Coeff[16199] <= 15'b111111111111011;
		Coeff[16200] <= 15'b111111111111011;
		Coeff[16201] <= 15'b111111111111011;
		Coeff[16202] <= 15'b111111111111011;
		Coeff[16203] <= 15'b111111111111011;
		Coeff[16204] <= 15'b111111111111011;
		Coeff[16205] <= 15'b111111111111011;
		Coeff[16206] <= 15'b111111111111011;
		Coeff[16207] <= 15'b111111111111011;
		Coeff[16208] <= 15'b111111111111011;
		Coeff[16209] <= 15'b111111111111011;
		Coeff[16210] <= 15'b111111111111011;
		Coeff[16211] <= 15'b111111111111011;
		Coeff[16212] <= 15'b111111111111100;
		Coeff[16213] <= 15'b111111111111100;
		Coeff[16214] <= 15'b111111111111100;
		Coeff[16215] <= 15'b111111111111100;
		Coeff[16216] <= 15'b111111111111100;
		Coeff[16217] <= 15'b111111111111100;
		Coeff[16218] <= 15'b111111111111100;
		Coeff[16219] <= 15'b111111111111100;
		Coeff[16220] <= 15'b111111111111100;
		Coeff[16221] <= 15'b111111111111100;
		Coeff[16222] <= 15'b111111111111100;
		Coeff[16223] <= 15'b111111111111100;
		Coeff[16224] <= 15'b111111111111100;
		Coeff[16225] <= 15'b111111111111100;
		Coeff[16226] <= 15'b111111111111100;
		Coeff[16227] <= 15'b111111111111100;
		Coeff[16228] <= 15'b111111111111100;
		Coeff[16229] <= 15'b111111111111100;
		Coeff[16230] <= 15'b111111111111100;
		Coeff[16231] <= 15'b111111111111100;
		Coeff[16232] <= 15'b111111111111101;
		Coeff[16233] <= 15'b111111111111101;
		Coeff[16234] <= 15'b111111111111101;
		Coeff[16235] <= 15'b111111111111101;
		Coeff[16236] <= 15'b111111111111101;
		Coeff[16237] <= 15'b111111111111101;
		Coeff[16238] <= 15'b111111111111101;
		Coeff[16239] <= 15'b111111111111101;
		Coeff[16240] <= 15'b111111111111101;
		Coeff[16241] <= 15'b111111111111101;
		Coeff[16242] <= 15'b111111111111101;
		Coeff[16243] <= 15'b111111111111101;
		Coeff[16244] <= 15'b111111111111101;
		Coeff[16245] <= 15'b111111111111101;
		Coeff[16246] <= 15'b111111111111101;
		Coeff[16247] <= 15'b111111111111101;
		Coeff[16248] <= 15'b111111111111101;
		Coeff[16249] <= 15'b111111111111101;
		Coeff[16250] <= 15'b111111111111101;
		Coeff[16251] <= 15'b111111111111101;
		Coeff[16252] <= 15'b111111111111101;
		Coeff[16253] <= 15'b111111111111101;
		Coeff[16254] <= 15'b111111111111101;
		Coeff[16255] <= 15'b111111111111101;
		Coeff[16256] <= 15'b111111111111110;
		Coeff[16257] <= 15'b111111111111110;
		Coeff[16258] <= 15'b111111111111110;
		Coeff[16259] <= 15'b111111111111110;
		Coeff[16260] <= 15'b111111111111110;
		Coeff[16261] <= 15'b111111111111110;
		Coeff[16262] <= 15'b111111111111110;
		Coeff[16263] <= 15'b111111111111110;
		Coeff[16264] <= 15'b111111111111110;
		Coeff[16265] <= 15'b111111111111110;
		Coeff[16266] <= 15'b111111111111110;
		Coeff[16267] <= 15'b111111111111110;
		Coeff[16268] <= 15'b111111111111110;
		Coeff[16269] <= 15'b111111111111110;
		Coeff[16270] <= 15'b111111111111110;
		Coeff[16271] <= 15'b111111111111110;
		Coeff[16272] <= 15'b111111111111110;
		Coeff[16273] <= 15'b111111111111110;
		Coeff[16274] <= 15'b111111111111110;
		Coeff[16275] <= 15'b111111111111110;
		Coeff[16276] <= 15'b111111111111110;
		Coeff[16277] <= 15'b111111111111110;
		Coeff[16278] <= 15'b111111111111110;
		Coeff[16279] <= 15'b111111111111110;
		Coeff[16280] <= 15'b111111111111110;
		Coeff[16281] <= 15'b111111111111110;
		Coeff[16282] <= 15'b111111111111110;
		Coeff[16283] <= 15'b111111111111110;
		Coeff[16284] <= 15'b111111111111110;
		Coeff[16285] <= 15'b111111111111111;
		Coeff[16286] <= 15'b111111111111111;
		Coeff[16287] <= 15'b111111111111111;
		Coeff[16288] <= 15'b111111111111111;
		Coeff[16289] <= 15'b111111111111111;
		Coeff[16290] <= 15'b111111111111111;
		Coeff[16291] <= 15'b111111111111111;
		Coeff[16292] <= 15'b111111111111111;
		Coeff[16293] <= 15'b111111111111111;
		Coeff[16294] <= 15'b111111111111111;
		Coeff[16295] <= 15'b111111111111111;
		Coeff[16296] <= 15'b111111111111111;
		Coeff[16297] <= 15'b111111111111111;
		Coeff[16298] <= 15'b111111111111111;
		Coeff[16299] <= 15'b111111111111111;
		Coeff[16300] <= 15'b111111111111111;
		Coeff[16301] <= 15'b111111111111111;
		Coeff[16302] <= 15'b111111111111111;
		Coeff[16303] <= 15'b111111111111111;
		Coeff[16304] <= 15'b111111111111111;
		Coeff[16305] <= 15'b111111111111111;
		Coeff[16306] <= 15'b111111111111111;
		Coeff[16307] <= 15'b111111111111111;
		Coeff[16308] <= 15'b111111111111111;
		Coeff[16309] <= 15'b111111111111111;
		Coeff[16310] <= 15'b111111111111111;
		Coeff[16311] <= 15'b111111111111111;
		Coeff[16312] <= 15'b111111111111111;
		Coeff[16313] <= 15'b111111111111111;
		Coeff[16314] <= 15'b111111111111111;
		Coeff[16315] <= 15'b111111111111111;
		Coeff[16316] <= 15'b111111111111111;
		Coeff[16317] <= 15'b111111111111111;
		Coeff[16318] <= 15'b111111111111111;
		Coeff[16319] <= 15'b111111111111111;
		Coeff[16320] <= 15'b111111111111111;
		Coeff[16321] <= 15'b111111111111111;
		Coeff[16322] <= 15'b111111111111111;
		Coeff[16323] <= 15'b111111111111111;
		Coeff[16324] <= 15'b111111111111111;
		Coeff[16325] <= 15'b111111111111111;
		Coeff[16326] <= 15'b111111111111111;
		Coeff[16327] <= 15'b111111111111111;
		Coeff[16328] <= 15'b111111111111111;
		Coeff[16329] <= 15'b111111111111111;
		Coeff[16330] <= 15'b111111111111111;
		Coeff[16331] <= 15'b111111111111111;
		Coeff[16332] <= 15'b111111111111111;
		Coeff[16333] <= 15'b111111111111111;
		Coeff[16334] <= 15'b111111111111111;
		Coeff[16335] <= 15'b111111111111111;
		Coeff[16336] <= 15'b111111111111111;
		Coeff[16337] <= 15'b111111111111111;
		Coeff[16338] <= 15'b111111111111111;
		Coeff[16339] <= 15'b111111111111111;
		Coeff[16340] <= 15'b111111111111111;
		Coeff[16341] <= 15'b111111111111111;
		Coeff[16342] <= 15'b111111111111111;
		Coeff[16343] <= 15'b111111111111111;
		Coeff[16344] <= 15'b111111111111111;
		Coeff[16345] <= 15'b111111111111111;
		Coeff[16346] <= 15'b111111111111111;
		Coeff[16347] <= 15'b111111111111111;
		Coeff[16348] <= 15'b111111111111111;
		Coeff[16349] <= 15'b111111111111111;
		Coeff[16350] <= 15'b111111111111111;
		Coeff[16351] <= 15'b111111111111111;
		Coeff[16352] <= 15'b111111111111111;
		Coeff[16353] <= 15'b111111111111111;
		Coeff[16354] <= 15'b111111111111111;
		Coeff[16355] <= 15'b111111111111111;
		Coeff[16356] <= 15'b111111111111111;
		Coeff[16357] <= 15'b111111111111111;
		Coeff[16358] <= 15'b111111111111111;
		Coeff[16359] <= 15'b111111111111111;
		Coeff[16360] <= 15'b111111111111111;
		Coeff[16361] <= 15'b111111111111111;
		Coeff[16362] <= 15'b111111111111111;
		Coeff[16363] <= 15'b111111111111111;
		Coeff[16364] <= 15'b111111111111111;
		Coeff[16365] <= 15'b111111111111111;
		Coeff[16366] <= 15'b111111111111111;
		Coeff[16367] <= 15'b111111111111111;
		Coeff[16368] <= 15'b111111111111111;
		Coeff[16369] <= 15'b111111111111111;
		Coeff[16370] <= 15'b111111111111111;
		Coeff[16371] <= 15'b111111111111111;
		Coeff[16372] <= 15'b111111111111111;
		Coeff[16373] <= 15'b111111111111111;
		Coeff[16374] <= 15'b111111111111111;
		Coeff[16375] <= 15'b111111111111111;
		Coeff[16376] <= 15'b111111111111111;
		Coeff[16377] <= 15'b111111111111111;
		Coeff[16378] <= 15'b111111111111111;
		Coeff[16379] <= 15'b111111111111111;
		Coeff[16380] <= 15'b111111111111111;
		Coeff[16381] <= 15'b111111111111111;
		Coeff[16382] <= 15'b111111111111111;
		Coeff[16383] <= 15'b111111111111111;
	
	end
end

endmodule
