/* Module to calculate sin of the input signal (16,16) bits 

Func - 	0 for sine
	1 for Cosine

Latency = 2 clock cycle

*/

module SinBlock(input clk, input reset, input func, input [15:0] x, output reg [15:0] sinValue);

reg [11:0] Sin_C1[128];
reg [18:0] Sin_C0[128];

reg [25:0] Term1;
reg [32:0] Term2;
reg sValue;

always @(posedge clk)
begin
	if(!reset)
	begin
		
		// Cycle 1
		Term1 <= Sin_C1[x[14:8]] * x[13:0];
		Term2 <= Sin_C0[x[14:8]];

		// Cycle 2
		sinValue [14:0] <= Term1[25:11] + Term2[32:18];
		sinValue [15] <= sValue;

		case( {func, x[15:14]} )
		// Sine Calculation
	
		3'b000 : begin
				sValue <= 1'b0;
			end

		3'b001 : begin
				sValue <= 1'b0;
			end
	
		3'b010 : begin
				sValue <= 1'b1;
			end
	
		3'b011 : begin
				sValue <= 1'b1;
			end

		// Cosine Calculation

		3'b100 : begin
				sValue <= 1'b0;
			end

		3'b101 : begin
				sValue <= 1'b1;
			end

		3'b110 : begin
				sValue <= 1'b1;
			end
	
		3'b111 : begin
				sValue <= 1'b0;
			end	

		endcase


	end // reset

	else
	begin

		Sin_C0[0] <= 19'b1000000000000000011;
		Sin_C0[1] <= 19'b1000000000000101011;
		Sin_C0[2] <= 19'b1000000000001111010;
		Sin_C0[3] <= 19'b1000000000011110000;
		Sin_C0[4] <= 19'b1000000000110001110;
		Sin_C0[5] <= 19'b1000000001001010011;
		Sin_C0[6] <= 19'b1000000001100111111;
		Sin_C0[7] <= 19'b1000000010001010010;
		Sin_C0[8] <= 19'b1000000010110001101;
		Sin_C0[9] <= 19'b1000000011011101110;
		Sin_C0[10] <= 19'b1000000100001110110;
		Sin_C0[11] <= 19'b1000000101000100100;
		Sin_C0[12] <= 19'b1000000101111111000;
		Sin_C0[13] <= 19'b1000000110111110011;
		Sin_C0[14] <= 19'b1000001000000010100;
		Sin_C0[15] <= 19'b1000001001001011010;
		Sin_C0[16] <= 19'b1000001010011000101;
		Sin_C0[17] <= 19'b1000001011101010110;
		Sin_C0[18] <= 19'b1000001101000001011;
		Sin_C0[19] <= 19'b1000001110011100101;
		Sin_C0[20] <= 19'b1000001111111100011;
		Sin_C0[21] <= 19'b1000010001100000101;
		Sin_C0[22] <= 19'b1000010011001001010;
		Sin_C0[23] <= 19'b1000010100110110010;
		Sin_C0[24] <= 19'b1000010110100111100;
		Sin_C0[25] <= 19'b1000011000011101001;
		Sin_C0[26] <= 19'b1000011010010111000;
		Sin_C0[27] <= 19'b1000011100010101000;
		Sin_C0[28] <= 19'b1000011110010111000;
		Sin_C0[29] <= 19'b1000100000011101010;
		Sin_C0[30] <= 19'b1000100010100111011;
		Sin_C0[31] <= 19'b1000100100110101011;
		Sin_C0[32] <= 19'b1000100111000111010;
		Sin_C0[33] <= 19'b1000101001011100111;
		Sin_C0[34] <= 19'b1000101011110110010;
		Sin_C0[35] <= 19'b1000101110010011011;
		Sin_C0[36] <= 19'b1000110000110011111;
		Sin_C0[37] <= 19'b1000110011011000000;
		Sin_C0[38] <= 19'b1000110101111111100;
		Sin_C0[39] <= 19'b1000111000101010011;
		Sin_C0[40] <= 19'b1000111011011000011;
		Sin_C0[41] <= 19'b1000111110001001101;
		Sin_C0[42] <= 19'b1001000000111110000;
		Sin_C0[43] <= 19'b1001000011110101011;
		Sin_C0[44] <= 19'b1001000110101111100;
		Sin_C0[45] <= 19'b1001001001101100101;
		Sin_C0[46] <= 19'b1001001100101100011;
		Sin_C0[47] <= 19'b1001001111101110110;
		Sin_C0[48] <= 19'b1001010010110011110;
		Sin_C0[49] <= 19'b1001010101111011001;
		Sin_C0[50] <= 19'b1001011001000100111;
		Sin_C0[51] <= 19'b1001011100010000111;
		Sin_C0[52] <= 19'b1001011111011110111;
		Sin_C0[53] <= 19'b1001100010101111001;
		Sin_C0[54] <= 19'b1001100110000001001;
		Sin_C0[55] <= 19'b1001101001010101000;
		Sin_C0[56] <= 19'b1001101100101010101;
		Sin_C0[57] <= 19'b1001110000000001111;
		Sin_C0[58] <= 19'b1001110011011010101;
		Sin_C0[59] <= 19'b1001110110110100110;
		Sin_C0[60] <= 19'b1001111010010000001;
		Sin_C0[61] <= 19'b1001111101101100101;
		Sin_C0[62] <= 19'b1010000001001010010;
		Sin_C0[63] <= 19'b1010000100101000110;
		Sin_C0[64] <= 19'b1010001000001000000;
		Sin_C0[65] <= 19'b1010001011101000001;
		Sin_C0[66] <= 19'b1010001111001000101;
		Sin_C0[67] <= 19'b1010010010101001101;
		Sin_C0[68] <= 19'b1010010110001011000;
		Sin_C0[69] <= 19'b1010011001101100100;
		Sin_C0[70] <= 19'b1010011101001110001;
		Sin_C0[71] <= 19'b1010100000101111110;
		Sin_C0[72] <= 19'b1010100100010001001;
		Sin_C0[73] <= 19'b1010100111110010010;
		Sin_C0[74] <= 19'b1010101011010010111;
		Sin_C0[75] <= 19'b1010101110110011000;
		Sin_C0[76] <= 19'b1010110010010010011;
		Sin_C0[77] <= 19'b1010110101110001000;
		Sin_C0[78] <= 19'b1010111001001110101;
		Sin_C0[79] <= 19'b1010111100101011001;
		Sin_C0[80] <= 19'b1011000000000110100;
		Sin_C0[81] <= 19'b1011000011100000100;
		Sin_C0[82] <= 19'b1011000110111001000;
		Sin_C0[83] <= 19'b1011001010001111111;
		Sin_C0[84] <= 19'b1011001101100100111;
		Sin_C0[85] <= 19'b1011010000111000001;
		Sin_C0[86] <= 19'b1011010100001001010;
		Sin_C0[87] <= 19'b1011010111011000011;
		Sin_C0[88] <= 19'b1011011010100101000;
		Sin_C0[89] <= 19'b1011011101101111010;
		Sin_C0[90] <= 19'b1011100000110111000;
		Sin_C0[91] <= 19'b1011100011111011111;
		Sin_C0[92] <= 19'b1011100110111110000;
		Sin_C0[93] <= 19'b1011101001111101001;
		Sin_C0[94] <= 19'b1011101100111001001;
		Sin_C0[95] <= 19'b1011101111110001111;
		Sin_C0[96] <= 19'b1011110010100111001;
		Sin_C0[97] <= 19'b1011110101011000111;
		Sin_C0[98] <= 19'b1011111000000110111;
		Sin_C0[99] <= 19'b1011111010110001001;
		Sin_C0[100] <= 19'b1011111101010111011;
		Sin_C0[101] <= 19'b1011111111111001100;
		Sin_C0[102] <= 19'b1100000010010111011;
		Sin_C0[103] <= 19'b1100000100110000111;
		Sin_C0[104] <= 19'b1100000111000101111;
		Sin_C0[105] <= 19'b1100001001010110001;
		Sin_C0[106] <= 19'b1100001011100001101;
		Sin_C0[107] <= 19'b1100001101101000010;
		Sin_C0[108] <= 19'b1100001111101001110;
		Sin_C0[109] <= 19'b1100010001100110000;
		Sin_C0[110] <= 19'b1100010011011100111;
		Sin_C0[111] <= 19'b1100010101001110011;
		Sin_C0[112] <= 19'b1100010110111010010;
		Sin_C0[113] <= 19'b1100011000100000010;
		Sin_C0[114] <= 19'b1100011010000000011;
		Sin_C0[115] <= 19'b1100011011011010101;
		Sin_C0[116] <= 19'b1100011100101110100;
		Sin_C0[117] <= 19'b1100011101111100010;
		Sin_C0[118] <= 19'b1100011111000011100;
		Sin_C0[119] <= 19'b1100100000000100010;
		Sin_C0[120] <= 19'b1100100000111110010;
		Sin_C0[121] <= 19'b1100100001110001100;
		Sin_C0[122] <= 19'b1100100010011101110;
		Sin_C0[123] <= 19'b1100100011000011000;
		Sin_C0[124] <= 19'b1100100011100001000;
		Sin_C0[125] <= 19'b1100100011110111110;
		Sin_C0[126] <= 19'b1100100100000111000;
		Sin_C0[127] <= 19'b1100100100001110101;

		Sin_C1[0] <= 12'b000000001101;
		Sin_C1[1] <= 12'b000000100110;
		Sin_C1[2] <= 12'b000000111111;
		Sin_C1[3] <= 12'b000001011000;
		Sin_C1[4] <= 12'b000001110001;
		Sin_C1[5] <= 12'b000010001010;
		Sin_C1[6] <= 12'b000010100011;
		Sin_C1[7] <= 12'b000010111100;
		Sin_C1[8] <= 12'b000011010101;
		Sin_C1[9] <= 12'b000011101110;
		Sin_C1[10] <= 12'b000100000111;
		Sin_C1[11] <= 12'b000100100000;
		Sin_C1[12] <= 12'b000100111001;
		Sin_C1[13] <= 12'b000101010010;
		Sin_C1[14] <= 12'b000101101011;
		Sin_C1[15] <= 12'b000110000011;
		Sin_C1[16] <= 12'b000110011100;
		Sin_C1[17] <= 12'b000110110100;
		Sin_C1[18] <= 12'b000111001101;
		Sin_C1[19] <= 12'b000111100101;
		Sin_C1[20] <= 12'b000111111110;
		Sin_C1[21] <= 12'b001000010110;
		Sin_C1[22] <= 12'b001000101110;
		Sin_C1[23] <= 12'b001001000110;
		Sin_C1[24] <= 12'b001001011111;
		Sin_C1[25] <= 12'b001001110110;
		Sin_C1[26] <= 12'b001010001110;
		Sin_C1[27] <= 12'b001010100110;
		Sin_C1[28] <= 12'b001010111110;
		Sin_C1[29] <= 12'b001011010101;
		Sin_C1[30] <= 12'b001011101101;
		Sin_C1[31] <= 12'b001100000100;
		Sin_C1[32] <= 12'b001100011011;
		Sin_C1[33] <= 12'b001100110010;
		Sin_C1[34] <= 12'b001101001001;
		Sin_C1[35] <= 12'b001101100000;
		Sin_C1[36] <= 12'b001101110111;
		Sin_C1[37] <= 12'b001110001110;
		Sin_C1[38] <= 12'b001110100100;
		Sin_C1[39] <= 12'b001110111010;
		Sin_C1[40] <= 12'b001111010000;
		Sin_C1[41] <= 12'b001111100110;
		Sin_C1[42] <= 12'b001111111100;
		Sin_C1[43] <= 12'b010000010010;
		Sin_C1[44] <= 12'b010000101000;
		Sin_C1[45] <= 12'b010000111101;
		Sin_C1[46] <= 12'b010001010010;
		Sin_C1[47] <= 12'b010001100111;
		Sin_C1[48] <= 12'b010001111100;
		Sin_C1[49] <= 12'b010010010001;
		Sin_C1[50] <= 12'b010010100110;
		Sin_C1[51] <= 12'b010010111010;
		Sin_C1[52] <= 12'b010011001110;
		Sin_C1[53] <= 12'b010011100010;
		Sin_C1[54] <= 12'b010011110110;
		Sin_C1[55] <= 12'b010100001001;
		Sin_C1[56] <= 12'b010100011101;
		Sin_C1[57] <= 12'b010100110000;
		Sin_C1[58] <= 12'b010101000011;
		Sin_C1[59] <= 12'b010101010110;
		Sin_C1[60] <= 12'b010101101001;
		Sin_C1[61] <= 12'b010101111011;
		Sin_C1[62] <= 12'b010110001101;
		Sin_C1[63] <= 12'b010110011111;
		Sin_C1[64] <= 12'b010110110001;
		Sin_C1[65] <= 12'b010111000011;
		Sin_C1[66] <= 12'b010111010100;
		Sin_C1[67] <= 12'b010111100101;
		Sin_C1[68] <= 12'b010111110110;
		Sin_C1[69] <= 12'b011000000111;
		Sin_C1[70] <= 12'b011000010111;
		Sin_C1[71] <= 12'b011000100111;
		Sin_C1[72] <= 12'b011000110111;
		Sin_C1[73] <= 12'b011001000111;
		Sin_C1[74] <= 12'b011001010110;
		Sin_C1[75] <= 12'b011001100101;
		Sin_C1[76] <= 12'b011001110100;
		Sin_C1[77] <= 12'b011010000011;
		Sin_C1[78] <= 12'b011010010010;
		Sin_C1[79] <= 12'b011010100000;
		Sin_C1[80] <= 12'b011010101110;
		Sin_C1[81] <= 12'b011010111011;
		Sin_C1[82] <= 12'b011011001001;
		Sin_C1[83] <= 12'b011011010110;
		Sin_C1[84] <= 12'b011011100011;
		Sin_C1[85] <= 12'b011011110000;
		Sin_C1[86] <= 12'b011011111100;
		Sin_C1[87] <= 12'b011100001000;
		Sin_C1[88] <= 12'b011100010100;
		Sin_C1[89] <= 12'b011100100000;
		Sin_C1[90] <= 12'b011100101011;
		Sin_C1[91] <= 12'b011100110110;
		Sin_C1[92] <= 12'b011101000001;
		Sin_C1[93] <= 12'b011101001011;
		Sin_C1[94] <= 12'b011101010101;
		Sin_C1[95] <= 12'b011101011111;
		Sin_C1[96] <= 12'b011101101001;
		Sin_C1[97] <= 12'b011101110010;
		Sin_C1[98] <= 12'b011101111011;
		Sin_C1[99] <= 12'b011110000100;
		Sin_C1[100] <= 12'b011110001100;
		Sin_C1[101] <= 12'b011110010101;
		Sin_C1[102] <= 12'b011110011101;
		Sin_C1[103] <= 12'b011110100100;
		Sin_C1[104] <= 12'b011110101011;
		Sin_C1[105] <= 12'b011110110010;
		Sin_C1[106] <= 12'b011110111001;
		Sin_C1[107] <= 12'b011111000000;
		Sin_C1[108] <= 12'b011111000110;
		Sin_C1[109] <= 12'b011111001011;
		Sin_C1[110] <= 12'b011111010001;
		Sin_C1[111] <= 12'b011111010110;
		Sin_C1[112] <= 12'b011111011011;
		Sin_C1[113] <= 12'b011111100000;
		Sin_C1[114] <= 12'b011111100100;
		Sin_C1[115] <= 12'b011111101000;
		Sin_C1[116] <= 12'b011111101100;
		Sin_C1[117] <= 12'b011111101111;
		Sin_C1[118] <= 12'b011111110010;
		Sin_C1[119] <= 12'b011111110101;
		Sin_C1[120] <= 12'b011111110111;
		Sin_C1[121] <= 12'b011111111001;
		Sin_C1[122] <= 12'b011111111011;
		Sin_C1[123] <= 12'b011111111101;
		Sin_C1[124] <= 12'b011111111110;
		Sin_C1[125] <= 12'b011111111111;
		Sin_C1[126] <= 12'b100000000000;
		Sin_C1[127] <= 12'b100000000000;
	end
end

endmodule
